-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTranspose is -- 
  generic (tag_length : integer); 
  port ( -- 
    Block0_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block0_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block0_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block1_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block1_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block1_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block2_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block2_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block2_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block3_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block3_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block3_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block1_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block1_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block1_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    Block0_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block0_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block0_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    Block3_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block3_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block3_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    Block2_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block2_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block2_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    elapsed_time_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_write_data : out  std_logic_vector(63 downto 0);
    testConfigure_call_reqs : out  std_logic_vector(0 downto 0);
    testConfigure_call_acks : in   std_logic_vector(0 downto 0);
    testConfigure_call_tag  :  out  std_logic_vector(0 downto 0);
    testConfigure_return_reqs : out  std_logic_vector(0 downto 0);
    testConfigure_return_acks : in   std_logic_vector(0 downto 0);
    testConfigure_return_data : in   std_logic_vector(15 downto 0);
    testConfigure_return_tag :  in   std_logic_vector(0 downto 0);
    sendOutput_call_reqs : out  std_logic_vector(0 downto 0);
    sendOutput_call_acks : in   std_logic_vector(0 downto 0);
    sendOutput_call_tag  :  out  std_logic_vector(0 downto 0);
    sendOutput_return_reqs : out  std_logic_vector(0 downto 0);
    sendOutput_return_acks : in   std_logic_vector(0 downto 0);
    sendOutput_return_tag :  in   std_logic_vector(0 downto 0);
    timer_call_reqs : out  std_logic_vector(0 downto 0);
    timer_call_acks : in   std_logic_vector(0 downto 0);
    timer_call_tag  :  out  std_logic_vector(1 downto 0);
    timer_return_reqs : out  std_logic_vector(0 downto 0);
    timer_return_acks : in   std_logic_vector(0 downto 0);
    timer_return_data : in   std_logic_vector(31 downto 0);
    timer_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTranspose;
architecture convTranspose_arch of convTranspose is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTranspose_CP_3766_start: Boolean;
  signal convTranspose_CP_3766_symbol: Boolean;
  -- volatile/operator module components. 
  component testConfigure is -- 
    generic (tag_length : integer); 
    port ( -- 
      ret_val_x_x : out  std_logic_vector(15 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sr_addr : out  std_logic_vector(10 downto 0);
      memory_space_5_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_5_sr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_6_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_6_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_7_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_7_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_7_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_8_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_8_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_8_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_8_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_8_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_8_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_4_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_4_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sc_tag :  in  std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component sendOutput is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_6_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_6_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(2 downto 0);
      ConvTranspose_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      c : out  std_logic_vector(31 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal WPIPE_Block3_start_1340_inst_req_0 : boolean;
  signal RPIPE_Block1_done_1348_inst_ack_1 : boolean;
  signal call_stmt_1358_call_ack_0 : boolean;
  signal RPIPE_Block1_done_1348_inst_req_0 : boolean;
  signal call_stmt_1358_call_ack_1 : boolean;
  signal call_stmt_1358_call_req_1 : boolean;
  signal WPIPE_Block2_start_1336_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1336_inst_req_0 : boolean;
  signal RPIPE_Block1_done_1348_inst_ack_0 : boolean;
  signal RPIPE_Block3_done_1354_inst_ack_1 : boolean;
  signal RPIPE_Block3_done_1354_inst_req_1 : boolean;
  signal RPIPE_Block1_done_1348_inst_req_1 : boolean;
  signal RPIPE_Block2_done_1351_inst_req_0 : boolean;
  signal WPIPE_elapsed_time_pipe_1368_inst_req_1 : boolean;
  signal RPIPE_Block0_done_1345_inst_req_1 : boolean;
  signal RPIPE_Block2_done_1351_inst_ack_0 : boolean;
  signal call_stmt_1358_call_req_0 : boolean;
  signal WPIPE_Block2_start_1336_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1336_inst_req_1 : boolean;
  signal WPIPE_Block3_start_1340_inst_ack_0 : boolean;
  signal call_stmt_1327_call_req_0 : boolean;
  signal call_stmt_1327_call_ack_0 : boolean;
  signal type_cast_1366_inst_ack_1 : boolean;
  signal type_cast_1366_inst_req_1 : boolean;
  signal type_cast_1366_inst_ack_0 : boolean;
  signal type_cast_1366_inst_req_0 : boolean;
  signal RPIPE_Block2_done_1351_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1332_inst_ack_1 : boolean;
  signal RPIPE_Block0_done_1345_inst_ack_0 : boolean;
  signal RPIPE_Block0_done_1345_inst_req_0 : boolean;
  signal WPIPE_elapsed_time_pipe_1368_inst_ack_1 : boolean;
  signal call_stmt_1324_call_ack_1 : boolean;
  signal call_stmt_1324_call_req_1 : boolean;
  signal WPIPE_Block1_start_1332_inst_req_1 : boolean;
  signal RPIPE_Block3_done_1354_inst_ack_0 : boolean;
  signal call_stmt_1327_call_ack_1 : boolean;
  signal WPIPE_elapsed_time_pipe_1368_inst_ack_0 : boolean;
  signal WPIPE_Block1_start_1332_inst_ack_0 : boolean;
  signal RPIPE_Block2_done_1351_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1332_inst_req_0 : boolean;
  signal RPIPE_Block3_done_1354_inst_req_0 : boolean;
  signal call_stmt_1324_call_ack_0 : boolean;
  signal call_stmt_1327_call_req_1 : boolean;
  signal RPIPE_Block0_done_1345_inst_ack_1 : boolean;
  signal call_stmt_1324_call_req_0 : boolean;
  signal call_stmt_1371_call_ack_1 : boolean;
  signal call_stmt_1371_call_req_1 : boolean;
  signal WPIPE_elapsed_time_pipe_1368_inst_req_0 : boolean;
  signal WPIPE_Block0_start_1328_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1328_inst_req_1 : boolean;
  signal call_stmt_1371_call_ack_0 : boolean;
  signal call_stmt_1371_call_req_0 : boolean;
  signal WPIPE_Block0_start_1328_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_1328_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1340_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1340_inst_req_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTranspose_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTranspose_CP_3766_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTranspose_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTranspose_CP_3766_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTranspose_CP_3766_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTranspose_CP_3766_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTranspose_CP_3766: Block -- control-path 
    signal convTranspose_CP_3766_elements: BooleanArray(30 downto 0);
    -- 
  begin -- 
    convTranspose_CP_3766_elements(0) <= convTranspose_CP_3766_start;
    convTranspose_CP_3766_symbol <= convTranspose_CP_3766_elements(30);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (11) 
      -- CP-element group 0: 	 branch_block_stmt_1322/call_stmt_1324__entry__
      -- CP-element group 0: 	 branch_block_stmt_1322/call_stmt_1324/call_stmt_1324_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1322/call_stmt_1324/call_stmt_1324_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1322/call_stmt_1324/call_stmt_1324_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1322/call_stmt_1324/$entry
      -- CP-element group 0: 	 branch_block_stmt_1322/$entry
      -- CP-element group 0: 	 branch_block_stmt_1322/call_stmt_1324/call_stmt_1324_Update/ccr
      -- CP-element group 0: 	 branch_block_stmt_1322/call_stmt_1324/call_stmt_1324_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1322/call_stmt_1324/call_stmt_1324_Sample/crr
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1322/branch_block_stmt_1322__entry__
      -- 
    ccr_3797_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3797_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3766_elements(0), ack => call_stmt_1324_call_req_1); -- 
    crr_3792_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3792_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3766_elements(0), ack => call_stmt_1324_call_req_0); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 branch_block_stmt_1322/call_stmt_1324/call_stmt_1324_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_1322/call_stmt_1324/call_stmt_1324_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_1322/call_stmt_1324/call_stmt_1324_Sample/cra
      -- 
    cra_3793_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1324_call_ack_0, ack => convTranspose_CP_3766_elements(1)); -- 
    -- CP-element group 2:  fork  transition  place  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	5 
    -- CP-element group 2: 	7 
    -- CP-element group 2: 	4 
    -- CP-element group 2: 	9 
    -- CP-element group 2: 	13 
    -- CP-element group 2: 	19 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	15 
    -- CP-element group 2: 	11 
    -- CP-element group 2: 	17 
    -- CP-element group 2:  members (37) 
      -- CP-element group 2: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/WPIPE_Block3_start_1340_Sample/req
      -- CP-element group 2: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/RPIPE_Block1_done_1348_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/WPIPE_Block2_start_1336_Sample/req
      -- CP-element group 2: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/WPIPE_Block3_start_1340_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/WPIPE_Block2_start_1336_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/RPIPE_Block1_done_1348_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355__entry__
      -- CP-element group 2: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/call_stmt_1327_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/WPIPE_Block3_start_1340_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/RPIPE_Block2_done_1351_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/RPIPE_Block2_done_1351_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/call_stmt_1327_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/call_stmt_1327_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/call_stmt_1327_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1322/call_stmt_1324__exit__
      -- CP-element group 2: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/call_stmt_1327_Sample/crr
      -- CP-element group 2: 	 branch_block_stmt_1322/call_stmt_1324/call_stmt_1324_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/$entry
      -- CP-element group 2: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/WPIPE_Block2_start_1336_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1322/call_stmt_1324/$exit
      -- CP-element group 2: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/RPIPE_Block0_done_1345_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_1322/call_stmt_1324/call_stmt_1324_Update/cca
      -- CP-element group 2: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/WPIPE_Block0_start_1328_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/RPIPE_Block2_done_1351_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/RPIPE_Block1_done_1348_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1322/call_stmt_1324/call_stmt_1324_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/RPIPE_Block0_done_1345_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/WPIPE_Block1_start_1332_Sample/req
      -- CP-element group 2: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/RPIPE_Block3_done_1354_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/call_stmt_1327_Update/ccr
      -- CP-element group 2: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/RPIPE_Block3_done_1354_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/WPIPE_Block1_start_1332_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/WPIPE_Block1_start_1332_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/RPIPE_Block3_done_1354_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/RPIPE_Block0_done_1345_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/WPIPE_Block0_start_1328_Sample/req
      -- CP-element group 2: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/WPIPE_Block0_start_1328_Sample/$entry
      -- 
    cca_3798_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1324_call_ack_1, ack => convTranspose_CP_3766_elements(2)); -- 
    req_3865_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3865_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3766_elements(2), ack => WPIPE_Block3_start_1340_inst_req_0); -- 
    rr_3893_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3893_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3766_elements(2), ack => RPIPE_Block1_done_1348_inst_req_0); -- 
    req_3851_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3851_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3766_elements(2), ack => WPIPE_Block2_start_1336_inst_req_0); -- 
    rr_3907_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3907_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3766_elements(2), ack => RPIPE_Block2_done_1351_inst_req_0); -- 
    crr_3809_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3809_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3766_elements(2), ack => call_stmt_1327_call_req_0); -- 
    rr_3879_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3879_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3766_elements(2), ack => RPIPE_Block0_done_1345_inst_req_0); -- 
    req_3837_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3837_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3766_elements(2), ack => WPIPE_Block1_start_1332_inst_req_0); -- 
    rr_3921_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3921_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3766_elements(2), ack => RPIPE_Block3_done_1354_inst_req_0); -- 
    ccr_3814_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3814_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3766_elements(2), ack => call_stmt_1327_call_req_1); -- 
    req_3823_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3823_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3766_elements(2), ack => WPIPE_Block0_start_1328_inst_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/call_stmt_1327_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/call_stmt_1327_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/call_stmt_1327_Sample/cra
      -- 
    cra_3810_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1327_call_ack_0, ack => convTranspose_CP_3766_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	2 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	21 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/call_stmt_1327_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/call_stmt_1327_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/call_stmt_1327_Update/cca
      -- 
    cca_3815_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1327_call_ack_1, ack => convTranspose_CP_3766_elements(4)); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/WPIPE_Block0_start_1328_update_start_
      -- CP-element group 5: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/WPIPE_Block0_start_1328_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/WPIPE_Block0_start_1328_Update/req
      -- CP-element group 5: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/WPIPE_Block0_start_1328_Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/WPIPE_Block0_start_1328_Sample/ack
      -- CP-element group 5: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/WPIPE_Block0_start_1328_Sample/$exit
      -- 
    ack_3824_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1328_inst_ack_0, ack => convTranspose_CP_3766_elements(5)); -- 
    req_3828_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3828_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3766_elements(5), ack => WPIPE_Block0_start_1328_inst_req_1); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	21 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/WPIPE_Block0_start_1328_Update/ack
      -- CP-element group 6: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/WPIPE_Block0_start_1328_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/WPIPE_Block0_start_1328_update_completed_
      -- 
    ack_3829_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1328_inst_ack_1, ack => convTranspose_CP_3766_elements(6)); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	2 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/WPIPE_Block1_start_1332_Update/req
      -- CP-element group 7: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/WPIPE_Block1_start_1332_Update/$entry
      -- CP-element group 7: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/WPIPE_Block1_start_1332_Sample/ack
      -- CP-element group 7: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/WPIPE_Block1_start_1332_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/WPIPE_Block1_start_1332_update_start_
      -- CP-element group 7: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/WPIPE_Block1_start_1332_sample_completed_
      -- 
    ack_3838_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1332_inst_ack_0, ack => convTranspose_CP_3766_elements(7)); -- 
    req_3842_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3842_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3766_elements(7), ack => WPIPE_Block1_start_1332_inst_req_1); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	21 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/WPIPE_Block1_start_1332_Update/ack
      -- CP-element group 8: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/WPIPE_Block1_start_1332_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/WPIPE_Block1_start_1332_update_completed_
      -- 
    ack_3843_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1332_inst_ack_1, ack => convTranspose_CP_3766_elements(8)); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	2 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/WPIPE_Block2_start_1336_Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/WPIPE_Block2_start_1336_Sample/ack
      -- CP-element group 9: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/WPIPE_Block2_start_1336_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/WPIPE_Block2_start_1336_Update/req
      -- CP-element group 9: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/WPIPE_Block2_start_1336_update_start_
      -- CP-element group 9: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/WPIPE_Block2_start_1336_sample_completed_
      -- 
    ack_3852_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1336_inst_ack_0, ack => convTranspose_CP_3766_elements(9)); -- 
    req_3856_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3856_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3766_elements(9), ack => WPIPE_Block2_start_1336_inst_req_1); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	21 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/WPIPE_Block2_start_1336_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/WPIPE_Block2_start_1336_Update/ack
      -- CP-element group 10: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/WPIPE_Block2_start_1336_Update/$exit
      -- 
    ack_3857_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1336_inst_ack_1, ack => convTranspose_CP_3766_elements(10)); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	2 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/WPIPE_Block3_start_1340_update_start_
      -- CP-element group 11: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/WPIPE_Block3_start_1340_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/WPIPE_Block3_start_1340_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/WPIPE_Block3_start_1340_Sample/ack
      -- CP-element group 11: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/WPIPE_Block3_start_1340_Update/$entry
      -- CP-element group 11: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/WPIPE_Block3_start_1340_Update/req
      -- 
    ack_3866_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1340_inst_ack_0, ack => convTranspose_CP_3766_elements(11)); -- 
    req_3870_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3870_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3766_elements(11), ack => WPIPE_Block3_start_1340_inst_req_1); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	21 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/WPIPE_Block3_start_1340_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/WPIPE_Block3_start_1340_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/WPIPE_Block3_start_1340_Update/ack
      -- 
    ack_3871_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1340_inst_ack_1, ack => convTranspose_CP_3766_elements(12)); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	2 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/RPIPE_Block0_done_1345_Update/cr
      -- CP-element group 13: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/RPIPE_Block0_done_1345_Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/RPIPE_Block0_done_1345_Sample/ra
      -- CP-element group 13: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/RPIPE_Block0_done_1345_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/RPIPE_Block0_done_1345_update_start_
      -- CP-element group 13: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/RPIPE_Block0_done_1345_sample_completed_
      -- 
    ra_3880_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_done_1345_inst_ack_0, ack => convTranspose_CP_3766_elements(13)); -- 
    cr_3884_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3884_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3766_elements(13), ack => RPIPE_Block0_done_1345_inst_req_1); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	21 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/RPIPE_Block0_done_1345_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/RPIPE_Block0_done_1345_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/RPIPE_Block0_done_1345_Update/ca
      -- 
    ca_3885_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_done_1345_inst_ack_1, ack => convTranspose_CP_3766_elements(14)); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	2 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/RPIPE_Block1_done_1348_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/RPIPE_Block1_done_1348_Sample/ra
      -- CP-element group 15: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/RPIPE_Block1_done_1348_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/RPIPE_Block1_done_1348_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/RPIPE_Block1_done_1348_update_start_
      -- CP-element group 15: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/RPIPE_Block1_done_1348_sample_completed_
      -- 
    ra_3894_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_done_1348_inst_ack_0, ack => convTranspose_CP_3766_elements(15)); -- 
    cr_3898_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3898_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3766_elements(15), ack => RPIPE_Block1_done_1348_inst_req_1); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	21 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/RPIPE_Block1_done_1348_Update/ca
      -- CP-element group 16: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/RPIPE_Block1_done_1348_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/RPIPE_Block1_done_1348_update_completed_
      -- 
    ca_3899_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_done_1348_inst_ack_1, ack => convTranspose_CP_3766_elements(16)); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	2 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/RPIPE_Block2_done_1351_update_start_
      -- CP-element group 17: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/RPIPE_Block2_done_1351_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/RPIPE_Block2_done_1351_Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/RPIPE_Block2_done_1351_Update/cr
      -- CP-element group 17: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/RPIPE_Block2_done_1351_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/RPIPE_Block2_done_1351_Update/$entry
      -- 
    ra_3908_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_done_1351_inst_ack_0, ack => convTranspose_CP_3766_elements(17)); -- 
    cr_3912_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3912_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3766_elements(17), ack => RPIPE_Block2_done_1351_inst_req_1); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	21 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/RPIPE_Block2_done_1351_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/RPIPE_Block2_done_1351_Update/ca
      -- CP-element group 18: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/RPIPE_Block2_done_1351_Update/$exit
      -- 
    ca_3913_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_done_1351_inst_ack_1, ack => convTranspose_CP_3766_elements(18)); -- 
    -- CP-element group 19:  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	2 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (6) 
      -- CP-element group 19: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/RPIPE_Block3_done_1354_Update/cr
      -- CP-element group 19: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/RPIPE_Block3_done_1354_Update/$entry
      -- CP-element group 19: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/RPIPE_Block3_done_1354_Sample/ra
      -- CP-element group 19: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/RPIPE_Block3_done_1354_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/RPIPE_Block3_done_1354_update_start_
      -- CP-element group 19: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/RPIPE_Block3_done_1354_sample_completed_
      -- 
    ra_3922_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_done_1354_inst_ack_0, ack => convTranspose_CP_3766_elements(19)); -- 
    cr_3926_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3926_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3766_elements(19), ack => RPIPE_Block3_done_1354_inst_req_1); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/RPIPE_Block3_done_1354_Update/ca
      -- CP-element group 20: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/RPIPE_Block3_done_1354_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/RPIPE_Block3_done_1354_update_completed_
      -- 
    ca_3927_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_done_1354_inst_ack_1, ack => convTranspose_CP_3766_elements(20)); -- 
    -- CP-element group 21:  join  fork  transition  place  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	6 
    -- CP-element group 21: 	4 
    -- CP-element group 21: 	8 
    -- CP-element group 21: 	20 
    -- CP-element group 21: 	14 
    -- CP-element group 21: 	10 
    -- CP-element group 21: 	18 
    -- CP-element group 21: 	12 
    -- CP-element group 21: 	16 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	23 
    -- CP-element group 21: 	25 
    -- CP-element group 21: 	28 
    -- CP-element group 21: 	29 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (19) 
      -- CP-element group 21: 	 branch_block_stmt_1322/call_stmt_1358_to_call_stmt_1371/call_stmt_1358_Update/$entry
      -- CP-element group 21: 	 branch_block_stmt_1322/call_stmt_1358_to_call_stmt_1371/call_stmt_1358_Update/ccr
      -- CP-element group 21: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355/$exit
      -- CP-element group 21: 	 branch_block_stmt_1322/call_stmt_1327_to_assign_stmt_1355__exit__
      -- CP-element group 21: 	 branch_block_stmt_1322/call_stmt_1358_to_call_stmt_1371/call_stmt_1358_Sample/crr
      -- CP-element group 21: 	 branch_block_stmt_1322/call_stmt_1358_to_call_stmt_1371/call_stmt_1358_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_1322/call_stmt_1358_to_call_stmt_1371/type_cast_1366_update_start_
      -- CP-element group 21: 	 branch_block_stmt_1322/call_stmt_1358_to_call_stmt_1371__entry__
      -- CP-element group 21: 	 branch_block_stmt_1322/call_stmt_1358_to_call_stmt_1371/call_stmt_1371_update_start_
      -- CP-element group 21: 	 branch_block_stmt_1322/call_stmt_1358_to_call_stmt_1371/type_cast_1366_Update/cr
      -- CP-element group 21: 	 branch_block_stmt_1322/call_stmt_1358_to_call_stmt_1371/type_cast_1366_Update/$entry
      -- CP-element group 21: 	 branch_block_stmt_1322/call_stmt_1358_to_call_stmt_1371/call_stmt_1358_update_start_
      -- CP-element group 21: 	 branch_block_stmt_1322/call_stmt_1358_to_call_stmt_1371/call_stmt_1358_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_1322/call_stmt_1358_to_call_stmt_1371/$entry
      -- CP-element group 21: 	 branch_block_stmt_1322/call_stmt_1358_to_call_stmt_1371/call_stmt_1371_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_1322/call_stmt_1358_to_call_stmt_1371/call_stmt_1371_Update/ccr
      -- CP-element group 21: 	 branch_block_stmt_1322/call_stmt_1358_to_call_stmt_1371/call_stmt_1371_Update/$entry
      -- CP-element group 21: 	 branch_block_stmt_1322/call_stmt_1358_to_call_stmt_1371/call_stmt_1371_Sample/crr
      -- CP-element group 21: 	 branch_block_stmt_1322/call_stmt_1358_to_call_stmt_1371/call_stmt_1371_Sample/$entry
      -- 
    ccr_3943_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3943_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3766_elements(21), ack => call_stmt_1358_call_req_1); -- 
    crr_3938_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3938_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3766_elements(21), ack => call_stmt_1358_call_req_0); -- 
    cr_3957_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3957_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3766_elements(21), ack => type_cast_1366_inst_req_1); -- 
    ccr_3985_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3985_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3766_elements(21), ack => call_stmt_1371_call_req_1); -- 
    crr_3980_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3980_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3766_elements(21), ack => call_stmt_1371_call_req_0); -- 
    convTranspose_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convTranspose_CP_3766_elements(6) & convTranspose_CP_3766_elements(4) & convTranspose_CP_3766_elements(8) & convTranspose_CP_3766_elements(20) & convTranspose_CP_3766_elements(14) & convTranspose_CP_3766_elements(10) & convTranspose_CP_3766_elements(18) & convTranspose_CP_3766_elements(12) & convTranspose_CP_3766_elements(16);
      gj_convTranspose_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_3766_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_1322/call_stmt_1358_to_call_stmt_1371/call_stmt_1358_Sample/cra
      -- CP-element group 22: 	 branch_block_stmt_1322/call_stmt_1358_to_call_stmt_1371/call_stmt_1358_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_1322/call_stmt_1358_to_call_stmt_1371/call_stmt_1358_sample_completed_
      -- 
    cra_3939_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1358_call_ack_0, ack => convTranspose_CP_3766_elements(22)); -- 
    -- CP-element group 23:  transition  input  output  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	21 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23:  members (6) 
      -- CP-element group 23: 	 branch_block_stmt_1322/call_stmt_1358_to_call_stmt_1371/call_stmt_1358_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_1322/call_stmt_1358_to_call_stmt_1371/call_stmt_1358_Update/cca
      -- CP-element group 23: 	 branch_block_stmt_1322/call_stmt_1358_to_call_stmt_1371/type_cast_1366_sample_start_
      -- CP-element group 23: 	 branch_block_stmt_1322/call_stmt_1358_to_call_stmt_1371/type_cast_1366_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_1322/call_stmt_1358_to_call_stmt_1371/call_stmt_1358_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_1322/call_stmt_1358_to_call_stmt_1371/type_cast_1366_Sample/rr
      -- 
    cca_3944_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1358_call_ack_1, ack => convTranspose_CP_3766_elements(23)); -- 
    rr_3952_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3952_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3766_elements(23), ack => type_cast_1366_inst_req_0); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_1322/call_stmt_1358_to_call_stmt_1371/type_cast_1366_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_1322/call_stmt_1358_to_call_stmt_1371/type_cast_1366_Sample/ra
      -- CP-element group 24: 	 branch_block_stmt_1322/call_stmt_1358_to_call_stmt_1371/type_cast_1366_Sample/$exit
      -- 
    ra_3953_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1366_inst_ack_0, ack => convTranspose_CP_3766_elements(24)); -- 
    -- CP-element group 25:  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	21 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25:  members (6) 
      -- CP-element group 25: 	 branch_block_stmt_1322/call_stmt_1358_to_call_stmt_1371/WPIPE_elapsed_time_pipe_1368_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_1322/call_stmt_1358_to_call_stmt_1371/type_cast_1366_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_1322/call_stmt_1358_to_call_stmt_1371/type_cast_1366_Update/ca
      -- CP-element group 25: 	 branch_block_stmt_1322/call_stmt_1358_to_call_stmt_1371/type_cast_1366_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_1322/call_stmt_1358_to_call_stmt_1371/WPIPE_elapsed_time_pipe_1368_Sample/req
      -- CP-element group 25: 	 branch_block_stmt_1322/call_stmt_1358_to_call_stmt_1371/WPIPE_elapsed_time_pipe_1368_Sample/$entry
      -- 
    ca_3958_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1366_inst_ack_1, ack => convTranspose_CP_3766_elements(25)); -- 
    req_3966_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3966_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3766_elements(25), ack => WPIPE_elapsed_time_pipe_1368_inst_req_0); -- 
    -- CP-element group 26:  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (6) 
      -- CP-element group 26: 	 branch_block_stmt_1322/call_stmt_1358_to_call_stmt_1371/WPIPE_elapsed_time_pipe_1368_update_start_
      -- CP-element group 26: 	 branch_block_stmt_1322/call_stmt_1358_to_call_stmt_1371/WPIPE_elapsed_time_pipe_1368_Update/req
      -- CP-element group 26: 	 branch_block_stmt_1322/call_stmt_1358_to_call_stmt_1371/WPIPE_elapsed_time_pipe_1368_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_1322/call_stmt_1358_to_call_stmt_1371/WPIPE_elapsed_time_pipe_1368_Sample/ack
      -- CP-element group 26: 	 branch_block_stmt_1322/call_stmt_1358_to_call_stmt_1371/WPIPE_elapsed_time_pipe_1368_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_1322/call_stmt_1358_to_call_stmt_1371/WPIPE_elapsed_time_pipe_1368_Update/$entry
      -- 
    ack_3967_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_elapsed_time_pipe_1368_inst_ack_0, ack => convTranspose_CP_3766_elements(26)); -- 
    req_3971_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3971_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3766_elements(26), ack => WPIPE_elapsed_time_pipe_1368_inst_req_1); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	30 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1322/call_stmt_1358_to_call_stmt_1371/WPIPE_elapsed_time_pipe_1368_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_1322/call_stmt_1358_to_call_stmt_1371/WPIPE_elapsed_time_pipe_1368_Update/ack
      -- CP-element group 27: 	 branch_block_stmt_1322/call_stmt_1358_to_call_stmt_1371/WPIPE_elapsed_time_pipe_1368_Update/$exit
      -- 
    ack_3972_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_elapsed_time_pipe_1368_inst_ack_1, ack => convTranspose_CP_3766_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	21 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_1322/call_stmt_1358_to_call_stmt_1371/call_stmt_1371_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_1322/call_stmt_1358_to_call_stmt_1371/call_stmt_1371_Sample/cra
      -- CP-element group 28: 	 branch_block_stmt_1322/call_stmt_1358_to_call_stmt_1371/call_stmt_1371_Sample/$exit
      -- 
    cra_3981_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1371_call_ack_0, ack => convTranspose_CP_3766_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	21 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_1322/call_stmt_1358_to_call_stmt_1371/call_stmt_1371_Update/cca
      -- CP-element group 29: 	 branch_block_stmt_1322/call_stmt_1358_to_call_stmt_1371/call_stmt_1371_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_1322/call_stmt_1358_to_call_stmt_1371/call_stmt_1371_update_completed_
      -- 
    cca_3986_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1371_call_ack_1, ack => convTranspose_CP_3766_elements(29)); -- 
    -- CP-element group 30:  join  transition  place  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	27 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (13) 
      -- CP-element group 30: 	 branch_block_stmt_1322/branch_block_stmt_1322__exit__
      -- CP-element group 30: 	 branch_block_stmt_1322/$exit
      -- CP-element group 30: 	 branch_block_stmt_1322/merge_stmt_1373_PhiReqMerge
      -- CP-element group 30: 	 branch_block_stmt_1322/merge_stmt_1373__exit__
      -- CP-element group 30: 	 branch_block_stmt_1322/return__
      -- CP-element group 30: 	 $exit
      -- CP-element group 30: 	 branch_block_stmt_1322/call_stmt_1358_to_call_stmt_1371__exit__
      -- CP-element group 30: 	 branch_block_stmt_1322/call_stmt_1358_to_call_stmt_1371/$exit
      -- CP-element group 30: 	 branch_block_stmt_1322/merge_stmt_1373_PhiAck/dummy
      -- CP-element group 30: 	 branch_block_stmt_1322/merge_stmt_1373_PhiAck/$entry
      -- CP-element group 30: 	 branch_block_stmt_1322/merge_stmt_1373_PhiAck/$exit
      -- CP-element group 30: 	 branch_block_stmt_1322/return___PhiReq/$entry
      -- CP-element group 30: 	 branch_block_stmt_1322/return___PhiReq/$exit
      -- 
    convTranspose_cp_element_group_30: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_30"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTranspose_CP_3766_elements(27) & convTranspose_CP_3766_elements(29);
      gj_convTranspose_cp_element_group_30 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_3766_elements(30), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal call10_1352 : std_logic_vector(15 downto 0);
    signal call12_1355 : std_logic_vector(15 downto 0);
    signal call14_1358 : std_logic_vector(31 downto 0);
    signal call1_1327 : std_logic_vector(31 downto 0);
    signal call6_1346 : std_logic_vector(15 downto 0);
    signal call8_1349 : std_logic_vector(15 downto 0);
    signal call_1324 : std_logic_vector(15 downto 0);
    signal conv_1367 : std_logic_vector(63 downto 0);
    signal sub_1363 : std_logic_vector(31 downto 0);
    signal type_cast_1330_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1334_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1338_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1342_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    type_cast_1330_wire_constant <= "0000000000000001";
    type_cast_1334_wire_constant <= "0000000000000001";
    type_cast_1338_wire_constant <= "0000000000000001";
    type_cast_1342_wire_constant <= "0000000000000001";
    type_cast_1366_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1366_inst_req_0;
      type_cast_1366_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1366_inst_req_1;
      type_cast_1366_inst_ack_1<= rack(0);
      type_cast_1366_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1366_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub_1363,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_1367,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- binary operator SUB_u32_u32_1362_inst
    process(call14_1358, call1_1327) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(call14_1358, call1_1327, tmp_var);
      sub_1363 <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_Block0_done_1345_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block0_done_1345_inst_req_0;
      RPIPE_Block0_done_1345_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block0_done_1345_inst_req_1;
      RPIPE_Block0_done_1345_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call6_1346 <= data_out(15 downto 0);
      Block0_done_read_0_gI: SplitGuardInterface generic map(name => "Block0_done_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block0_done_read_0: InputPortRevised -- 
        generic map ( name => "Block0_done_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block0_done_pipe_read_req(0),
          oack => Block0_done_pipe_read_ack(0),
          odata => Block0_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_Block1_done_1348_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block1_done_1348_inst_req_0;
      RPIPE_Block1_done_1348_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block1_done_1348_inst_req_1;
      RPIPE_Block1_done_1348_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call8_1349 <= data_out(15 downto 0);
      Block1_done_read_1_gI: SplitGuardInterface generic map(name => "Block1_done_read_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block1_done_read_1: InputPortRevised -- 
        generic map ( name => "Block1_done_read_1", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block1_done_pipe_read_req(0),
          oack => Block1_done_pipe_read_ack(0),
          odata => Block1_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : RPIPE_Block2_done_1351_inst 
    InportGroup_2: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block2_done_1351_inst_req_0;
      RPIPE_Block2_done_1351_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block2_done_1351_inst_req_1;
      RPIPE_Block2_done_1351_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call10_1352 <= data_out(15 downto 0);
      Block2_done_read_2_gI: SplitGuardInterface generic map(name => "Block2_done_read_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block2_done_read_2: InputPortRevised -- 
        generic map ( name => "Block2_done_read_2", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block2_done_pipe_read_req(0),
          oack => Block2_done_pipe_read_ack(0),
          odata => Block2_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : RPIPE_Block3_done_1354_inst 
    InportGroup_3: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block3_done_1354_inst_req_0;
      RPIPE_Block3_done_1354_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block3_done_1354_inst_req_1;
      RPIPE_Block3_done_1354_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call12_1355 <= data_out(15 downto 0);
      Block3_done_read_3_gI: SplitGuardInterface generic map(name => "Block3_done_read_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block3_done_read_3: InputPortRevised -- 
        generic map ( name => "Block3_done_read_3", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block3_done_pipe_read_req(0),
          oack => Block3_done_pipe_read_ack(0),
          odata => Block3_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- shared outport operator group (0) : WPIPE_Block0_start_1328_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block0_start_1328_inst_req_0;
      WPIPE_Block0_start_1328_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block0_start_1328_inst_req_1;
      WPIPE_Block0_start_1328_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_1330_wire_constant;
      Block0_start_write_0_gI: SplitGuardInterface generic map(name => "Block0_start_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block0_start_write_0: OutputPortRevised -- 
        generic map ( name => "Block0_start", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block0_start_pipe_write_req(0),
          oack => Block0_start_pipe_write_ack(0),
          odata => Block0_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_Block1_start_1332_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block1_start_1332_inst_req_0;
      WPIPE_Block1_start_1332_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block1_start_1332_inst_req_1;
      WPIPE_Block1_start_1332_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_1334_wire_constant;
      Block1_start_write_1_gI: SplitGuardInterface generic map(name => "Block1_start_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block1_start_write_1: OutputPortRevised -- 
        generic map ( name => "Block1_start", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block1_start_pipe_write_req(0),
          oack => Block1_start_pipe_write_ack(0),
          odata => Block1_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_Block2_start_1336_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block2_start_1336_inst_req_0;
      WPIPE_Block2_start_1336_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block2_start_1336_inst_req_1;
      WPIPE_Block2_start_1336_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_1338_wire_constant;
      Block2_start_write_2_gI: SplitGuardInterface generic map(name => "Block2_start_write_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block2_start_write_2: OutputPortRevised -- 
        generic map ( name => "Block2_start", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block2_start_pipe_write_req(0),
          oack => Block2_start_pipe_write_ack(0),
          odata => Block2_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_Block3_start_1340_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block3_start_1340_inst_req_0;
      WPIPE_Block3_start_1340_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block3_start_1340_inst_req_1;
      WPIPE_Block3_start_1340_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_1342_wire_constant;
      Block3_start_write_3_gI: SplitGuardInterface generic map(name => "Block3_start_write_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block3_start_write_3: OutputPortRevised -- 
        generic map ( name => "Block3_start", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block3_start_pipe_write_req(0),
          oack => Block3_start_pipe_write_ack(0),
          odata => Block3_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- shared outport operator group (4) : WPIPE_elapsed_time_pipe_1368_inst 
    OutportGroup_4: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_elapsed_time_pipe_1368_inst_req_0;
      WPIPE_elapsed_time_pipe_1368_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_elapsed_time_pipe_1368_inst_req_1;
      WPIPE_elapsed_time_pipe_1368_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= conv_1367;
      elapsed_time_pipe_write_4_gI: SplitGuardInterface generic map(name => "elapsed_time_pipe_write_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      elapsed_time_pipe_write_4: OutputPortRevised -- 
        generic map ( name => "elapsed_time_pipe", data_width => 64, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => elapsed_time_pipe_pipe_write_req(0),
          oack => elapsed_time_pipe_pipe_write_ack(0),
          odata => elapsed_time_pipe_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 4
    -- shared call operator group (0) : call_stmt_1324_call 
    testConfigure_call_group_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1324_call_req_0;
      call_stmt_1324_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1324_call_req_1;
      call_stmt_1324_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      testConfigure_call_group_0_gI: SplitGuardInterface generic map(name => "testConfigure_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      call_1324 <= data_out(15 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 1,
        nreqs => 1,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => testConfigure_call_reqs(0),
          ackR => testConfigure_call_acks(0),
          tagR => testConfigure_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 16,
          owidth => 16,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => testConfigure_return_acks(0), -- cross-over
          ackL => testConfigure_return_reqs(0), -- cross-over
          dataL => testConfigure_return_data(15 downto 0),
          tagL => testConfigure_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_1358_call call_stmt_1327_call 
    timer_call_group_1: Block -- 
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_1358_call_req_0;
      reqL_unguarded(0) <= call_stmt_1327_call_req_0;
      call_stmt_1358_call_ack_0 <= ackL_unguarded(1);
      call_stmt_1327_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_1358_call_req_1;
      reqR_unguarded(0) <= call_stmt_1327_call_req_1;
      call_stmt_1358_call_ack_1 <= ackR_unguarded(1);
      call_stmt_1327_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      timer_call_group_1_accessRegulator_0: access_regulator_base generic map (name => "timer_call_group_1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      timer_call_group_1_accessRegulator_1: access_regulator_base generic map (name => "timer_call_group_1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      timer_call_group_1_gI: SplitGuardInterface generic map(name => "timer_call_group_1_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      call14_1358 <= data_out(63 downto 32);
      call1_1327 <= data_out(31 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 2,
        nreqs => 2,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => timer_call_reqs(0),
          ackR => timer_call_acks(0),
          tagR => timer_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => timer_return_acks(0), -- cross-over
          ackL => timer_return_reqs(0), -- cross-over
          dataL => timer_return_data(31 downto 0),
          tagL => timer_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- shared call operator group (2) : call_stmt_1371_call 
    sendOutput_call_group_2: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1371_call_req_0;
      call_stmt_1371_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1371_call_req_1;
      call_stmt_1371_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      sendOutput_call_group_2_gI: SplitGuardInterface generic map(name => "sendOutput_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 1,
        nreqs => 1,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => sendOutput_call_reqs(0),
          ackR => sendOutput_call_acks(0),
          tagR => sendOutput_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => sendOutput_return_acks(0), -- cross-over
          ackL => sendOutput_return_reqs(0), -- cross-over
          tagL => sendOutput_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- 
  end Block; -- data_path
  -- 
end convTranspose_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeA is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_7_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_8_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_8_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_8_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_8_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_8_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_8_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_4_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_4_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_6_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_6_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_sc_tag :  in  std_logic_vector(0 downto 0);
    Block0_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block0_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block0_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block0_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block0_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block0_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeA;
architecture convTransposeA_arch of convTransposeA is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeA_CP_3995_start: Boolean;
  signal convTransposeA_CP_3995_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal ptr_deref_1505_load_0_ack_1 : boolean;
  signal array_obj_ref_1729_index_offset_req_1 : boolean;
  signal array_obj_ref_1698_index_offset_ack_0 : boolean;
  signal ptr_deref_1703_load_0_req_1 : boolean;
  signal array_obj_ref_1729_index_offset_ack_1 : boolean;
  signal ptr_deref_1703_load_0_ack_1 : boolean;
  signal ptr_deref_1733_store_0_ack_1 : boolean;
  signal type_cast_1739_inst_ack_0 : boolean;
  signal if_stmt_1752_branch_req_0 : boolean;
  signal addr_of_1730_final_reg_ack_0 : boolean;
  signal type_cast_1739_inst_req_0 : boolean;
  signal type_cast_1739_inst_req_1 : boolean;
  signal addr_of_1730_final_reg_req_0 : boolean;
  signal ptr_deref_1733_store_0_ack_0 : boolean;
  signal ptr_deref_1733_store_0_req_1 : boolean;
  signal type_cast_1723_inst_req_0 : boolean;
  signal array_obj_ref_1698_index_offset_req_0 : boolean;
  signal array_obj_ref_1698_index_offset_ack_1 : boolean;
  signal array_obj_ref_1729_index_offset_req_0 : boolean;
  signal ptr_deref_1505_load_0_req_1 : boolean;
  signal array_obj_ref_1729_index_offset_ack_0 : boolean;
  signal type_cast_1739_inst_ack_1 : boolean;
  signal type_cast_1723_inst_ack_0 : boolean;
  signal addr_of_1730_final_reg_req_1 : boolean;
  signal addr_of_1730_final_reg_ack_1 : boolean;
  signal ptr_deref_1733_store_0_req_0 : boolean;
  signal if_stmt_1752_branch_ack_1 : boolean;
  signal array_obj_ref_1698_index_offset_req_1 : boolean;
  signal type_cast_1534_inst_ack_1 : boolean;
  signal type_cast_1534_inst_req_1 : boolean;
  signal type_cast_1534_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1379_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1379_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1379_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1379_inst_ack_1 : boolean;
  signal type_cast_1534_inst_req_0 : boolean;
  signal ptr_deref_1703_load_0_ack_0 : boolean;
  signal ptr_deref_1703_load_0_req_0 : boolean;
  signal type_cast_1692_inst_ack_1 : boolean;
  signal ptr_deref_1392_load_0_req_0 : boolean;
  signal type_cast_1692_inst_req_1 : boolean;
  signal ptr_deref_1392_load_0_ack_0 : boolean;
  signal ptr_deref_1392_load_0_req_1 : boolean;
  signal ptr_deref_1392_load_0_ack_1 : boolean;
  signal ptr_deref_1505_load_0_ack_0 : boolean;
  signal ptr_deref_1487_load_0_ack_1 : boolean;
  signal ptr_deref_1505_load_0_req_0 : boolean;
  signal type_cast_1692_inst_ack_0 : boolean;
  signal type_cast_1692_inst_req_0 : boolean;
  signal ptr_deref_1487_load_0_req_1 : boolean;
  signal ptr_deref_1404_load_0_req_0 : boolean;
  signal ptr_deref_1404_load_0_ack_0 : boolean;
  signal ptr_deref_1404_load_0_req_1 : boolean;
  signal ptr_deref_1404_load_0_ack_1 : boolean;
  signal addr_of_1699_final_reg_ack_1 : boolean;
  signal type_cast_1661_inst_ack_1 : boolean;
  signal type_cast_1661_inst_req_1 : boolean;
  signal type_cast_1661_inst_ack_0 : boolean;
  signal type_cast_1661_inst_req_0 : boolean;
  signal addr_of_1699_final_reg_req_1 : boolean;
  signal ptr_deref_1414_load_0_req_0 : boolean;
  signal ptr_deref_1414_load_0_ack_0 : boolean;
  signal ptr_deref_1414_load_0_req_1 : boolean;
  signal ptr_deref_1414_load_0_ack_1 : boolean;
  signal type_cast_1723_inst_ack_1 : boolean;
  signal addr_of_1699_final_reg_ack_0 : boolean;
  signal type_cast_1539_inst_ack_1 : boolean;
  signal type_cast_1539_inst_req_1 : boolean;
  signal addr_of_1699_final_reg_req_0 : boolean;
  signal type_cast_1723_inst_req_1 : boolean;
  signal type_cast_1418_inst_req_0 : boolean;
  signal type_cast_1418_inst_ack_0 : boolean;
  signal type_cast_1418_inst_req_1 : boolean;
  signal type_cast_1418_inst_ack_1 : boolean;
  signal type_cast_1539_inst_ack_0 : boolean;
  signal type_cast_1539_inst_req_0 : boolean;
  signal ptr_deref_1430_load_0_req_0 : boolean;
  signal ptr_deref_1430_load_0_ack_0 : boolean;
  signal ptr_deref_1430_load_0_req_1 : boolean;
  signal ptr_deref_1430_load_0_ack_1 : boolean;
  signal LOAD_padding_1433_load_0_req_0 : boolean;
  signal LOAD_padding_1433_load_0_ack_0 : boolean;
  signal LOAD_padding_1433_load_0_req_1 : boolean;
  signal LOAD_padding_1433_load_0_ack_1 : boolean;
  signal type_cast_1437_inst_req_0 : boolean;
  signal type_cast_1437_inst_ack_0 : boolean;
  signal type_cast_1437_inst_req_1 : boolean;
  signal type_cast_1437_inst_ack_1 : boolean;
  signal ptr_deref_1447_load_0_req_0 : boolean;
  signal ptr_deref_1447_load_0_ack_0 : boolean;
  signal ptr_deref_1447_load_0_req_1 : boolean;
  signal ptr_deref_1447_load_0_ack_1 : boolean;
  signal type_cast_1451_inst_req_0 : boolean;
  signal type_cast_1451_inst_ack_0 : boolean;
  signal type_cast_1451_inst_req_1 : boolean;
  signal type_cast_1451_inst_ack_1 : boolean;
  signal ptr_deref_1463_load_0_req_0 : boolean;
  signal ptr_deref_1463_load_0_ack_0 : boolean;
  signal ptr_deref_1463_load_0_req_1 : boolean;
  signal ptr_deref_1463_load_0_ack_1 : boolean;
  signal ptr_deref_1475_load_0_req_0 : boolean;
  signal ptr_deref_1475_load_0_ack_0 : boolean;
  signal ptr_deref_1475_load_0_req_1 : boolean;
  signal ptr_deref_1475_load_0_ack_1 : boolean;
  signal ptr_deref_1487_load_0_req_0 : boolean;
  signal ptr_deref_1487_load_0_ack_0 : boolean;
  signal if_stmt_1752_branch_ack_0 : boolean;
  signal type_cast_1776_inst_req_0 : boolean;
  signal type_cast_1776_inst_ack_0 : boolean;
  signal type_cast_1776_inst_req_1 : boolean;
  signal type_cast_1776_inst_ack_1 : boolean;
  signal type_cast_1785_inst_req_0 : boolean;
  signal type_cast_1785_inst_ack_0 : boolean;
  signal type_cast_1785_inst_req_1 : boolean;
  signal type_cast_1785_inst_ack_1 : boolean;
  signal type_cast_1802_inst_req_0 : boolean;
  signal type_cast_1802_inst_ack_0 : boolean;
  signal type_cast_1802_inst_req_1 : boolean;
  signal type_cast_1802_inst_ack_1 : boolean;
  signal if_stmt_1809_branch_req_0 : boolean;
  signal if_stmt_1809_branch_ack_1 : boolean;
  signal if_stmt_1809_branch_ack_0 : boolean;
  signal WPIPE_Block0_done_1817_inst_req_0 : boolean;
  signal WPIPE_Block0_done_1817_inst_ack_0 : boolean;
  signal WPIPE_Block0_done_1817_inst_req_1 : boolean;
  signal WPIPE_Block0_done_1817_inst_ack_1 : boolean;
  signal phi_stmt_1515_req_0 : boolean;
  signal phi_stmt_1522_req_0 : boolean;
  signal type_cast_1521_inst_req_0 : boolean;
  signal type_cast_1521_inst_ack_0 : boolean;
  signal type_cast_1521_inst_req_1 : boolean;
  signal type_cast_1521_inst_ack_1 : boolean;
  signal phi_stmt_1515_req_1 : boolean;
  signal type_cast_1528_inst_req_0 : boolean;
  signal type_cast_1528_inst_ack_0 : boolean;
  signal type_cast_1528_inst_req_1 : boolean;
  signal type_cast_1528_inst_ack_1 : boolean;
  signal phi_stmt_1522_req_1 : boolean;
  signal phi_stmt_1515_ack_0 : boolean;
  signal phi_stmt_1522_ack_0 : boolean;
  signal type_cast_1651_inst_req_0 : boolean;
  signal type_cast_1651_inst_ack_0 : boolean;
  signal type_cast_1651_inst_req_1 : boolean;
  signal type_cast_1651_inst_ack_1 : boolean;
  signal phi_stmt_1645_req_1 : boolean;
  signal phi_stmt_1645_req_0 : boolean;
  signal phi_stmt_1645_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeA_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeA_CP_3995_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeA_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeA_CP_3995_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeA_CP_3995_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeA_CP_3995_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeA_CP_3995: Block -- control-path 
    signal convTransposeA_CP_3995_elements: BooleanArray(88 downto 0);
    -- 
  begin -- 
    convTransposeA_CP_3995_elements(0) <= convTransposeA_CP_3995_start;
    convTransposeA_CP_3995_symbol <= convTransposeA_CP_3995_elements(68);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1377/$entry
      -- CP-element group 0: 	 branch_block_stmt_1377/branch_block_stmt_1377__entry__
      -- CP-element group 0: 	 branch_block_stmt_1377/assign_stmt_1380__entry__
      -- CP-element group 0: 	 branch_block_stmt_1377/assign_stmt_1380/$entry
      -- CP-element group 0: 	 branch_block_stmt_1377/assign_stmt_1380/RPIPE_Block0_start_1379_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1377/assign_stmt_1380/RPIPE_Block0_start_1379_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1377/assign_stmt_1380/RPIPE_Block0_start_1379_Sample/rr
      -- 
    rr_4043_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4043_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(0), ack => RPIPE_Block0_start_1379_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_1377/assign_stmt_1380/RPIPE_Block0_start_1379_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_1377/assign_stmt_1380/RPIPE_Block0_start_1379_update_start_
      -- CP-element group 1: 	 branch_block_stmt_1377/assign_stmt_1380/RPIPE_Block0_start_1379_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_1377/assign_stmt_1380/RPIPE_Block0_start_1379_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_1377/assign_stmt_1380/RPIPE_Block0_start_1379_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1377/assign_stmt_1380/RPIPE_Block0_start_1379_Update/cr
      -- 
    ra_4044_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1379_inst_ack_0, ack => convTransposeA_CP_3995_elements(1)); -- 
    cr_4048_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4048_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(1), ack => RPIPE_Block0_start_1379_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  place  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	20 
    -- CP-element group 2: 	21 
    -- CP-element group 2: 	22 
    -- CP-element group 2: 	17 
    -- CP-element group 2: 	18 
    -- CP-element group 2: 	28 
    -- CP-element group 2: 	23 
    -- CP-element group 2: 	24 
    -- CP-element group 2: 	25 
    -- CP-element group 2: 	26 
    -- CP-element group 2: 	27 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	4 
    -- CP-element group 2: 	5 
    -- CP-element group 2: 	6 
    -- CP-element group 2: 	7 
    -- CP-element group 2: 	8 
    -- CP-element group 2: 	10 
    -- CP-element group 2: 	11 
    -- CP-element group 2: 	12 
    -- CP-element group 2: 	13 
    -- CP-element group 2: 	14 
    -- CP-element group 2: 	16 
    -- CP-element group 2:  members (262) 
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1505_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1505_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1505_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1505_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1505_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1505_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1505_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1505_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1505_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1505_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1505_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1505_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1380__exit__
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512__entry__
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1505_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1505_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1505_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1380/$exit
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1380/RPIPE_Block0_start_1379_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1505_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1380/RPIPE_Block0_start_1379_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1380/RPIPE_Block0_start_1379_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1392_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1392_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1392_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1392_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1392_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1392_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1392_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1392_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1392_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1392_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1392_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1392_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1392_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1392_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1392_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1392_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1392_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1392_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1392_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1392_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1392_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1392_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1392_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1392_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1392_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1392_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1505_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1404_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1505_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1404_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1404_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1404_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1404_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1404_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1404_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1404_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1404_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1404_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1404_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1404_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1404_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1404_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1505_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1404_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1404_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1404_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1404_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1487_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1404_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1404_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1404_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1404_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1404_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1404_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1404_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1404_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1505_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1487_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1414_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1414_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1414_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1414_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1414_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1414_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1414_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1414_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1414_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1414_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1414_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1414_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1414_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1414_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1505_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1414_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1414_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1414_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1414_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1414_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1414_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1414_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1414_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1487_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1414_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1414_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1414_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1414_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1505_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1505_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/type_cast_1418_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1487_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/type_cast_1418_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/type_cast_1418_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1505_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1505_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1430_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1430_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1430_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1430_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1430_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1430_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1430_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1430_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1430_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1430_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1505_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1430_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1430_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1430_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1430_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1430_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1430_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1430_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1430_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1430_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1430_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1430_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1430_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1430_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1430_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1430_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1430_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/LOAD_padding_1433_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/LOAD_padding_1433_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/LOAD_padding_1433_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/LOAD_padding_1433_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/LOAD_padding_1433_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/LOAD_padding_1433_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/LOAD_padding_1433_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/LOAD_padding_1433_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/LOAD_padding_1433_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/LOAD_padding_1433_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/LOAD_padding_1433_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/LOAD_padding_1433_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/type_cast_1437_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/type_cast_1437_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/type_cast_1437_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1447_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1447_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1447_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1447_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1447_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1447_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1447_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1447_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1447_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1447_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1447_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1447_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1447_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1447_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1447_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1447_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1447_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1447_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1447_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1447_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1447_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1447_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1447_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1447_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1447_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1447_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/type_cast_1451_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/type_cast_1451_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/type_cast_1451_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1463_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1463_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1463_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1463_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1463_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1463_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1463_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1463_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1463_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1463_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1463_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1463_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1463_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1463_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1463_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1463_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1463_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1463_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1463_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1463_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1463_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1463_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1463_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1463_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1463_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1463_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1475_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1475_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1475_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1475_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1475_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1475_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1475_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1475_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1475_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1475_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1475_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1475_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1475_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1475_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1475_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1475_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1475_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1475_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1475_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1475_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1475_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1475_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1475_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1475_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1475_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1475_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1487_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1487_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1487_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1487_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1487_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1487_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1487_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1487_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1487_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1487_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1487_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1487_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1487_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1487_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1487_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1487_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1487_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1487_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1487_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1487_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1487_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1487_Sample/word_access_start/word_0/rr
      -- 
    ca_4049_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1379_inst_ack_1, ack => convTransposeA_CP_3995_elements(2)); -- 
    cr_4571_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4571_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(2), ack => ptr_deref_1505_load_0_req_1); -- 
    rr_4085_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4085_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(2), ack => ptr_deref_1392_load_0_req_0); -- 
    cr_4096_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4096_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(2), ack => ptr_deref_1392_load_0_req_1); -- 
    rr_4560_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4560_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(2), ack => ptr_deref_1505_load_0_req_0); -- 
    cr_4521_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4521_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(2), ack => ptr_deref_1487_load_0_req_1); -- 
    rr_4135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(2), ack => ptr_deref_1404_load_0_req_0); -- 
    cr_4146_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4146_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(2), ack => ptr_deref_1404_load_0_req_1); -- 
    rr_4185_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4185_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(2), ack => ptr_deref_1414_load_0_req_0); -- 
    cr_4196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(2), ack => ptr_deref_1414_load_0_req_1); -- 
    cr_4215_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4215_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(2), ack => type_cast_1418_inst_req_1); -- 
    rr_4249_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4249_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(2), ack => ptr_deref_1430_load_0_req_0); -- 
    cr_4260_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4260_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(2), ack => ptr_deref_1430_load_0_req_1); -- 
    rr_4282_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4282_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(2), ack => LOAD_padding_1433_load_0_req_0); -- 
    cr_4293_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4293_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(2), ack => LOAD_padding_1433_load_0_req_1); -- 
    cr_4312_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4312_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(2), ack => type_cast_1437_inst_req_1); -- 
    rr_4346_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4346_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(2), ack => ptr_deref_1447_load_0_req_0); -- 
    cr_4357_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4357_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(2), ack => ptr_deref_1447_load_0_req_1); -- 
    cr_4376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(2), ack => type_cast_1451_inst_req_1); -- 
    rr_4410_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4410_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(2), ack => ptr_deref_1463_load_0_req_0); -- 
    cr_4421_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4421_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(2), ack => ptr_deref_1463_load_0_req_1); -- 
    rr_4460_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4460_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(2), ack => ptr_deref_1475_load_0_req_0); -- 
    cr_4471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(2), ack => ptr_deref_1475_load_0_req_1); -- 
    rr_4510_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4510_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(2), ack => ptr_deref_1487_load_0_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (5) 
      -- CP-element group 3: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1392_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1392_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1392_Sample/word_access_start/$exit
      -- CP-element group 3: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1392_Sample/word_access_start/word_0/$exit
      -- CP-element group 3: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1392_Sample/word_access_start/word_0/ra
      -- 
    ra_4086_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1392_load_0_ack_0, ack => convTransposeA_CP_3995_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	2 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	29 
    -- CP-element group 4:  members (9) 
      -- CP-element group 4: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1392_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1392_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1392_Update/word_access_complete/$exit
      -- CP-element group 4: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1392_Update/word_access_complete/word_0/$exit
      -- CP-element group 4: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1392_Update/word_access_complete/word_0/ca
      -- CP-element group 4: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1392_Update/ptr_deref_1392_Merge/$entry
      -- CP-element group 4: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1392_Update/ptr_deref_1392_Merge/$exit
      -- CP-element group 4: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1392_Update/ptr_deref_1392_Merge/merge_req
      -- CP-element group 4: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1392_Update/ptr_deref_1392_Merge/merge_ack
      -- 
    ca_4097_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1392_load_0_ack_1, ack => convTransposeA_CP_3995_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (5) 
      -- CP-element group 5: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1404_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1404_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1404_Sample/word_access_start/$exit
      -- CP-element group 5: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1404_Sample/word_access_start/word_0/$exit
      -- CP-element group 5: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1404_Sample/word_access_start/word_0/ra
      -- 
    ra_4136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1404_load_0_ack_0, ack => convTransposeA_CP_3995_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	2 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	29 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1404_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1404_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1404_Update/word_access_complete/$exit
      -- CP-element group 6: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1404_Update/word_access_complete/word_0/$exit
      -- CP-element group 6: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1404_Update/word_access_complete/word_0/ca
      -- CP-element group 6: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1404_Update/ptr_deref_1404_Merge/$entry
      -- CP-element group 6: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1404_Update/ptr_deref_1404_Merge/$exit
      -- CP-element group 6: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1404_Update/ptr_deref_1404_Merge/merge_req
      -- CP-element group 6: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1404_Update/ptr_deref_1404_Merge/merge_ack
      -- 
    ca_4147_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1404_load_0_ack_1, ack => convTransposeA_CP_3995_elements(6)); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	2 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (5) 
      -- CP-element group 7: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1414_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1414_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1414_Sample/word_access_start/$exit
      -- CP-element group 7: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1414_Sample/word_access_start/word_0/$exit
      -- CP-element group 7: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1414_Sample/word_access_start/word_0/ra
      -- 
    ra_4186_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1414_load_0_ack_0, ack => convTransposeA_CP_3995_elements(7)); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (12) 
      -- CP-element group 8: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1414_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1414_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1414_Update/word_access_complete/$exit
      -- CP-element group 8: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1414_Update/word_access_complete/word_0/$exit
      -- CP-element group 8: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1414_Update/word_access_complete/word_0/ca
      -- CP-element group 8: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1414_Update/ptr_deref_1414_Merge/$entry
      -- CP-element group 8: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1414_Update/ptr_deref_1414_Merge/$exit
      -- CP-element group 8: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1414_Update/ptr_deref_1414_Merge/merge_req
      -- CP-element group 8: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1414_Update/ptr_deref_1414_Merge/merge_ack
      -- CP-element group 8: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/type_cast_1418_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/type_cast_1418_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/type_cast_1418_Sample/rr
      -- 
    ca_4197_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1414_load_0_ack_1, ack => convTransposeA_CP_3995_elements(8)); -- 
    rr_4210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(8), ack => type_cast_1418_inst_req_0); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/type_cast_1418_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/type_cast_1418_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/type_cast_1418_Sample/ra
      -- 
    ra_4211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1418_inst_ack_0, ack => convTransposeA_CP_3995_elements(9)); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	2 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	29 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/type_cast_1418_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/type_cast_1418_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/type_cast_1418_Update/ca
      -- 
    ca_4216_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1418_inst_ack_1, ack => convTransposeA_CP_3995_elements(10)); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	2 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (5) 
      -- CP-element group 11: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1430_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1430_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1430_Sample/word_access_start/$exit
      -- CP-element group 11: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1430_Sample/word_access_start/word_0/$exit
      -- CP-element group 11: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1430_Sample/word_access_start/word_0/ra
      -- 
    ra_4250_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1430_load_0_ack_0, ack => convTransposeA_CP_3995_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	2 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	29 
    -- CP-element group 12:  members (9) 
      -- CP-element group 12: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1430_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1430_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1430_Update/word_access_complete/$exit
      -- CP-element group 12: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1430_Update/word_access_complete/word_0/$exit
      -- CP-element group 12: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1430_Update/word_access_complete/word_0/ca
      -- CP-element group 12: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1430_Update/ptr_deref_1430_Merge/$entry
      -- CP-element group 12: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1430_Update/ptr_deref_1430_Merge/$exit
      -- CP-element group 12: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1430_Update/ptr_deref_1430_Merge/merge_req
      -- CP-element group 12: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1430_Update/ptr_deref_1430_Merge/merge_ack
      -- 
    ca_4261_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1430_load_0_ack_1, ack => convTransposeA_CP_3995_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	2 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (5) 
      -- CP-element group 13: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/LOAD_padding_1433_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/LOAD_padding_1433_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/LOAD_padding_1433_Sample/word_access_start/$exit
      -- CP-element group 13: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/LOAD_padding_1433_Sample/word_access_start/word_0/$exit
      -- CP-element group 13: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/LOAD_padding_1433_Sample/word_access_start/word_0/ra
      -- 
    ra_4283_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_padding_1433_load_0_ack_0, ack => convTransposeA_CP_3995_elements(13)); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	2 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (12) 
      -- CP-element group 14: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/LOAD_padding_1433_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/LOAD_padding_1433_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/LOAD_padding_1433_Update/word_access_complete/$exit
      -- CP-element group 14: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/LOAD_padding_1433_Update/word_access_complete/word_0/$exit
      -- CP-element group 14: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/LOAD_padding_1433_Update/word_access_complete/word_0/ca
      -- CP-element group 14: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/LOAD_padding_1433_Update/LOAD_padding_1433_Merge/$entry
      -- CP-element group 14: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/LOAD_padding_1433_Update/LOAD_padding_1433_Merge/$exit
      -- CP-element group 14: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/LOAD_padding_1433_Update/LOAD_padding_1433_Merge/merge_req
      -- CP-element group 14: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/LOAD_padding_1433_Update/LOAD_padding_1433_Merge/merge_ack
      -- CP-element group 14: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/type_cast_1437_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/type_cast_1437_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/type_cast_1437_Sample/rr
      -- 
    ca_4294_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_padding_1433_load_0_ack_1, ack => convTransposeA_CP_3995_elements(14)); -- 
    rr_4307_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4307_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(14), ack => type_cast_1437_inst_req_0); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/type_cast_1437_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/type_cast_1437_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/type_cast_1437_Sample/ra
      -- 
    ra_4308_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1437_inst_ack_0, ack => convTransposeA_CP_3995_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	2 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	29 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/type_cast_1437_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/type_cast_1437_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/type_cast_1437_Update/ca
      -- 
    ca_4313_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1437_inst_ack_1, ack => convTransposeA_CP_3995_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	2 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (5) 
      -- CP-element group 17: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1447_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1447_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1447_Sample/word_access_start/$exit
      -- CP-element group 17: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1447_Sample/word_access_start/word_0/$exit
      -- CP-element group 17: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1447_Sample/word_access_start/word_0/ra
      -- 
    ra_4347_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1447_load_0_ack_0, ack => convTransposeA_CP_3995_elements(17)); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	2 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (12) 
      -- CP-element group 18: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1447_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1447_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1447_Update/word_access_complete/$exit
      -- CP-element group 18: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1447_Update/word_access_complete/word_0/$exit
      -- CP-element group 18: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1447_Update/word_access_complete/word_0/ca
      -- CP-element group 18: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1447_Update/ptr_deref_1447_Merge/$entry
      -- CP-element group 18: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1447_Update/ptr_deref_1447_Merge/$exit
      -- CP-element group 18: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1447_Update/ptr_deref_1447_Merge/merge_req
      -- CP-element group 18: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1447_Update/ptr_deref_1447_Merge/merge_ack
      -- CP-element group 18: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/type_cast_1451_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/type_cast_1451_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/type_cast_1451_Sample/rr
      -- 
    ca_4358_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1447_load_0_ack_1, ack => convTransposeA_CP_3995_elements(18)); -- 
    rr_4371_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4371_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(18), ack => type_cast_1451_inst_req_0); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/type_cast_1451_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/type_cast_1451_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/type_cast_1451_Sample/ra
      -- 
    ra_4372_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1451_inst_ack_0, ack => convTransposeA_CP_3995_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	2 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	29 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/type_cast_1451_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/type_cast_1451_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/type_cast_1451_Update/ca
      -- 
    ca_4377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1451_inst_ack_1, ack => convTransposeA_CP_3995_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	2 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (5) 
      -- CP-element group 21: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1463_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1463_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1463_Sample/word_access_start/$exit
      -- CP-element group 21: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1463_Sample/word_access_start/word_0/$exit
      -- CP-element group 21: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1463_Sample/word_access_start/word_0/ra
      -- 
    ra_4411_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1463_load_0_ack_0, ack => convTransposeA_CP_3995_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	2 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	29 
    -- CP-element group 22:  members (9) 
      -- CP-element group 22: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1463_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1463_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1463_Update/word_access_complete/$exit
      -- CP-element group 22: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1463_Update/word_access_complete/word_0/$exit
      -- CP-element group 22: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1463_Update/word_access_complete/word_0/ca
      -- CP-element group 22: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1463_Update/ptr_deref_1463_Merge/$entry
      -- CP-element group 22: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1463_Update/ptr_deref_1463_Merge/$exit
      -- CP-element group 22: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1463_Update/ptr_deref_1463_Merge/merge_req
      -- CP-element group 22: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1463_Update/ptr_deref_1463_Merge/merge_ack
      -- 
    ca_4422_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1463_load_0_ack_1, ack => convTransposeA_CP_3995_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	2 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (5) 
      -- CP-element group 23: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1475_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1475_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1475_Sample/word_access_start/$exit
      -- CP-element group 23: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1475_Sample/word_access_start/word_0/$exit
      -- CP-element group 23: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1475_Sample/word_access_start/word_0/ra
      -- 
    ra_4461_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1475_load_0_ack_0, ack => convTransposeA_CP_3995_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	2 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	29 
    -- CP-element group 24:  members (9) 
      -- CP-element group 24: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1475_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1475_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1475_Update/word_access_complete/$exit
      -- CP-element group 24: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1475_Update/word_access_complete/word_0/$exit
      -- CP-element group 24: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1475_Update/word_access_complete/word_0/ca
      -- CP-element group 24: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1475_Update/ptr_deref_1475_Merge/$entry
      -- CP-element group 24: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1475_Update/ptr_deref_1475_Merge/$exit
      -- CP-element group 24: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1475_Update/ptr_deref_1475_Merge/merge_req
      -- CP-element group 24: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1475_Update/ptr_deref_1475_Merge/merge_ack
      -- 
    ca_4472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1475_load_0_ack_1, ack => convTransposeA_CP_3995_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	2 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (5) 
      -- CP-element group 25: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1487_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1487_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1487_Sample/word_access_start/$exit
      -- CP-element group 25: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1487_Sample/word_access_start/word_0/$exit
      -- CP-element group 25: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1487_Sample/word_access_start/word_0/ra
      -- 
    ra_4511_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1487_load_0_ack_0, ack => convTransposeA_CP_3995_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	2 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	29 
    -- CP-element group 26:  members (9) 
      -- CP-element group 26: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1487_Update/ptr_deref_1487_Merge/merge_ack
      -- CP-element group 26: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1487_Update/ptr_deref_1487_Merge/merge_req
      -- CP-element group 26: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1487_Update/ptr_deref_1487_Merge/$exit
      -- CP-element group 26: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1487_Update/ptr_deref_1487_Merge/$entry
      -- CP-element group 26: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1487_Update/word_access_complete/word_0/ca
      -- CP-element group 26: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1487_Update/word_access_complete/word_0/$exit
      -- CP-element group 26: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1487_Update/word_access_complete/$exit
      -- CP-element group 26: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1487_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1487_update_completed_
      -- 
    ca_4522_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1487_load_0_ack_1, ack => convTransposeA_CP_3995_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	2 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (5) 
      -- CP-element group 27: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1505_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1505_Sample/word_access_start/word_0/ra
      -- CP-element group 27: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1505_Sample/word_access_start/word_0/$exit
      -- CP-element group 27: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1505_Sample/word_access_start/$exit
      -- CP-element group 27: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1505_Sample/$exit
      -- 
    ra_4561_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1505_load_0_ack_0, ack => convTransposeA_CP_3995_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	2 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (9) 
      -- CP-element group 28: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1505_Update/word_access_complete/word_0/ca
      -- CP-element group 28: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1505_Update/ptr_deref_1505_Merge/merge_req
      -- CP-element group 28: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1505_Update/ptr_deref_1505_Merge/$entry
      -- CP-element group 28: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1505_Update/ptr_deref_1505_Merge/$exit
      -- CP-element group 28: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1505_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1505_Update/word_access_complete/word_0/$exit
      -- CP-element group 28: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1505_Update/word_access_complete/$exit
      -- CP-element group 28: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1505_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/ptr_deref_1505_Update/ptr_deref_1505_Merge/merge_ack
      -- 
    ca_4572_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1505_load_0_ack_1, ack => convTransposeA_CP_3995_elements(28)); -- 
    -- CP-element group 29:  join  fork  transition  place  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	20 
    -- CP-element group 29: 	22 
    -- CP-element group 29: 	28 
    -- CP-element group 29: 	24 
    -- CP-element group 29: 	26 
    -- CP-element group 29: 	4 
    -- CP-element group 29: 	6 
    -- CP-element group 29: 	10 
    -- CP-element group 29: 	12 
    -- CP-element group 29: 	16 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	69 
    -- CP-element group 29: 	70 
    -- CP-element group 29:  members (8) 
      -- CP-element group 29: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512__exit__
      -- CP-element group 29: 	 branch_block_stmt_1377/entry_whilex_xbodyx_xouter
      -- CP-element group 29: 	 branch_block_stmt_1377/assign_stmt_1389_to_assign_stmt_1512/$exit
      -- CP-element group 29: 	 branch_block_stmt_1377/entry_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 29: 	 branch_block_stmt_1377/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1515/$entry
      -- CP-element group 29: 	 branch_block_stmt_1377/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1515/phi_stmt_1515_sources/$entry
      -- CP-element group 29: 	 branch_block_stmt_1377/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1522/$entry
      -- CP-element group 29: 	 branch_block_stmt_1377/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1522/phi_stmt_1522_sources/$entry
      -- 
    convTransposeA_cp_element_group_29: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_29"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= convTransposeA_CP_3995_elements(20) & convTransposeA_CP_3995_elements(22) & convTransposeA_CP_3995_elements(28) & convTransposeA_CP_3995_elements(24) & convTransposeA_CP_3995_elements(26) & convTransposeA_CP_3995_elements(4) & convTransposeA_CP_3995_elements(6) & convTransposeA_CP_3995_elements(10) & convTransposeA_CP_3995_elements(12) & convTransposeA_CP_3995_elements(16);
      gj_convTransposeA_cp_element_group_29 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3995_elements(29), clk => clk, reset => reset); --
    end block;
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	82 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_1377/assign_stmt_1535_to_assign_stmt_1642/type_cast_1534_Sample/ra
      -- CP-element group 30: 	 branch_block_stmt_1377/assign_stmt_1535_to_assign_stmt_1642/type_cast_1534_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_1377/assign_stmt_1535_to_assign_stmt_1642/type_cast_1534_sample_completed_
      -- 
    ra_4589_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1534_inst_ack_0, ack => convTransposeA_CP_3995_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	82 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	34 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_1377/assign_stmt_1535_to_assign_stmt_1642/type_cast_1534_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_1377/assign_stmt_1535_to_assign_stmt_1642/type_cast_1534_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_1377/assign_stmt_1535_to_assign_stmt_1642/type_cast_1534_update_completed_
      -- 
    ca_4594_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1534_inst_ack_1, ack => convTransposeA_CP_3995_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	82 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_1377/assign_stmt_1535_to_assign_stmt_1642/type_cast_1539_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_1377/assign_stmt_1535_to_assign_stmt_1642/type_cast_1539_Sample/ra
      -- CP-element group 32: 	 branch_block_stmt_1377/assign_stmt_1535_to_assign_stmt_1642/type_cast_1539_Sample/$exit
      -- 
    ra_4603_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1539_inst_ack_0, ack => convTransposeA_CP_3995_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	82 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_1377/assign_stmt_1535_to_assign_stmt_1642/type_cast_1539_Update/ca
      -- CP-element group 33: 	 branch_block_stmt_1377/assign_stmt_1535_to_assign_stmt_1642/type_cast_1539_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_1377/assign_stmt_1535_to_assign_stmt_1642/type_cast_1539_update_completed_
      -- 
    ca_4608_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1539_inst_ack_1, ack => convTransposeA_CP_3995_elements(33)); -- 
    -- CP-element group 34:  join  transition  place  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	31 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	86 
    -- CP-element group 34:  members (6) 
      -- CP-element group 34: 	 branch_block_stmt_1377/assign_stmt_1535_to_assign_stmt_1642__exit__
      -- CP-element group 34: 	 branch_block_stmt_1377/whilex_xbodyx_xouter_whilex_xbody
      -- CP-element group 34: 	 branch_block_stmt_1377/assign_stmt_1535_to_assign_stmt_1642/$exit
      -- CP-element group 34: 	 branch_block_stmt_1377/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$entry
      -- CP-element group 34: 	 branch_block_stmt_1377/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1645/$entry
      -- CP-element group 34: 	 branch_block_stmt_1377/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1645/phi_stmt_1645_sources/$entry
      -- 
    convTransposeA_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3995_elements(31) & convTransposeA_CP_3995_elements(33);
      gj_convTransposeA_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3995_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	88 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/type_cast_1661_Sample/ra
      -- CP-element group 35: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/type_cast_1661_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/type_cast_1661_sample_completed_
      -- 
    ra_4620_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1661_inst_ack_0, ack => convTransposeA_CP_3995_elements(35)); -- 
    -- CP-element group 36:  fork  transition  input  output  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	88 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	37 
    -- CP-element group 36: 	45 
    -- CP-element group 36:  members (9) 
      -- CP-element group 36: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/type_cast_1723_Sample/$entry
      -- CP-element group 36: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/type_cast_1723_Sample/rr
      -- CP-element group 36: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/type_cast_1692_Sample/rr
      -- CP-element group 36: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/type_cast_1692_Sample/$entry
      -- CP-element group 36: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/type_cast_1692_sample_start_
      -- CP-element group 36: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/type_cast_1723_sample_start_
      -- CP-element group 36: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/type_cast_1661_Update/ca
      -- CP-element group 36: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/type_cast_1661_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/type_cast_1661_update_completed_
      -- 
    ca_4625_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1661_inst_ack_1, ack => convTransposeA_CP_3995_elements(36)); -- 
    rr_4633_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4633_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(36), ack => type_cast_1692_inst_req_0); -- 
    rr_4743_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4743_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(36), ack => type_cast_1723_inst_req_0); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	36 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/type_cast_1692_Sample/ra
      -- CP-element group 37: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/type_cast_1692_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/type_cast_1692_sample_completed_
      -- 
    ra_4634_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1692_inst_ack_0, ack => convTransposeA_CP_3995_elements(37)); -- 
    -- CP-element group 38:  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	88 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (16) 
      -- CP-element group 38: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/array_obj_ref_1698_index_scale_1/scale_rename_req
      -- CP-element group 38: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/array_obj_ref_1698_index_resized_1
      -- CP-element group 38: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/array_obj_ref_1698_index_resize_1/index_resize_req
      -- CP-element group 38: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/array_obj_ref_1698_final_index_sum_regn_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/array_obj_ref_1698_index_scaled_1
      -- CP-element group 38: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/array_obj_ref_1698_index_resize_1/index_resize_ack
      -- CP-element group 38: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/array_obj_ref_1698_index_computed_1
      -- CP-element group 38: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/array_obj_ref_1698_index_scale_1/$entry
      -- CP-element group 38: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/array_obj_ref_1698_index_scale_1/$exit
      -- CP-element group 38: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/array_obj_ref_1698_index_resize_1/$exit
      -- CP-element group 38: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/array_obj_ref_1698_final_index_sum_regn_Sample/req
      -- CP-element group 38: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/array_obj_ref_1698_index_scale_1/scale_rename_ack
      -- CP-element group 38: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/array_obj_ref_1698_index_resize_1/$entry
      -- CP-element group 38: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/type_cast_1692_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/type_cast_1692_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/type_cast_1692_update_completed_
      -- 
    ca_4639_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1692_inst_ack_1, ack => convTransposeA_CP_3995_elements(38)); -- 
    req_4664_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4664_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(38), ack => array_obj_ref_1698_index_offset_req_0); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	56 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/array_obj_ref_1698_final_index_sum_regn_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/array_obj_ref_1698_final_index_sum_regn_Sample/ack
      -- CP-element group 39: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/array_obj_ref_1698_final_index_sum_regn_sample_complete
      -- 
    ack_4665_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1698_index_offset_ack_0, ack => convTransposeA_CP_3995_elements(39)); -- 
    -- CP-element group 40:  transition  input  output  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	88 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (11) 
      -- CP-element group 40: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/array_obj_ref_1698_offset_calculated
      -- CP-element group 40: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/array_obj_ref_1698_base_plus_offset/$entry
      -- CP-element group 40: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/array_obj_ref_1698_base_plus_offset/$exit
      -- CP-element group 40: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/array_obj_ref_1698_base_plus_offset/sum_rename_req
      -- CP-element group 40: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/array_obj_ref_1698_final_index_sum_regn_Update/ack
      -- CP-element group 40: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/array_obj_ref_1698_base_plus_offset/sum_rename_ack
      -- CP-element group 40: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/array_obj_ref_1698_root_address_calculated
      -- CP-element group 40: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/array_obj_ref_1698_final_index_sum_regn_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/addr_of_1699_sample_start_
      -- CP-element group 40: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/addr_of_1699_request/req
      -- CP-element group 40: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/addr_of_1699_request/$entry
      -- 
    ack_4670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1698_index_offset_ack_1, ack => convTransposeA_CP_3995_elements(40)); -- 
    req_4679_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4679_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(40), ack => addr_of_1699_final_reg_req_0); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/addr_of_1699_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/addr_of_1699_request/ack
      -- CP-element group 41: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/addr_of_1699_request/$exit
      -- 
    ack_4680_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1699_final_reg_ack_0, ack => convTransposeA_CP_3995_elements(41)); -- 
    -- CP-element group 42:  join  fork  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	88 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (24) 
      -- CP-element group 42: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1703_word_addrgen/root_register_req
      -- CP-element group 42: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1703_base_plus_offset/sum_rename_ack
      -- CP-element group 42: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1703_base_plus_offset/sum_rename_req
      -- CP-element group 42: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1703_word_addrgen/$entry
      -- CP-element group 42: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1703_base_plus_offset/$exit
      -- CP-element group 42: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1703_base_plus_offset/$entry
      -- CP-element group 42: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1703_base_addr_resize/base_resize_ack
      -- CP-element group 42: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1703_word_addrgen/$exit
      -- CP-element group 42: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1703_base_addr_resize/base_resize_req
      -- CP-element group 42: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1703_base_addr_resize/$exit
      -- CP-element group 42: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1703_base_addr_resize/$entry
      -- CP-element group 42: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1703_base_address_resized
      -- CP-element group 42: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1703_Sample/word_access_start/word_0/rr
      -- CP-element group 42: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1703_Sample/word_access_start/word_0/$entry
      -- CP-element group 42: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1703_root_address_calculated
      -- CP-element group 42: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/addr_of_1699_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1703_word_address_calculated
      -- CP-element group 42: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1703_base_address_calculated
      -- CP-element group 42: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1703_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/addr_of_1699_complete/ack
      -- CP-element group 42: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1703_Sample/word_access_start/$entry
      -- CP-element group 42: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/addr_of_1699_complete/$exit
      -- CP-element group 42: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1703_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1703_word_addrgen/root_register_ack
      -- 
    ack_4685_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1699_final_reg_ack_1, ack => convTransposeA_CP_3995_elements(42)); -- 
    rr_4718_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4718_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(42), ack => ptr_deref_1703_load_0_req_0); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (5) 
      -- CP-element group 43: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1703_Sample/word_access_start/word_0/ra
      -- CP-element group 43: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1703_Sample/word_access_start/word_0/$exit
      -- CP-element group 43: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1703_Sample/word_access_start/$exit
      -- CP-element group 43: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1703_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1703_Sample/$exit
      -- 
    ra_4719_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1703_load_0_ack_0, ack => convTransposeA_CP_3995_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	88 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	51 
    -- CP-element group 44:  members (9) 
      -- CP-element group 44: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1703_Update/word_access_complete/word_0/ca
      -- CP-element group 44: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1703_Update/ptr_deref_1703_Merge/$entry
      -- CP-element group 44: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1703_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1703_Update/word_access_complete/$exit
      -- CP-element group 44: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1703_Update/ptr_deref_1703_Merge/merge_ack
      -- CP-element group 44: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1703_Update/word_access_complete/word_0/$exit
      -- CP-element group 44: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1703_Update/ptr_deref_1703_Merge/merge_req
      -- CP-element group 44: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1703_Update/ptr_deref_1703_Merge/$exit
      -- CP-element group 44: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1703_update_completed_
      -- 
    ca_4730_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1703_load_0_ack_1, ack => convTransposeA_CP_3995_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	36 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/type_cast_1723_Sample/ra
      -- CP-element group 45: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/type_cast_1723_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/type_cast_1723_sample_completed_
      -- 
    ra_4744_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1723_inst_ack_0, ack => convTransposeA_CP_3995_elements(45)); -- 
    -- CP-element group 46:  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	88 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (16) 
      -- CP-element group 46: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/array_obj_ref_1729_index_resized_1
      -- CP-element group 46: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/array_obj_ref_1729_index_computed_1
      -- CP-element group 46: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/array_obj_ref_1729_index_scale_1/scale_rename_ack
      -- CP-element group 46: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/array_obj_ref_1729_final_index_sum_regn_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/array_obj_ref_1729_final_index_sum_regn_Sample/req
      -- CP-element group 46: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/array_obj_ref_1729_index_scale_1/scale_rename_req
      -- CP-element group 46: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/array_obj_ref_1729_index_scale_1/$exit
      -- CP-element group 46: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/array_obj_ref_1729_index_scaled_1
      -- CP-element group 46: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/array_obj_ref_1729_index_scale_1/$entry
      -- CP-element group 46: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/array_obj_ref_1729_index_resize_1/index_resize_ack
      -- CP-element group 46: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/array_obj_ref_1729_index_resize_1/index_resize_req
      -- CP-element group 46: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/array_obj_ref_1729_index_resize_1/$exit
      -- CP-element group 46: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/array_obj_ref_1729_index_resize_1/$entry
      -- CP-element group 46: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/type_cast_1723_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/type_cast_1723_Update/ca
      -- CP-element group 46: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/type_cast_1723_Update/$exit
      -- 
    ca_4749_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1723_inst_ack_1, ack => convTransposeA_CP_3995_elements(46)); -- 
    req_4774_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4774_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(46), ack => array_obj_ref_1729_index_offset_req_0); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	56 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/array_obj_ref_1729_final_index_sum_regn_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/array_obj_ref_1729_final_index_sum_regn_sample_complete
      -- CP-element group 47: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/array_obj_ref_1729_final_index_sum_regn_Sample/ack
      -- 
    ack_4775_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1729_index_offset_ack_0, ack => convTransposeA_CP_3995_elements(47)); -- 
    -- CP-element group 48:  transition  input  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	88 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (11) 
      -- CP-element group 48: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/array_obj_ref_1729_final_index_sum_regn_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/array_obj_ref_1729_final_index_sum_regn_Update/ack
      -- CP-element group 48: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/array_obj_ref_1729_base_plus_offset/$entry
      -- CP-element group 48: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/array_obj_ref_1729_base_plus_offset/$exit
      -- CP-element group 48: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/array_obj_ref_1729_base_plus_offset/sum_rename_req
      -- CP-element group 48: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/addr_of_1730_request/req
      -- CP-element group 48: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/array_obj_ref_1729_root_address_calculated
      -- CP-element group 48: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/array_obj_ref_1729_offset_calculated
      -- CP-element group 48: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/array_obj_ref_1729_base_plus_offset/sum_rename_ack
      -- CP-element group 48: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/addr_of_1730_sample_start_
      -- CP-element group 48: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/addr_of_1730_request/$entry
      -- 
    ack_4780_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1729_index_offset_ack_1, ack => convTransposeA_CP_3995_elements(48)); -- 
    req_4789_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4789_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(48), ack => addr_of_1730_final_reg_req_0); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/addr_of_1730_request/ack
      -- CP-element group 49: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/addr_of_1730_request/$exit
      -- CP-element group 49: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/addr_of_1730_sample_completed_
      -- 
    ack_4790_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1730_final_reg_ack_0, ack => convTransposeA_CP_3995_elements(49)); -- 
    -- CP-element group 50:  fork  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	88 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (19) 
      -- CP-element group 50: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1733_base_addr_resize/base_resize_req
      -- CP-element group 50: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1733_base_addr_resize/base_resize_ack
      -- CP-element group 50: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/addr_of_1730_complete/$exit
      -- CP-element group 50: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1733_word_address_calculated
      -- CP-element group 50: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1733_base_address_calculated
      -- CP-element group 50: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1733_word_addrgen/root_register_ack
      -- CP-element group 50: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1733_base_address_resized
      -- CP-element group 50: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1733_base_addr_resize/$entry
      -- CP-element group 50: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1733_base_plus_offset/sum_rename_req
      -- CP-element group 50: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1733_root_address_calculated
      -- CP-element group 50: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1733_base_addr_resize/$exit
      -- CP-element group 50: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1733_word_addrgen/root_register_req
      -- CP-element group 50: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1733_word_addrgen/$entry
      -- CP-element group 50: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1733_word_addrgen/$exit
      -- CP-element group 50: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1733_base_plus_offset/sum_rename_ack
      -- CP-element group 50: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1733_base_plus_offset/$entry
      -- CP-element group 50: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1733_base_plus_offset/$exit
      -- CP-element group 50: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/addr_of_1730_complete/ack
      -- CP-element group 50: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/addr_of_1730_update_completed_
      -- 
    ack_4795_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1730_final_reg_ack_1, ack => convTransposeA_CP_3995_elements(50)); -- 
    -- CP-element group 51:  join  transition  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	44 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (9) 
      -- CP-element group 51: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1733_Sample/word_access_start/word_0/$entry
      -- CP-element group 51: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1733_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1733_Sample/ptr_deref_1733_Split/split_ack
      -- CP-element group 51: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1733_Sample/ptr_deref_1733_Split/$entry
      -- CP-element group 51: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1733_Sample/ptr_deref_1733_Split/$exit
      -- CP-element group 51: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1733_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1733_Sample/ptr_deref_1733_Split/split_req
      -- CP-element group 51: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1733_Sample/word_access_start/$entry
      -- CP-element group 51: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1733_Sample/word_access_start/word_0/rr
      -- 
    rr_4833_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4833_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(51), ack => ptr_deref_1733_store_0_req_0); -- 
    convTransposeA_cp_element_group_51: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_51"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3995_elements(44) & convTransposeA_CP_3995_elements(50);
      gj_convTransposeA_cp_element_group_51 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3995_elements(51), clk => clk, reset => reset); --
    end block;
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (5) 
      -- CP-element group 52: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1733_Sample/word_access_start/word_0/$exit
      -- CP-element group 52: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1733_Sample/word_access_start/word_0/ra
      -- CP-element group 52: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1733_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1733_Sample/word_access_start/$exit
      -- CP-element group 52: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1733_sample_completed_
      -- 
    ra_4834_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1733_store_0_ack_0, ack => convTransposeA_CP_3995_elements(52)); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	88 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	56 
    -- CP-element group 53:  members (5) 
      -- CP-element group 53: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1733_Update/word_access_complete/word_0/ca
      -- CP-element group 53: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1733_Update/word_access_complete/word_0/$exit
      -- CP-element group 53: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1733_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1733_Update/word_access_complete/$exit
      -- CP-element group 53: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1733_update_completed_
      -- 
    ca_4845_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1733_store_0_ack_1, ack => convTransposeA_CP_3995_elements(53)); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	88 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/type_cast_1739_Sample/ra
      -- CP-element group 54: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/type_cast_1739_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/type_cast_1739_sample_completed_
      -- 
    ra_4854_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1739_inst_ack_0, ack => convTransposeA_CP_3995_elements(54)); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	88 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/type_cast_1739_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/type_cast_1739_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/type_cast_1739_Update/ca
      -- 
    ca_4859_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1739_inst_ack_1, ack => convTransposeA_CP_3995_elements(55)); -- 
    -- CP-element group 56:  branch  join  transition  place  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	39 
    -- CP-element group 56: 	47 
    -- CP-element group 56: 	53 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56: 	58 
    -- CP-element group 56:  members (10) 
      -- CP-element group 56: 	 branch_block_stmt_1377/if_stmt_1752_eval_test/$exit
      -- CP-element group 56: 	 branch_block_stmt_1377/if_stmt_1752_eval_test/branch_req
      -- CP-element group 56: 	 branch_block_stmt_1377/if_stmt_1752_if_link/$entry
      -- CP-element group 56: 	 branch_block_stmt_1377/if_stmt_1752_dead_link/$entry
      -- CP-element group 56: 	 branch_block_stmt_1377/if_stmt_1752_eval_test/$entry
      -- CP-element group 56: 	 branch_block_stmt_1377/if_stmt_1752_else_link/$entry
      -- CP-element group 56: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751__exit__
      -- CP-element group 56: 	 branch_block_stmt_1377/if_stmt_1752__entry__
      -- CP-element group 56: 	 branch_block_stmt_1377/R_cmp_1753_place
      -- CP-element group 56: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/$exit
      -- 
    branch_req_4867_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4867_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(56), ack => if_stmt_1752_branch_req_0); -- 
    convTransposeA_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_3995_elements(39) & convTransposeA_CP_3995_elements(47) & convTransposeA_CP_3995_elements(53) & convTransposeA_CP_3995_elements(55);
      gj_convTransposeA_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3995_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	83 
    -- CP-element group 57: 	84 
    -- CP-element group 57:  members (24) 
      -- CP-element group 57: 	 branch_block_stmt_1377/if_stmt_1752_if_link/$exit
      -- CP-element group 57: 	 branch_block_stmt_1377/if_stmt_1752_if_link/if_choice_transition
      -- CP-element group 57: 	 branch_block_stmt_1377/merge_stmt_1758__exit__
      -- CP-element group 57: 	 branch_block_stmt_1377/whilex_xbody_ifx_xthen
      -- CP-element group 57: 	 branch_block_stmt_1377/assign_stmt_1764__entry__
      -- CP-element group 57: 	 branch_block_stmt_1377/assign_stmt_1764__exit__
      -- CP-element group 57: 	 branch_block_stmt_1377/ifx_xthen_whilex_xbody
      -- CP-element group 57: 	 branch_block_stmt_1377/assign_stmt_1764/$entry
      -- CP-element group 57: 	 branch_block_stmt_1377/assign_stmt_1764/$exit
      -- CP-element group 57: 	 branch_block_stmt_1377/ifx_xthen_whilex_xbody_PhiReq/$entry
      -- CP-element group 57: 	 branch_block_stmt_1377/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1645/$entry
      -- CP-element group 57: 	 branch_block_stmt_1377/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1645/phi_stmt_1645_sources/$entry
      -- CP-element group 57: 	 branch_block_stmt_1377/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1645/phi_stmt_1645_sources/type_cast_1651/$entry
      -- CP-element group 57: 	 branch_block_stmt_1377/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1645/phi_stmt_1645_sources/type_cast_1651/SplitProtocol/$entry
      -- CP-element group 57: 	 branch_block_stmt_1377/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1645/phi_stmt_1645_sources/type_cast_1651/SplitProtocol/Sample/$entry
      -- CP-element group 57: 	 branch_block_stmt_1377/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1645/phi_stmt_1645_sources/type_cast_1651/SplitProtocol/Sample/rr
      -- CP-element group 57: 	 branch_block_stmt_1377/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1645/phi_stmt_1645_sources/type_cast_1651/SplitProtocol/Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_1377/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1645/phi_stmt_1645_sources/type_cast_1651/SplitProtocol/Update/cr
      -- CP-element group 57: 	 branch_block_stmt_1377/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 57: 	 branch_block_stmt_1377/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 57: 	 branch_block_stmt_1377/merge_stmt_1758_PhiReqMerge
      -- CP-element group 57: 	 branch_block_stmt_1377/merge_stmt_1758_PhiAck/$entry
      -- CP-element group 57: 	 branch_block_stmt_1377/merge_stmt_1758_PhiAck/$exit
      -- CP-element group 57: 	 branch_block_stmt_1377/merge_stmt_1758_PhiAck/dummy
      -- 
    if_choice_transition_4872_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1752_branch_ack_1, ack => convTransposeA_CP_3995_elements(57)); -- 
    rr_5055_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5055_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(57), ack => type_cast_1651_inst_req_0); -- 
    cr_5060_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5060_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(57), ack => type_cast_1651_inst_req_1); -- 
    -- CP-element group 58:  fork  transition  place  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	56 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58: 	60 
    -- CP-element group 58: 	62 
    -- CP-element group 58: 	64 
    -- CP-element group 58:  members (24) 
      -- CP-element group 58: 	 branch_block_stmt_1377/whilex_xbody_ifx_xelse
      -- CP-element group 58: 	 branch_block_stmt_1377/if_stmt_1752_else_link/$exit
      -- CP-element group 58: 	 branch_block_stmt_1377/merge_stmt_1766__exit__
      -- CP-element group 58: 	 branch_block_stmt_1377/assign_stmt_1772_to_assign_stmt_1808__entry__
      -- CP-element group 58: 	 branch_block_stmt_1377/if_stmt_1752_else_link/else_choice_transition
      -- CP-element group 58: 	 branch_block_stmt_1377/assign_stmt_1772_to_assign_stmt_1808/$entry
      -- CP-element group 58: 	 branch_block_stmt_1377/assign_stmt_1772_to_assign_stmt_1808/type_cast_1776_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_1377/assign_stmt_1772_to_assign_stmt_1808/type_cast_1776_update_start_
      -- CP-element group 58: 	 branch_block_stmt_1377/assign_stmt_1772_to_assign_stmt_1808/type_cast_1776_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_1377/assign_stmt_1772_to_assign_stmt_1808/type_cast_1776_Sample/rr
      -- CP-element group 58: 	 branch_block_stmt_1377/assign_stmt_1772_to_assign_stmt_1808/type_cast_1776_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_1377/assign_stmt_1772_to_assign_stmt_1808/type_cast_1776_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_1377/assign_stmt_1772_to_assign_stmt_1808/type_cast_1785_update_start_
      -- CP-element group 58: 	 branch_block_stmt_1377/assign_stmt_1772_to_assign_stmt_1808/type_cast_1785_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_1377/assign_stmt_1772_to_assign_stmt_1808/type_cast_1785_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_1377/assign_stmt_1772_to_assign_stmt_1808/type_cast_1802_update_start_
      -- CP-element group 58: 	 branch_block_stmt_1377/assign_stmt_1772_to_assign_stmt_1808/type_cast_1802_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_1377/assign_stmt_1772_to_assign_stmt_1808/type_cast_1802_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_1377/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 58: 	 branch_block_stmt_1377/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 58: 	 branch_block_stmt_1377/merge_stmt_1766_PhiReqMerge
      -- CP-element group 58: 	 branch_block_stmt_1377/merge_stmt_1766_PhiAck/$entry
      -- CP-element group 58: 	 branch_block_stmt_1377/merge_stmt_1766_PhiAck/$exit
      -- CP-element group 58: 	 branch_block_stmt_1377/merge_stmt_1766_PhiAck/dummy
      -- 
    else_choice_transition_4876_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1752_branch_ack_0, ack => convTransposeA_CP_3995_elements(58)); -- 
    rr_4892_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4892_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(58), ack => type_cast_1776_inst_req_0); -- 
    cr_4897_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4897_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(58), ack => type_cast_1776_inst_req_1); -- 
    cr_4911_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4911_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(58), ack => type_cast_1785_inst_req_1); -- 
    cr_4925_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4925_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(58), ack => type_cast_1802_inst_req_1); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_1377/assign_stmt_1772_to_assign_stmt_1808/type_cast_1776_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_1377/assign_stmt_1772_to_assign_stmt_1808/type_cast_1776_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_1377/assign_stmt_1772_to_assign_stmt_1808/type_cast_1776_Sample/ra
      -- 
    ra_4893_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1776_inst_ack_0, ack => convTransposeA_CP_3995_elements(59)); -- 
    -- CP-element group 60:  transition  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	58 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (6) 
      -- CP-element group 60: 	 branch_block_stmt_1377/assign_stmt_1772_to_assign_stmt_1808/type_cast_1776_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_1377/assign_stmt_1772_to_assign_stmt_1808/type_cast_1776_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_1377/assign_stmt_1772_to_assign_stmt_1808/type_cast_1776_Update/ca
      -- CP-element group 60: 	 branch_block_stmt_1377/assign_stmt_1772_to_assign_stmt_1808/type_cast_1785_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_1377/assign_stmt_1772_to_assign_stmt_1808/type_cast_1785_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_1377/assign_stmt_1772_to_assign_stmt_1808/type_cast_1785_Sample/rr
      -- 
    ca_4898_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1776_inst_ack_1, ack => convTransposeA_CP_3995_elements(60)); -- 
    rr_4906_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4906_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(60), ack => type_cast_1785_inst_req_0); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_1377/assign_stmt_1772_to_assign_stmt_1808/type_cast_1785_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_1377/assign_stmt_1772_to_assign_stmt_1808/type_cast_1785_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_1377/assign_stmt_1772_to_assign_stmt_1808/type_cast_1785_Sample/ra
      -- 
    ra_4907_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1785_inst_ack_0, ack => convTransposeA_CP_3995_elements(61)); -- 
    -- CP-element group 62:  transition  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	58 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (6) 
      -- CP-element group 62: 	 branch_block_stmt_1377/assign_stmt_1772_to_assign_stmt_1808/type_cast_1785_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_1377/assign_stmt_1772_to_assign_stmt_1808/type_cast_1785_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_1377/assign_stmt_1772_to_assign_stmt_1808/type_cast_1785_Update/ca
      -- CP-element group 62: 	 branch_block_stmt_1377/assign_stmt_1772_to_assign_stmt_1808/type_cast_1802_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_1377/assign_stmt_1772_to_assign_stmt_1808/type_cast_1802_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_1377/assign_stmt_1772_to_assign_stmt_1808/type_cast_1802_Sample/rr
      -- 
    ca_4912_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1785_inst_ack_1, ack => convTransposeA_CP_3995_elements(62)); -- 
    rr_4920_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4920_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(62), ack => type_cast_1802_inst_req_0); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_1377/assign_stmt_1772_to_assign_stmt_1808/type_cast_1802_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_1377/assign_stmt_1772_to_assign_stmt_1808/type_cast_1802_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_1377/assign_stmt_1772_to_assign_stmt_1808/type_cast_1802_Sample/ra
      -- 
    ra_4921_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1802_inst_ack_0, ack => convTransposeA_CP_3995_elements(63)); -- 
    -- CP-element group 64:  branch  transition  place  input  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	58 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64: 	66 
    -- CP-element group 64:  members (13) 
      -- CP-element group 64: 	 branch_block_stmt_1377/R_cmp77_1810_place
      -- CP-element group 64: 	 branch_block_stmt_1377/assign_stmt_1772_to_assign_stmt_1808__exit__
      -- CP-element group 64: 	 branch_block_stmt_1377/if_stmt_1809__entry__
      -- CP-element group 64: 	 branch_block_stmt_1377/assign_stmt_1772_to_assign_stmt_1808/$exit
      -- CP-element group 64: 	 branch_block_stmt_1377/assign_stmt_1772_to_assign_stmt_1808/type_cast_1802_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_1377/assign_stmt_1772_to_assign_stmt_1808/type_cast_1802_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_1377/assign_stmt_1772_to_assign_stmt_1808/type_cast_1802_Update/ca
      -- CP-element group 64: 	 branch_block_stmt_1377/if_stmt_1809_dead_link/$entry
      -- CP-element group 64: 	 branch_block_stmt_1377/if_stmt_1809_eval_test/$entry
      -- CP-element group 64: 	 branch_block_stmt_1377/if_stmt_1809_eval_test/$exit
      -- CP-element group 64: 	 branch_block_stmt_1377/if_stmt_1809_eval_test/branch_req
      -- CP-element group 64: 	 branch_block_stmt_1377/if_stmt_1809_if_link/$entry
      -- CP-element group 64: 	 branch_block_stmt_1377/if_stmt_1809_else_link/$entry
      -- 
    ca_4926_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1802_inst_ack_1, ack => convTransposeA_CP_3995_elements(64)); -- 
    branch_req_4934_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4934_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(64), ack => if_stmt_1809_branch_req_0); -- 
    -- CP-element group 65:  merge  transition  place  input  output  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	67 
    -- CP-element group 65:  members (15) 
      -- CP-element group 65: 	 branch_block_stmt_1377/ifx_xelse_whilex_xend
      -- CP-element group 65: 	 branch_block_stmt_1377/merge_stmt_1815__exit__
      -- CP-element group 65: 	 branch_block_stmt_1377/assign_stmt_1819__entry__
      -- CP-element group 65: 	 branch_block_stmt_1377/if_stmt_1809_if_link/$exit
      -- CP-element group 65: 	 branch_block_stmt_1377/if_stmt_1809_if_link/if_choice_transition
      -- CP-element group 65: 	 branch_block_stmt_1377/assign_stmt_1819/$entry
      -- CP-element group 65: 	 branch_block_stmt_1377/assign_stmt_1819/WPIPE_Block0_done_1817_sample_start_
      -- CP-element group 65: 	 branch_block_stmt_1377/assign_stmt_1819/WPIPE_Block0_done_1817_Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_1377/assign_stmt_1819/WPIPE_Block0_done_1817_Sample/req
      -- CP-element group 65: 	 branch_block_stmt_1377/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 65: 	 branch_block_stmt_1377/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 65: 	 branch_block_stmt_1377/merge_stmt_1815_PhiReqMerge
      -- CP-element group 65: 	 branch_block_stmt_1377/merge_stmt_1815_PhiAck/$entry
      -- CP-element group 65: 	 branch_block_stmt_1377/merge_stmt_1815_PhiAck/$exit
      -- CP-element group 65: 	 branch_block_stmt_1377/merge_stmt_1815_PhiAck/dummy
      -- 
    if_choice_transition_4939_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1809_branch_ack_1, ack => convTransposeA_CP_3995_elements(65)); -- 
    req_4956_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4956_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(65), ack => WPIPE_Block0_done_1817_inst_req_0); -- 
    -- CP-element group 66:  fork  transition  place  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	64 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	72 
    -- CP-element group 66: 	73 
    -- CP-element group 66: 	75 
    -- CP-element group 66: 	76 
    -- CP-element group 66:  members (20) 
      -- CP-element group 66: 	 branch_block_stmt_1377/ifx_xelse_whilex_xbodyx_xouter
      -- CP-element group 66: 	 branch_block_stmt_1377/if_stmt_1809_else_link/$exit
      -- CP-element group 66: 	 branch_block_stmt_1377/if_stmt_1809_else_link/else_choice_transition
      -- CP-element group 66: 	 branch_block_stmt_1377/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 66: 	 branch_block_stmt_1377/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1515/$entry
      -- CP-element group 66: 	 branch_block_stmt_1377/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1515/phi_stmt_1515_sources/$entry
      -- CP-element group 66: 	 branch_block_stmt_1377/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1515/phi_stmt_1515_sources/type_cast_1521/$entry
      -- CP-element group 66: 	 branch_block_stmt_1377/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1515/phi_stmt_1515_sources/type_cast_1521/SplitProtocol/$entry
      -- CP-element group 66: 	 branch_block_stmt_1377/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1515/phi_stmt_1515_sources/type_cast_1521/SplitProtocol/Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_1377/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1515/phi_stmt_1515_sources/type_cast_1521/SplitProtocol/Sample/rr
      -- CP-element group 66: 	 branch_block_stmt_1377/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1515/phi_stmt_1515_sources/type_cast_1521/SplitProtocol/Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_1377/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1515/phi_stmt_1515_sources/type_cast_1521/SplitProtocol/Update/cr
      -- CP-element group 66: 	 branch_block_stmt_1377/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1522/$entry
      -- CP-element group 66: 	 branch_block_stmt_1377/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1522/phi_stmt_1522_sources/$entry
      -- CP-element group 66: 	 branch_block_stmt_1377/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1522/phi_stmt_1522_sources/type_cast_1528/$entry
      -- CP-element group 66: 	 branch_block_stmt_1377/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1522/phi_stmt_1522_sources/type_cast_1528/SplitProtocol/$entry
      -- CP-element group 66: 	 branch_block_stmt_1377/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1522/phi_stmt_1522_sources/type_cast_1528/SplitProtocol/Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_1377/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1522/phi_stmt_1522_sources/type_cast_1528/SplitProtocol/Sample/rr
      -- CP-element group 66: 	 branch_block_stmt_1377/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1522/phi_stmt_1522_sources/type_cast_1528/SplitProtocol/Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_1377/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1522/phi_stmt_1522_sources/type_cast_1528/SplitProtocol/Update/cr
      -- 
    else_choice_transition_4943_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1809_branch_ack_0, ack => convTransposeA_CP_3995_elements(66)); -- 
    rr_5000_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5000_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(66), ack => type_cast_1521_inst_req_0); -- 
    cr_5005_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5005_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(66), ack => type_cast_1521_inst_req_1); -- 
    rr_5023_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5023_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(66), ack => type_cast_1528_inst_req_0); -- 
    cr_5028_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5028_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(66), ack => type_cast_1528_inst_req_1); -- 
    -- CP-element group 67:  transition  input  output  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	65 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (6) 
      -- CP-element group 67: 	 branch_block_stmt_1377/assign_stmt_1819/WPIPE_Block0_done_1817_sample_completed_
      -- CP-element group 67: 	 branch_block_stmt_1377/assign_stmt_1819/WPIPE_Block0_done_1817_update_start_
      -- CP-element group 67: 	 branch_block_stmt_1377/assign_stmt_1819/WPIPE_Block0_done_1817_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_1377/assign_stmt_1819/WPIPE_Block0_done_1817_Sample/ack
      -- CP-element group 67: 	 branch_block_stmt_1377/assign_stmt_1819/WPIPE_Block0_done_1817_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_1377/assign_stmt_1819/WPIPE_Block0_done_1817_Update/req
      -- 
    ack_4957_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_done_1817_inst_ack_0, ack => convTransposeA_CP_3995_elements(67)); -- 
    req_4961_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4961_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(67), ack => WPIPE_Block0_done_1817_inst_req_1); -- 
    -- CP-element group 68:  transition  place  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (16) 
      -- CP-element group 68: 	 $exit
      -- CP-element group 68: 	 branch_block_stmt_1377/$exit
      -- CP-element group 68: 	 branch_block_stmt_1377/branch_block_stmt_1377__exit__
      -- CP-element group 68: 	 branch_block_stmt_1377/assign_stmt_1819__exit__
      -- CP-element group 68: 	 branch_block_stmt_1377/return__
      -- CP-element group 68: 	 branch_block_stmt_1377/merge_stmt_1821__exit__
      -- CP-element group 68: 	 branch_block_stmt_1377/assign_stmt_1819/$exit
      -- CP-element group 68: 	 branch_block_stmt_1377/assign_stmt_1819/WPIPE_Block0_done_1817_update_completed_
      -- CP-element group 68: 	 branch_block_stmt_1377/assign_stmt_1819/WPIPE_Block0_done_1817_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_1377/assign_stmt_1819/WPIPE_Block0_done_1817_Update/ack
      -- CP-element group 68: 	 branch_block_stmt_1377/return___PhiReq/$entry
      -- CP-element group 68: 	 branch_block_stmt_1377/return___PhiReq/$exit
      -- CP-element group 68: 	 branch_block_stmt_1377/merge_stmt_1821_PhiReqMerge
      -- CP-element group 68: 	 branch_block_stmt_1377/merge_stmt_1821_PhiAck/$entry
      -- CP-element group 68: 	 branch_block_stmt_1377/merge_stmt_1821_PhiAck/$exit
      -- CP-element group 68: 	 branch_block_stmt_1377/merge_stmt_1821_PhiAck/dummy
      -- 
    ack_4962_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_done_1817_inst_ack_1, ack => convTransposeA_CP_3995_elements(68)); -- 
    -- CP-element group 69:  transition  output  delay-element  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	29 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	71 
    -- CP-element group 69:  members (4) 
      -- CP-element group 69: 	 branch_block_stmt_1377/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1515/$exit
      -- CP-element group 69: 	 branch_block_stmt_1377/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1515/phi_stmt_1515_sources/$exit
      -- CP-element group 69: 	 branch_block_stmt_1377/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1515/phi_stmt_1515_sources/type_cast_1519_konst_delay_trans
      -- CP-element group 69: 	 branch_block_stmt_1377/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1515/phi_stmt_1515_req
      -- 
    phi_stmt_1515_req_4973_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1515_req_4973_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(69), ack => phi_stmt_1515_req_0); -- 
    -- Element group convTransposeA_CP_3995_elements(69) is a control-delay.
    cp_element_69_delay: control_delay_element  generic map(name => " 69_delay", delay_value => 1)  port map(req => convTransposeA_CP_3995_elements(29), ack => convTransposeA_CP_3995_elements(69), clk => clk, reset =>reset);
    -- CP-element group 70:  transition  output  delay-element  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	29 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70:  members (4) 
      -- CP-element group 70: 	 branch_block_stmt_1377/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1522/$exit
      -- CP-element group 70: 	 branch_block_stmt_1377/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1522/phi_stmt_1522_sources/$exit
      -- CP-element group 70: 	 branch_block_stmt_1377/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1522/phi_stmt_1522_sources/type_cast_1526_konst_delay_trans
      -- CP-element group 70: 	 branch_block_stmt_1377/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1522/phi_stmt_1522_req
      -- 
    phi_stmt_1522_req_4981_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1522_req_4981_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(70), ack => phi_stmt_1522_req_0); -- 
    -- Element group convTransposeA_CP_3995_elements(70) is a control-delay.
    cp_element_70_delay: control_delay_element  generic map(name => " 70_delay", delay_value => 1)  port map(req => convTransposeA_CP_3995_elements(29), ack => convTransposeA_CP_3995_elements(70), clk => clk, reset =>reset);
    -- CP-element group 71:  join  transition  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	69 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	79 
    -- CP-element group 71:  members (1) 
      -- CP-element group 71: 	 branch_block_stmt_1377/entry_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3995_elements(69) & convTransposeA_CP_3995_elements(70);
      gj_convTransposeA_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3995_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	66 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	74 
    -- CP-element group 72:  members (2) 
      -- CP-element group 72: 	 branch_block_stmt_1377/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1515/phi_stmt_1515_sources/type_cast_1521/SplitProtocol/Sample/$exit
      -- CP-element group 72: 	 branch_block_stmt_1377/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1515/phi_stmt_1515_sources/type_cast_1521/SplitProtocol/Sample/ra
      -- 
    ra_5001_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1521_inst_ack_0, ack => convTransposeA_CP_3995_elements(72)); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	66 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (2) 
      -- CP-element group 73: 	 branch_block_stmt_1377/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1515/phi_stmt_1515_sources/type_cast_1521/SplitProtocol/Update/$exit
      -- CP-element group 73: 	 branch_block_stmt_1377/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1515/phi_stmt_1515_sources/type_cast_1521/SplitProtocol/Update/ca
      -- 
    ca_5006_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1521_inst_ack_1, ack => convTransposeA_CP_3995_elements(73)); -- 
    -- CP-element group 74:  join  transition  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	72 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	78 
    -- CP-element group 74:  members (5) 
      -- CP-element group 74: 	 branch_block_stmt_1377/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1515/$exit
      -- CP-element group 74: 	 branch_block_stmt_1377/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1515/phi_stmt_1515_sources/$exit
      -- CP-element group 74: 	 branch_block_stmt_1377/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1515/phi_stmt_1515_sources/type_cast_1521/$exit
      -- CP-element group 74: 	 branch_block_stmt_1377/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1515/phi_stmt_1515_sources/type_cast_1521/SplitProtocol/$exit
      -- CP-element group 74: 	 branch_block_stmt_1377/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1515/phi_stmt_1515_req
      -- 
    phi_stmt_1515_req_5007_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1515_req_5007_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(74), ack => phi_stmt_1515_req_1); -- 
    convTransposeA_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3995_elements(72) & convTransposeA_CP_3995_elements(73);
      gj_convTransposeA_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3995_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	66 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (2) 
      -- CP-element group 75: 	 branch_block_stmt_1377/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1522/phi_stmt_1522_sources/type_cast_1528/SplitProtocol/Sample/$exit
      -- CP-element group 75: 	 branch_block_stmt_1377/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1522/phi_stmt_1522_sources/type_cast_1528/SplitProtocol/Sample/ra
      -- 
    ra_5024_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1528_inst_ack_0, ack => convTransposeA_CP_3995_elements(75)); -- 
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	66 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76:  members (2) 
      -- CP-element group 76: 	 branch_block_stmt_1377/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1522/phi_stmt_1522_sources/type_cast_1528/SplitProtocol/Update/$exit
      -- CP-element group 76: 	 branch_block_stmt_1377/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1522/phi_stmt_1522_sources/type_cast_1528/SplitProtocol/Update/ca
      -- 
    ca_5029_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1528_inst_ack_1, ack => convTransposeA_CP_3995_elements(76)); -- 
    -- CP-element group 77:  join  transition  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: 	76 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (5) 
      -- CP-element group 77: 	 branch_block_stmt_1377/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1522/$exit
      -- CP-element group 77: 	 branch_block_stmt_1377/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1522/phi_stmt_1522_sources/$exit
      -- CP-element group 77: 	 branch_block_stmt_1377/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1522/phi_stmt_1522_sources/type_cast_1528/$exit
      -- CP-element group 77: 	 branch_block_stmt_1377/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1522/phi_stmt_1522_sources/type_cast_1528/SplitProtocol/$exit
      -- CP-element group 77: 	 branch_block_stmt_1377/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1522/phi_stmt_1522_req
      -- 
    phi_stmt_1522_req_5030_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1522_req_5030_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(77), ack => phi_stmt_1522_req_1); -- 
    convTransposeA_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3995_elements(75) & convTransposeA_CP_3995_elements(76);
      gj_convTransposeA_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3995_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  join  transition  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	74 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_1377/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_78: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_78"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3995_elements(74) & convTransposeA_CP_3995_elements(77);
      gj_convTransposeA_cp_element_group_78 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3995_elements(78), clk => clk, reset => reset); --
    end block;
    -- CP-element group 79:  merge  fork  transition  place  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	71 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79: 	81 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_1377/merge_stmt_1514_PhiReqMerge
      -- CP-element group 79: 	 branch_block_stmt_1377/merge_stmt_1514_PhiAck/$entry
      -- 
    convTransposeA_CP_3995_elements(79) <= OrReduce(convTransposeA_CP_3995_elements(71) & convTransposeA_CP_3995_elements(78));
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	82 
    -- CP-element group 80:  members (1) 
      -- CP-element group 80: 	 branch_block_stmt_1377/merge_stmt_1514_PhiAck/phi_stmt_1515_ack
      -- 
    phi_stmt_1515_ack_5035_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1515_ack_0, ack => convTransposeA_CP_3995_elements(80)); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	79 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	82 
    -- CP-element group 81:  members (1) 
      -- CP-element group 81: 	 branch_block_stmt_1377/merge_stmt_1514_PhiAck/phi_stmt_1522_ack
      -- 
    phi_stmt_1522_ack_5036_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1522_ack_0, ack => convTransposeA_CP_3995_elements(81)); -- 
    -- CP-element group 82:  join  fork  transition  place  output  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	80 
    -- CP-element group 82: 	81 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	30 
    -- CP-element group 82: 	31 
    -- CP-element group 82: 	32 
    -- CP-element group 82: 	33 
    -- CP-element group 82:  members (16) 
      -- CP-element group 82: 	 branch_block_stmt_1377/assign_stmt_1535_to_assign_stmt_1642/type_cast_1539_update_start_
      -- CP-element group 82: 	 branch_block_stmt_1377/assign_stmt_1535_to_assign_stmt_1642/type_cast_1539_sample_start_
      -- CP-element group 82: 	 branch_block_stmt_1377/merge_stmt_1514__exit__
      -- CP-element group 82: 	 branch_block_stmt_1377/assign_stmt_1535_to_assign_stmt_1642__entry__
      -- CP-element group 82: 	 branch_block_stmt_1377/assign_stmt_1535_to_assign_stmt_1642/type_cast_1534_Update/cr
      -- CP-element group 82: 	 branch_block_stmt_1377/assign_stmt_1535_to_assign_stmt_1642/type_cast_1534_Update/$entry
      -- CP-element group 82: 	 branch_block_stmt_1377/assign_stmt_1535_to_assign_stmt_1642/type_cast_1534_Sample/rr
      -- CP-element group 82: 	 branch_block_stmt_1377/assign_stmt_1535_to_assign_stmt_1642/type_cast_1534_Sample/$entry
      -- CP-element group 82: 	 branch_block_stmt_1377/assign_stmt_1535_to_assign_stmt_1642/type_cast_1534_update_start_
      -- CP-element group 82: 	 branch_block_stmt_1377/assign_stmt_1535_to_assign_stmt_1642/type_cast_1534_sample_start_
      -- CP-element group 82: 	 branch_block_stmt_1377/assign_stmt_1535_to_assign_stmt_1642/$entry
      -- CP-element group 82: 	 branch_block_stmt_1377/assign_stmt_1535_to_assign_stmt_1642/type_cast_1539_Update/cr
      -- CP-element group 82: 	 branch_block_stmt_1377/assign_stmt_1535_to_assign_stmt_1642/type_cast_1539_Update/$entry
      -- CP-element group 82: 	 branch_block_stmt_1377/assign_stmt_1535_to_assign_stmt_1642/type_cast_1539_Sample/rr
      -- CP-element group 82: 	 branch_block_stmt_1377/assign_stmt_1535_to_assign_stmt_1642/type_cast_1539_Sample/$entry
      -- CP-element group 82: 	 branch_block_stmt_1377/merge_stmt_1514_PhiAck/$exit
      -- 
    cr_4593_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4593_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(82), ack => type_cast_1534_inst_req_1); -- 
    rr_4588_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4588_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(82), ack => type_cast_1534_inst_req_0); -- 
    cr_4607_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4607_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(82), ack => type_cast_1539_inst_req_1); -- 
    rr_4602_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4602_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(82), ack => type_cast_1539_inst_req_0); -- 
    convTransposeA_cp_element_group_82: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_82"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3995_elements(80) & convTransposeA_CP_3995_elements(81);
      gj_convTransposeA_cp_element_group_82 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3995_elements(82), clk => clk, reset => reset); --
    end block;
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	57 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	85 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_1377/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1645/phi_stmt_1645_sources/type_cast_1651/SplitProtocol/Sample/$exit
      -- CP-element group 83: 	 branch_block_stmt_1377/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1645/phi_stmt_1645_sources/type_cast_1651/SplitProtocol/Sample/ra
      -- 
    ra_5056_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1651_inst_ack_0, ack => convTransposeA_CP_3995_elements(83)); -- 
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	57 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84:  members (2) 
      -- CP-element group 84: 	 branch_block_stmt_1377/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1645/phi_stmt_1645_sources/type_cast_1651/SplitProtocol/Update/$exit
      -- CP-element group 84: 	 branch_block_stmt_1377/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1645/phi_stmt_1645_sources/type_cast_1651/SplitProtocol/Update/ca
      -- 
    ca_5061_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1651_inst_ack_1, ack => convTransposeA_CP_3995_elements(84)); -- 
    -- CP-element group 85:  join  transition  output  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	83 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (6) 
      -- CP-element group 85: 	 branch_block_stmt_1377/ifx_xthen_whilex_xbody_PhiReq/$exit
      -- CP-element group 85: 	 branch_block_stmt_1377/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1645/$exit
      -- CP-element group 85: 	 branch_block_stmt_1377/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1645/phi_stmt_1645_sources/$exit
      -- CP-element group 85: 	 branch_block_stmt_1377/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1645/phi_stmt_1645_sources/type_cast_1651/$exit
      -- CP-element group 85: 	 branch_block_stmt_1377/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1645/phi_stmt_1645_sources/type_cast_1651/SplitProtocol/$exit
      -- CP-element group 85: 	 branch_block_stmt_1377/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1645/phi_stmt_1645_req
      -- 
    phi_stmt_1645_req_5062_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1645_req_5062_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(85), ack => phi_stmt_1645_req_1); -- 
    convTransposeA_cp_element_group_85: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_85"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_3995_elements(83) & convTransposeA_CP_3995_elements(84);
      gj_convTransposeA_cp_element_group_85 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_3995_elements(85), clk => clk, reset => reset); --
    end block;
    -- CP-element group 86:  transition  output  delay-element  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	34 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (5) 
      -- CP-element group 86: 	 branch_block_stmt_1377/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$exit
      -- CP-element group 86: 	 branch_block_stmt_1377/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1645/$exit
      -- CP-element group 86: 	 branch_block_stmt_1377/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1645/phi_stmt_1645_sources/$exit
      -- CP-element group 86: 	 branch_block_stmt_1377/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1645/phi_stmt_1645_sources/type_cast_1649_konst_delay_trans
      -- CP-element group 86: 	 branch_block_stmt_1377/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1645/phi_stmt_1645_req
      -- 
    phi_stmt_1645_req_5073_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1645_req_5073_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(86), ack => phi_stmt_1645_req_0); -- 
    -- Element group convTransposeA_CP_3995_elements(86) is a control-delay.
    cp_element_86_delay: control_delay_element  generic map(name => " 86_delay", delay_value => 1)  port map(req => convTransposeA_CP_3995_elements(34), ack => convTransposeA_CP_3995_elements(86), clk => clk, reset =>reset);
    -- CP-element group 87:  merge  transition  place  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (2) 
      -- CP-element group 87: 	 branch_block_stmt_1377/merge_stmt_1644_PhiReqMerge
      -- CP-element group 87: 	 branch_block_stmt_1377/merge_stmt_1644_PhiAck/$entry
      -- 
    convTransposeA_CP_3995_elements(87) <= OrReduce(convTransposeA_CP_3995_elements(85) & convTransposeA_CP_3995_elements(86));
    -- CP-element group 88:  fork  transition  place  input  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	35 
    -- CP-element group 88: 	36 
    -- CP-element group 88: 	38 
    -- CP-element group 88: 	40 
    -- CP-element group 88: 	42 
    -- CP-element group 88: 	44 
    -- CP-element group 88: 	46 
    -- CP-element group 88: 	48 
    -- CP-element group 88: 	50 
    -- CP-element group 88: 	53 
    -- CP-element group 88: 	54 
    -- CP-element group 88: 	55 
    -- CP-element group 88:  members (45) 
      -- CP-element group 88: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/array_obj_ref_1729_final_index_sum_regn_Update/req
      -- CP-element group 88: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/array_obj_ref_1698_final_index_sum_regn_update_start
      -- CP-element group 88: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/type_cast_1723_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1703_Update/word_access_complete/word_0/cr
      -- CP-element group 88: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/array_obj_ref_1729_final_index_sum_regn_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1703_Update/word_access_complete/word_0/$entry
      -- CP-element group 88: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/array_obj_ref_1698_final_index_sum_regn_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1733_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/type_cast_1739_Sample/rr
      -- CP-element group 88: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/type_cast_1739_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/type_cast_1739_Update/cr
      -- CP-element group 88: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/type_cast_1739_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1733_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/array_obj_ref_1729_final_index_sum_regn_update_start
      -- CP-element group 88: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1733_Update/word_access_complete/word_0/cr
      -- CP-element group 88: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/type_cast_1739_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1733_Update/word_access_complete/word_0/$entry
      -- CP-element group 88: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1703_Update/word_access_complete/$entry
      -- CP-element group 88: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1733_Update/word_access_complete/$entry
      -- CP-element group 88: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/type_cast_1739_Sample/$entry
      -- CP-element group 88: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/addr_of_1730_complete/req
      -- CP-element group 88: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/addr_of_1730_complete/$entry
      -- CP-element group 88: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/array_obj_ref_1698_final_index_sum_regn_Update/req
      -- CP-element group 88: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/addr_of_1730_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1377/merge_stmt_1644__exit__
      -- CP-element group 88: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751__entry__
      -- CP-element group 88: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1703_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/type_cast_1723_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/addr_of_1699_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/type_cast_1692_Update/cr
      -- CP-element group 88: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/type_cast_1692_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/ptr_deref_1703_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/type_cast_1692_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/type_cast_1661_Update/cr
      -- CP-element group 88: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/type_cast_1661_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/type_cast_1661_Sample/rr
      -- CP-element group 88: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/addr_of_1699_complete/req
      -- CP-element group 88: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/type_cast_1661_Sample/$entry
      -- CP-element group 88: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/type_cast_1661_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/addr_of_1699_complete/$entry
      -- CP-element group 88: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/type_cast_1661_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/$entry
      -- CP-element group 88: 	 branch_block_stmt_1377/assign_stmt_1658_to_assign_stmt_1751/type_cast_1723_Update/cr
      -- CP-element group 88: 	 branch_block_stmt_1377/merge_stmt_1644_PhiAck/$exit
      -- CP-element group 88: 	 branch_block_stmt_1377/merge_stmt_1644_PhiAck/phi_stmt_1645_ack
      -- 
    phi_stmt_1645_ack_5078_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1645_ack_0, ack => convTransposeA_CP_3995_elements(88)); -- 
    req_4779_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4779_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(88), ack => array_obj_ref_1729_index_offset_req_1); -- 
    cr_4729_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4729_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(88), ack => ptr_deref_1703_load_0_req_1); -- 
    rr_4853_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4853_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(88), ack => type_cast_1739_inst_req_0); -- 
    cr_4858_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4858_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(88), ack => type_cast_1739_inst_req_1); -- 
    cr_4844_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4844_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(88), ack => ptr_deref_1733_store_0_req_1); -- 
    req_4794_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4794_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(88), ack => addr_of_1730_final_reg_req_1); -- 
    req_4669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(88), ack => array_obj_ref_1698_index_offset_req_1); -- 
    cr_4638_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4638_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(88), ack => type_cast_1692_inst_req_1); -- 
    cr_4624_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4624_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(88), ack => type_cast_1661_inst_req_1); -- 
    rr_4619_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4619_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(88), ack => type_cast_1661_inst_req_0); -- 
    req_4684_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4684_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(88), ack => addr_of_1699_final_reg_req_1); -- 
    cr_4748_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4748_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_3995_elements(88), ack => type_cast_1723_inst_req_1); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i32_i32_1604_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1625_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1685_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1717_wire : std_logic_vector(31 downto 0);
    signal LOAD_padding_1433_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_padding_1433_word_address_0 : std_logic_vector(0 downto 0);
    signal R_idxprom52_1728_resized : std_logic_vector(13 downto 0);
    signal R_idxprom52_1728_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_1697_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_1697_scaled : std_logic_vector(13 downto 0);
    signal add16_1565 : std_logic_vector(31 downto 0);
    signal add27_1580 : std_logic_vector(31 downto 0);
    signal add42_1637 : std_logic_vector(31 downto 0);
    signal add44_1672 : std_logic_vector(31 downto 0);
    signal add57_1746 : std_logic_vector(31 downto 0);
    signal add8_1667 : std_logic_vector(31 downto 0);
    signal add_1550 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1698_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1698_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1698_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1698_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1698_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1698_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1729_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1729_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1729_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1729_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1729_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1729_root_address : std_logic_vector(13 downto 0);
    signal arrayidx53_1731 : std_logic_vector(31 downto 0);
    signal arrayidx_1700 : std_logic_vector(31 downto 0);
    signal call_1380 : std_logic_vector(15 downto 0);
    signal cmp68_1782 : std_logic_vector(0 downto 0);
    signal cmp77_1808 : std_logic_vector(0 downto 0);
    signal cmp_1751 : std_logic_vector(0 downto 0);
    signal conv13_1419 : std_logic_vector(31 downto 0);
    signal conv18_1438 : std_logic_vector(31 downto 0);
    signal conv24_1452 : std_logic_vector(31 downto 0);
    signal conv37_1606 : std_logic_vector(31 downto 0);
    signal conv3_1535 : std_logic_vector(31 downto 0);
    signal conv40_1627 : std_logic_vector(31 downto 0);
    signal conv56_1740 : std_logic_vector(31 downto 0);
    signal conv66_1777 : std_logic_vector(31 downto 0);
    signal conv6_1540 : std_logic_vector(31 downto 0);
    signal conv74_1803 : std_logic_vector(31 downto 0);
    signal conv90_1662 : std_logic_vector(31 downto 0);
    signal div76_1512 : std_logic_vector(31 downto 0);
    signal div_1494 : std_logic_vector(31 downto 0);
    signal iNsTr_10_1502 : std_logic_vector(31 downto 0);
    signal iNsTr_2_1389 : std_logic_vector(31 downto 0);
    signal iNsTr_3_1401 : std_logic_vector(31 downto 0);
    signal iNsTr_4_1411 : std_logic_vector(31 downto 0);
    signal iNsTr_5_1427 : std_logic_vector(31 downto 0);
    signal iNsTr_6_1444 : std_logic_vector(31 downto 0);
    signal iNsTr_7_1460 : std_logic_vector(31 downto 0);
    signal iNsTr_8_1472 : std_logic_vector(31 downto 0);
    signal iNsTr_9_1484 : std_logic_vector(31 downto 0);
    signal idxprom52_1724 : std_logic_vector(63 downto 0);
    signal idxprom_1693 : std_logic_vector(63 downto 0);
    signal inc72_1786 : std_logic_vector(15 downto 0);
    signal inc72x_xinput_dim0x_x2_1791 : std_logic_vector(15 downto 0);
    signal inc_1772 : std_logic_vector(15 downto 0);
    signal indvar_1645 : std_logic_vector(15 downto 0);
    signal indvarx_xnext_1764 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2x_xph_1522 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1x_xph_1515 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_1798 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_1658 : std_logic_vector(15 downto 0);
    signal mul14_1560 : std_logic_vector(31 downto 0);
    signal mul25_1575 : std_logic_vector(31 downto 0);
    signal mul41_1632 : std_logic_vector(31 downto 0);
    signal mul43_1642 : std_logic_vector(31 downto 0);
    signal mul7_1555 : std_logic_vector(31 downto 0);
    signal mul_1545 : std_logic_vector(31 downto 0);
    signal ptr_deref_1392_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1392_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1392_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1392_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1392_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1404_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1404_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1404_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1404_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1404_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1414_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1414_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1414_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1414_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1414_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1430_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1430_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1430_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1430_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1430_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1447_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1447_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1447_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1447_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1447_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1463_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1463_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1463_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1463_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1463_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1475_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1475_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1475_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1475_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1475_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1487_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1487_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1487_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1487_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1487_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1505_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1505_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1505_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1505_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1505_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1703_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1703_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1703_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1703_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1703_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1733_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1733_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1733_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1733_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1733_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1733_word_offset_0 : std_logic_vector(13 downto 0);
    signal sext91_1618 : std_logic_vector(31 downto 0);
    signal sext93_1678 : std_logic_vector(31 downto 0);
    signal sext94_1710 : std_logic_vector(31 downto 0);
    signal sext_1597 : std_logic_vector(31 downto 0);
    signal shr51_1719 : std_logic_vector(31 downto 0);
    signal shr_1687 : std_logic_vector(31 downto 0);
    signal sub19_1612 : std_logic_vector(31 downto 0);
    signal sub30_1585 : std_logic_vector(31 downto 0);
    signal sub31_1591 : std_logic_vector(31 downto 0);
    signal sub_1570 : std_logic_vector(31 downto 0);
    signal tmp12_1415 : std_logic_vector(7 downto 0);
    signal tmp15_1431 : std_logic_vector(31 downto 0);
    signal tmp17_1434 : std_logic_vector(7 downto 0);
    signal tmp1_1393 : std_logic_vector(31 downto 0);
    signal tmp23_1448 : std_logic_vector(7 downto 0);
    signal tmp26_1464 : std_logic_vector(31 downto 0);
    signal tmp35_1476 : std_logic_vector(31 downto 0);
    signal tmp38_1488 : std_logic_vector(31 downto 0);
    signal tmp48_1704 : std_logic_vector(63 downto 0);
    signal tmp4_1405 : std_logic_vector(31 downto 0);
    signal tmp75_1506 : std_logic_vector(31 downto 0);
    signal type_cast_1492_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1510_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1519_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1521_wire : std_logic_vector(15 downto 0);
    signal type_cast_1526_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1528_wire : std_logic_vector(15 downto 0);
    signal type_cast_1533_wire : std_logic_vector(31 downto 0);
    signal type_cast_1538_wire : std_logic_vector(31 downto 0);
    signal type_cast_1589_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1595_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1600_wire : std_logic_vector(31 downto 0);
    signal type_cast_1603_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1610_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1616_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1621_wire : std_logic_vector(31 downto 0);
    signal type_cast_1624_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1649_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1651_wire : std_logic_vector(15 downto 0);
    signal type_cast_1656_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1676_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1681_wire : std_logic_vector(31 downto 0);
    signal type_cast_1684_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1691_wire : std_logic_vector(63 downto 0);
    signal type_cast_1708_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1713_wire : std_logic_vector(31 downto 0);
    signal type_cast_1716_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1722_wire : std_logic_vector(63 downto 0);
    signal type_cast_1738_wire : std_logic_vector(31 downto 0);
    signal type_cast_1744_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1762_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1770_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1775_wire : std_logic_vector(31 downto 0);
    signal type_cast_1795_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1801_wire : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    LOAD_padding_1433_word_address_0 <= "0";
    array_obj_ref_1698_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1698_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1698_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1698_resized_base_address <= "00000000000000";
    array_obj_ref_1729_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1729_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1729_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1729_resized_base_address <= "00000000000000";
    iNsTr_10_1502 <= "00000000000000000000000000000011";
    iNsTr_2_1389 <= "00000000000000000000000000000101";
    iNsTr_3_1401 <= "00000000000000000000000000000100";
    iNsTr_4_1411 <= "00000000000000000000000000000000";
    iNsTr_5_1427 <= "00000000000000000000000000000100";
    iNsTr_6_1444 <= "00000000000000000000000000000001";
    iNsTr_7_1460 <= "00000000000000000000000000000101";
    iNsTr_8_1472 <= "00000000000000000000000000000101";
    iNsTr_9_1484 <= "00000000000000000000000000000100";
    ptr_deref_1392_word_offset_0 <= "0000000";
    ptr_deref_1404_word_offset_0 <= "0000000";
    ptr_deref_1414_word_offset_0 <= "0";
    ptr_deref_1430_word_offset_0 <= "0000000";
    ptr_deref_1447_word_offset_0 <= "0";
    ptr_deref_1463_word_offset_0 <= "0000000";
    ptr_deref_1475_word_offset_0 <= "0000000";
    ptr_deref_1487_word_offset_0 <= "0000000";
    ptr_deref_1505_word_offset_0 <= "0000000";
    ptr_deref_1703_word_offset_0 <= "00000000000000";
    ptr_deref_1733_word_offset_0 <= "00000000000000";
    type_cast_1492_wire_constant <= "00000000000000000000000000000001";
    type_cast_1510_wire_constant <= "00000000000000000000000000000001";
    type_cast_1519_wire_constant <= "0000000000000000";
    type_cast_1526_wire_constant <= "0000000000000000";
    type_cast_1589_wire_constant <= "00000000000000000000000000010000";
    type_cast_1595_wire_constant <= "11111111111111110000000000000000";
    type_cast_1603_wire_constant <= "00000000000000000000000000010000";
    type_cast_1610_wire_constant <= "00000000000000000000000000010000";
    type_cast_1616_wire_constant <= "11111111111111110000000000000000";
    type_cast_1624_wire_constant <= "00000000000000000000000000010000";
    type_cast_1649_wire_constant <= "0000000000000000";
    type_cast_1656_wire_constant <= "0000000000000100";
    type_cast_1676_wire_constant <= "00000000000000000000000000010000";
    type_cast_1684_wire_constant <= "00000000000000000000000000010010";
    type_cast_1708_wire_constant <= "00000000000000000000000000010000";
    type_cast_1716_wire_constant <= "00000000000000000000000000010010";
    type_cast_1744_wire_constant <= "00000000000000000000000000000100";
    type_cast_1762_wire_constant <= "0000000000000001";
    type_cast_1770_wire_constant <= "0000000000000001";
    type_cast_1795_wire_constant <= "0000000000000000";
    phi_stmt_1515: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1519_wire_constant & type_cast_1521_wire;
      req <= phi_stmt_1515_req_0 & phi_stmt_1515_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1515",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1515_ack_0,
          idata => idata,
          odata => input_dim1x_x1x_xph_1515,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1515
    phi_stmt_1522: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1526_wire_constant & type_cast_1528_wire;
      req <= phi_stmt_1522_req_0 & phi_stmt_1522_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1522",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1522_ack_0,
          idata => idata,
          odata => input_dim0x_x2x_xph_1522,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1522
    phi_stmt_1645: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1649_wire_constant & type_cast_1651_wire;
      req <= phi_stmt_1645_req_0 & phi_stmt_1645_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1645",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1645_ack_0,
          idata => idata,
          odata => indvar_1645,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1645
    -- flow-through select operator MUX_1797_inst
    input_dim1x_x2_1798 <= type_cast_1795_wire_constant when (cmp68_1782(0) /=  '0') else inc_1772;
    addr_of_1699_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1699_final_reg_req_0;
      addr_of_1699_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1699_final_reg_req_1;
      addr_of_1699_final_reg_ack_1<= rack(0);
      addr_of_1699_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1699_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1698_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_1700,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1730_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1730_final_reg_req_0;
      addr_of_1730_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1730_final_reg_req_1;
      addr_of_1730_final_reg_ack_1<= rack(0);
      addr_of_1730_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1730_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1729_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx53_1731,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1418_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1418_inst_req_0;
      type_cast_1418_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1418_inst_req_1;
      type_cast_1418_inst_ack_1<= rack(0);
      type_cast_1418_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1418_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp12_1415,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv13_1419,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1437_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1437_inst_req_0;
      type_cast_1437_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1437_inst_req_1;
      type_cast_1437_inst_ack_1<= rack(0);
      type_cast_1437_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1437_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp17_1434,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv18_1438,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1451_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1451_inst_req_0;
      type_cast_1451_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1451_inst_req_1;
      type_cast_1451_inst_ack_1<= rack(0);
      type_cast_1451_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1451_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp23_1448,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv24_1452,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1521_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1521_inst_req_0;
      type_cast_1521_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1521_inst_req_1;
      type_cast_1521_inst_ack_1<= rack(0);
      type_cast_1521_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1521_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_1798,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1521_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1528_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1528_inst_req_0;
      type_cast_1528_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1528_inst_req_1;
      type_cast_1528_inst_ack_1<= rack(0);
      type_cast_1528_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1528_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc72x_xinput_dim0x_x2_1791,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1528_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1534_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1534_inst_req_0;
      type_cast_1534_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1534_inst_req_1;
      type_cast_1534_inst_ack_1<= rack(0);
      type_cast_1534_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1534_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1533_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv3_1535,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1539_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1539_inst_req_0;
      type_cast_1539_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1539_inst_req_1;
      type_cast_1539_inst_ack_1<= rack(0);
      type_cast_1539_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1539_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1538_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv6_1540,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1600_inst
    process(sext_1597) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext_1597(31 downto 0);
      type_cast_1600_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1605_inst
    process(ASHR_i32_i32_1604_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1604_wire(31 downto 0);
      conv37_1606 <= tmp_var; -- 
    end process;
    -- interlock type_cast_1621_inst
    process(sext91_1618) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext91_1618(31 downto 0);
      type_cast_1621_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1626_inst
    process(ASHR_i32_i32_1625_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1625_wire(31 downto 0);
      conv40_1627 <= tmp_var; -- 
    end process;
    type_cast_1651_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1651_inst_req_0;
      type_cast_1651_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1651_inst_req_1;
      type_cast_1651_inst_ack_1<= rack(0);
      type_cast_1651_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1651_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1764,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1651_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1661_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1661_inst_req_0;
      type_cast_1661_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1661_inst_req_1;
      type_cast_1661_inst_ack_1<= rack(0);
      type_cast_1661_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1661_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_1658,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv90_1662,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1681_inst
    process(sext93_1678) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext93_1678(31 downto 0);
      type_cast_1681_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1686_inst
    process(ASHR_i32_i32_1685_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1685_wire(31 downto 0);
      shr_1687 <= tmp_var; -- 
    end process;
    type_cast_1692_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1692_inst_req_0;
      type_cast_1692_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1692_inst_req_1;
      type_cast_1692_inst_ack_1<= rack(0);
      type_cast_1692_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1692_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1691_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_1693,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1713_inst
    process(sext94_1710) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext94_1710(31 downto 0);
      type_cast_1713_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1718_inst
    process(ASHR_i32_i32_1717_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1717_wire(31 downto 0);
      shr51_1719 <= tmp_var; -- 
    end process;
    type_cast_1723_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1723_inst_req_0;
      type_cast_1723_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1723_inst_req_1;
      type_cast_1723_inst_ack_1<= rack(0);
      type_cast_1723_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1723_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1722_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom52_1724,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1739_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1739_inst_req_0;
      type_cast_1739_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1739_inst_req_1;
      type_cast_1739_inst_ack_1<= rack(0);
      type_cast_1739_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1739_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1738_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv56_1740,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1776_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1776_inst_req_0;
      type_cast_1776_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1776_inst_req_1;
      type_cast_1776_inst_ack_1<= rack(0);
      type_cast_1776_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1776_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1775_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv66_1777,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1785_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1785_inst_req_0;
      type_cast_1785_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1785_inst_req_1;
      type_cast_1785_inst_ack_1<= rack(0);
      type_cast_1785_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1785_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp68_1782,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc72_1786,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1802_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1802_inst_req_0;
      type_cast_1802_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1802_inst_req_1;
      type_cast_1802_inst_ack_1<= rack(0);
      type_cast_1802_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1802_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1801_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv74_1803,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence LOAD_padding_1433_gather_scatter
    process(LOAD_padding_1433_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_padding_1433_data_0;
      ov(7 downto 0) := iv;
      tmp17_1434 <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1698_index_1_rename
    process(R_idxprom_1697_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_1697_resized;
      ov(13 downto 0) := iv;
      R_idxprom_1697_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1698_index_1_resize
    process(idxprom_1693) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_1693;
      ov := iv(13 downto 0);
      R_idxprom_1697_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1698_root_address_inst
    process(array_obj_ref_1698_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1698_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1698_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1729_index_1_rename
    process(R_idxprom52_1728_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom52_1728_resized;
      ov(13 downto 0) := iv;
      R_idxprom52_1728_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1729_index_1_resize
    process(idxprom52_1724) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom52_1724;
      ov := iv(13 downto 0);
      R_idxprom52_1728_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1729_root_address_inst
    process(array_obj_ref_1729_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1729_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1729_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1392_addr_0
    process(ptr_deref_1392_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1392_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1392_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1392_base_resize
    process(iNsTr_2_1389) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_2_1389;
      ov := iv(6 downto 0);
      ptr_deref_1392_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1392_gather_scatter
    process(ptr_deref_1392_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1392_data_0;
      ov(31 downto 0) := iv;
      tmp1_1393 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1392_root_address_inst
    process(ptr_deref_1392_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1392_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1392_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1404_addr_0
    process(ptr_deref_1404_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1404_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1404_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1404_base_resize
    process(iNsTr_3_1401) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_3_1401;
      ov := iv(6 downto 0);
      ptr_deref_1404_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1404_gather_scatter
    process(ptr_deref_1404_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1404_data_0;
      ov(31 downto 0) := iv;
      tmp4_1405 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1404_root_address_inst
    process(ptr_deref_1404_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1404_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1404_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1414_addr_0
    process(ptr_deref_1414_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1414_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_1414_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1414_base_resize
    process(iNsTr_4_1411) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_4_1411;
      ov := iv(0 downto 0);
      ptr_deref_1414_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1414_gather_scatter
    process(ptr_deref_1414_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1414_data_0;
      ov(7 downto 0) := iv;
      tmp12_1415 <= ov(7 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1414_root_address_inst
    process(ptr_deref_1414_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1414_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_1414_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1430_addr_0
    process(ptr_deref_1430_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1430_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1430_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1430_base_resize
    process(iNsTr_5_1427) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_5_1427;
      ov := iv(6 downto 0);
      ptr_deref_1430_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1430_gather_scatter
    process(ptr_deref_1430_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1430_data_0;
      ov(31 downto 0) := iv;
      tmp15_1431 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1430_root_address_inst
    process(ptr_deref_1430_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1430_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1430_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1447_addr_0
    process(ptr_deref_1447_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1447_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_1447_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1447_base_resize
    process(iNsTr_6_1444) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_6_1444;
      ov := iv(0 downto 0);
      ptr_deref_1447_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1447_gather_scatter
    process(ptr_deref_1447_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1447_data_0;
      ov(7 downto 0) := iv;
      tmp23_1448 <= ov(7 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1447_root_address_inst
    process(ptr_deref_1447_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1447_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_1447_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1463_addr_0
    process(ptr_deref_1463_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1463_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1463_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1463_base_resize
    process(iNsTr_7_1460) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_7_1460;
      ov := iv(6 downto 0);
      ptr_deref_1463_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1463_gather_scatter
    process(ptr_deref_1463_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1463_data_0;
      ov(31 downto 0) := iv;
      tmp26_1464 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1463_root_address_inst
    process(ptr_deref_1463_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1463_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1463_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1475_addr_0
    process(ptr_deref_1475_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1475_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1475_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1475_base_resize
    process(iNsTr_8_1472) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_8_1472;
      ov := iv(6 downto 0);
      ptr_deref_1475_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1475_gather_scatter
    process(ptr_deref_1475_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1475_data_0;
      ov(31 downto 0) := iv;
      tmp35_1476 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1475_root_address_inst
    process(ptr_deref_1475_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1475_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1475_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1487_addr_0
    process(ptr_deref_1487_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1487_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1487_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1487_base_resize
    process(iNsTr_9_1484) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_9_1484;
      ov := iv(6 downto 0);
      ptr_deref_1487_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1487_gather_scatter
    process(ptr_deref_1487_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1487_data_0;
      ov(31 downto 0) := iv;
      tmp38_1488 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1487_root_address_inst
    process(ptr_deref_1487_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1487_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1487_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1505_addr_0
    process(ptr_deref_1505_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1505_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1505_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1505_base_resize
    process(iNsTr_10_1502) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_10_1502;
      ov := iv(6 downto 0);
      ptr_deref_1505_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1505_gather_scatter
    process(ptr_deref_1505_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1505_data_0;
      ov(31 downto 0) := iv;
      tmp75_1506 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1505_root_address_inst
    process(ptr_deref_1505_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1505_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1505_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1703_addr_0
    process(ptr_deref_1703_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1703_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1703_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1703_base_resize
    process(arrayidx_1700) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_1700;
      ov := iv(13 downto 0);
      ptr_deref_1703_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1703_gather_scatter
    process(ptr_deref_1703_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1703_data_0;
      ov(63 downto 0) := iv;
      tmp48_1704 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1703_root_address_inst
    process(ptr_deref_1703_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1703_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1703_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1733_addr_0
    process(ptr_deref_1733_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1733_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1733_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1733_base_resize
    process(arrayidx53_1731) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx53_1731;
      ov := iv(13 downto 0);
      ptr_deref_1733_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1733_gather_scatter
    process(tmp48_1704) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp48_1704;
      ov(63 downto 0) := iv;
      ptr_deref_1733_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1733_root_address_inst
    process(ptr_deref_1733_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1733_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1733_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1752_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_1751;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1752_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1752_branch_req_0,
          ack0 => if_stmt_1752_branch_ack_0,
          ack1 => if_stmt_1752_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1809_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp77_1808;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1809_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1809_branch_req_0,
          ack0 => if_stmt_1809_branch_ack_0,
          ack1 => if_stmt_1809_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1763_inst
    process(indvar_1645) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1645, type_cast_1762_wire_constant, tmp_var);
      indvarx_xnext_1764 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1771_inst
    process(input_dim1x_x1x_xph_1515) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_1515, type_cast_1770_wire_constant, tmp_var);
      inc_1772 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1790_inst
    process(inc72_1786, input_dim0x_x2x_xph_1522) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc72_1786, input_dim0x_x2x_xph_1522, tmp_var);
      inc72x_xinput_dim0x_x2_1791 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1549_inst
    process(mul_1545, conv3_1535) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul_1545, conv3_1535, tmp_var);
      add_1550 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1564_inst
    process(mul14_1560, tmp15_1431) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul14_1560, tmp15_1431, tmp_var);
      add16_1565 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1579_inst
    process(mul25_1575, tmp26_1464) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul25_1575, tmp26_1464, tmp_var);
      add27_1580 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1596_inst
    process(sub31_1591) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub31_1591, type_cast_1595_wire_constant, tmp_var);
      sext_1597 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1617_inst
    process(sub19_1612) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub19_1612, type_cast_1616_wire_constant, tmp_var);
      sext91_1618 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1636_inst
    process(conv37_1606, mul41_1632) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv37_1606, mul41_1632, tmp_var);
      add42_1637 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1666_inst
    process(mul7_1555, conv90_1662) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul7_1555, conv90_1662, tmp_var);
      add8_1667 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1671_inst
    process(mul43_1642, conv90_1662) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul43_1642, conv90_1662, tmp_var);
      add44_1672 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1745_inst
    process(conv56_1740) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv56_1740, type_cast_1744_wire_constant, tmp_var);
      add57_1746 <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1604_inst
    process(type_cast_1600_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1600_wire, type_cast_1603_wire_constant, tmp_var);
      ASHR_i32_i32_1604_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1625_inst
    process(type_cast_1621_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1621_wire, type_cast_1624_wire_constant, tmp_var);
      ASHR_i32_i32_1625_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1685_inst
    process(type_cast_1681_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1681_wire, type_cast_1684_wire_constant, tmp_var);
      ASHR_i32_i32_1685_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1717_inst
    process(type_cast_1713_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1713_wire, type_cast_1716_wire_constant, tmp_var);
      ASHR_i32_i32_1717_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1781_inst
    process(conv66_1777, div_1494) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv66_1777, div_1494, tmp_var);
      cmp68_1782 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1807_inst
    process(conv74_1803, div76_1512) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv74_1803, div76_1512, tmp_var);
      cmp77_1808 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1493_inst
    process(tmp4_1405) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_1405, type_cast_1492_wire_constant, tmp_var);
      div_1494 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1511_inst
    process(tmp75_1506) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp75_1506, type_cast_1510_wire_constant, tmp_var);
      div76_1512 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1657_inst
    process(indvar_1645) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_1645, type_cast_1656_wire_constant, tmp_var);
      input_dim2x_x1_1658 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1544_inst
    process(tmp4_1405, conv6_1540) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp4_1405, conv6_1540, tmp_var);
      mul_1545 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1554_inst
    process(add_1550, tmp1_1393) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add_1550, tmp1_1393, tmp_var);
      mul7_1555 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1559_inst
    process(conv13_1419, conv6_1540) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv13_1419, conv6_1540, tmp_var);
      mul14_1560 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1574_inst
    process(conv24_1452, conv3_1535) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv24_1452, conv3_1535, tmp_var);
      mul25_1575 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1631_inst
    process(tmp38_1488, conv40_1627) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp38_1488, conv40_1627, tmp_var);
      mul41_1632 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1641_inst
    process(add42_1637, tmp35_1476) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add42_1637, tmp35_1476, tmp_var);
      mul43_1642 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1590_inst
    process(sub30_1585) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(sub30_1585, type_cast_1589_wire_constant, tmp_var);
      sub31_1591 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1611_inst
    process(sub_1570) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(sub_1570, type_cast_1610_wire_constant, tmp_var);
      sub19_1612 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1677_inst
    process(add8_1667) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add8_1667, type_cast_1676_wire_constant, tmp_var);
      sext93_1678 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1709_inst
    process(add44_1672) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add44_1672, type_cast_1708_wire_constant, tmp_var);
      sext94_1710 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_1569_inst
    process(add16_1565, conv18_1438) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(add16_1565, conv18_1438, tmp_var);
      sub_1570 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_1584_inst
    process(add27_1580, conv18_1438) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(add27_1580, conv18_1438, tmp_var);
      sub30_1585 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_1750_inst
    process(add57_1746, tmp1_1393) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add57_1746, tmp1_1393, tmp_var);
      cmp_1751 <= tmp_var; --
    end process;
    -- shared split operator group (34) : array_obj_ref_1698_index_offset 
    ApIntAdd_group_34: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_1697_scaled;
      array_obj_ref_1698_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1698_index_offset_req_0;
      array_obj_ref_1698_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1698_index_offset_req_1;
      array_obj_ref_1698_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_34_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_34_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_34",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 34
    -- shared split operator group (35) : array_obj_ref_1729_index_offset 
    ApIntAdd_group_35: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom52_1728_scaled;
      array_obj_ref_1729_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1729_index_offset_req_0;
      array_obj_ref_1729_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1729_index_offset_req_1;
      array_obj_ref_1729_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_35_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_35_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_35",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 35
    -- unary operator type_cast_1533_inst
    process(input_dim1x_x1x_xph_1515) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim1x_x1x_xph_1515, tmp_var);
      type_cast_1533_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1538_inst
    process(input_dim0x_x2x_xph_1522) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim0x_x2x_xph_1522, tmp_var);
      type_cast_1538_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1691_inst
    process(shr_1687) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr_1687, tmp_var);
      type_cast_1691_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1722_inst
    process(shr51_1719) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr51_1719, tmp_var);
      type_cast_1722_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1738_inst
    process(input_dim2x_x1_1658) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim2x_x1_1658, tmp_var);
      type_cast_1738_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1775_inst
    process(inc_1772) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc_1772, tmp_var);
      type_cast_1775_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1801_inst
    process(inc72x_xinput_dim0x_x2_1791) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc72x_xinput_dim0x_x2_1791, tmp_var);
      type_cast_1801_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : LOAD_padding_1433_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_padding_1433_load_0_req_0;
      LOAD_padding_1433_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_padding_1433_load_0_req_1;
      LOAD_padding_1433_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_padding_1433_word_address_0;
      LOAD_padding_1433_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_7_lr_req(0),
          mack => memory_space_7_lr_ack(0),
          maddr => memory_space_7_lr_addr(0 downto 0),
          mtag => memory_space_7_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 8,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_7_lc_req(0),
          mack => memory_space_7_lc_ack(0),
          mdata => memory_space_7_lc_data(7 downto 0),
          mtag => memory_space_7_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_1392_load_0 ptr_deref_1404_load_0 ptr_deref_1505_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(20 downto 0);
      signal data_out: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_1392_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_1404_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1505_load_0_req_0;
      ptr_deref_1392_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_1404_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1505_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_1392_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_1404_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1505_load_0_req_1;
      ptr_deref_1392_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_1404_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1505_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      LoadGroup1_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1392_word_address_0 & ptr_deref_1404_word_address_0 & ptr_deref_1505_word_address_0;
      ptr_deref_1392_data_0 <= data_out(95 downto 64);
      ptr_deref_1404_data_0 <= data_out(63 downto 32);
      ptr_deref_1505_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 7,
        num_reqs => 3,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(6 downto 0),
          mtag => memory_space_1_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 32,
        num_reqs => 3,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(31 downto 0),
          mtag => memory_space_1_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : ptr_deref_1414_load_0 ptr_deref_1447_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1414_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1447_load_0_req_0;
      ptr_deref_1414_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1447_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1414_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1447_load_0_req_1;
      ptr_deref_1414_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1447_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup2_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup2_gI: SplitGuardInterface generic map(name => "LoadGroup2_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1414_word_address_0 & ptr_deref_1447_word_address_0;
      ptr_deref_1414_data_0 <= data_out(15 downto 8);
      ptr_deref_1447_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup2", addr_width => 1,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_8_lr_req(0),
          mack => memory_space_8_lr_ack(0),
          maddr => memory_space_8_lr_addr(0 downto 0),
          mtag => memory_space_8_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup2 load-complete ",
        data_width => 8,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_8_lc_req(0),
          mack => memory_space_8_lc_ack(0),
          mdata => memory_space_8_lc_data(7 downto 0),
          mtag => memory_space_8_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared load operator group (3) : ptr_deref_1430_load_0 ptr_deref_1463_load_0 
    LoadGroup3: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1430_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1463_load_0_req_0;
      ptr_deref_1430_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1463_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1430_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1463_load_0_req_1;
      ptr_deref_1430_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1463_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup3_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup3_gI: SplitGuardInterface generic map(name => "LoadGroup3_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1430_word_address_0 & ptr_deref_1463_word_address_0;
      ptr_deref_1430_data_0 <= data_out(63 downto 32);
      ptr_deref_1463_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup3", addr_width => 7,
        num_reqs => 2,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(6 downto 0),
          mtag => memory_space_2_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup3 load-complete ",
        data_width => 32,
        num_reqs => 2,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(31 downto 0),
          mtag => memory_space_2_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 3
    -- shared load operator group (4) : ptr_deref_1475_load_0 ptr_deref_1487_load_0 
    LoadGroup4: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1475_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1487_load_0_req_0;
      ptr_deref_1475_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1487_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1475_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1487_load_0_req_1;
      ptr_deref_1475_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1487_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup4_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup4_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup4_gI: SplitGuardInterface generic map(name => "LoadGroup4_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1475_word_address_0 & ptr_deref_1487_word_address_0;
      ptr_deref_1475_data_0 <= data_out(63 downto 32);
      ptr_deref_1487_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup4", addr_width => 7,
        num_reqs => 2,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(6 downto 0),
          mtag => memory_space_3_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup4 load-complete ",
        data_width => 32,
        num_reqs => 2,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(31 downto 0),
          mtag => memory_space_3_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 4
    -- shared load operator group (5) : ptr_deref_1703_load_0 
    LoadGroup5: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1703_load_0_req_0;
      ptr_deref_1703_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1703_load_0_req_1;
      ptr_deref_1703_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup5_gI: SplitGuardInterface generic map(name => "LoadGroup5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1703_word_address_0;
      ptr_deref_1703_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup5", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_4_lr_req(0),
          mack => memory_space_4_lr_ack(0),
          maddr => memory_space_4_lr_addr(13 downto 0),
          mtag => memory_space_4_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup5 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_4_lc_req(0),
          mack => memory_space_4_lc_ack(0),
          mdata => memory_space_4_lc_data(63 downto 0),
          mtag => memory_space_4_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 5
    -- shared store operator group (0) : ptr_deref_1733_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1733_store_0_req_0;
      ptr_deref_1733_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1733_store_0_req_1;
      ptr_deref_1733_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1733_word_address_0;
      data_in <= ptr_deref_1733_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_6_sr_req(0),
          mack => memory_space_6_sr_ack(0),
          maddr => memory_space_6_sr_addr(13 downto 0),
          mdata => memory_space_6_sr_data(63 downto 0),
          mtag => memory_space_6_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_6_sc_req(0),
          mack => memory_space_6_sc_ack(0),
          mtag => memory_space_6_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block0_start_1379_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block0_start_1379_inst_req_0;
      RPIPE_Block0_start_1379_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block0_start_1379_inst_req_1;
      RPIPE_Block0_start_1379_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call_1380 <= data_out(15 downto 0);
      Block0_start_read_0_gI: SplitGuardInterface generic map(name => "Block0_start_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block0_start_read_0: InputPortRevised -- 
        generic map ( name => "Block0_start_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block0_start_pipe_read_req(0),
          oack => Block0_start_pipe_read_ack(0),
          odata => Block0_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block0_done_1817_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block0_done_1817_inst_req_0;
      WPIPE_Block0_done_1817_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block0_done_1817_inst_req_1;
      WPIPE_Block0_done_1817_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= call_1380;
      Block0_done_write_0_gI: SplitGuardInterface generic map(name => "Block0_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block0_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block0_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block0_done_pipe_write_req(0),
          oack => Block0_done_pipe_write_ack(0),
          odata => Block0_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeA_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeB is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_7_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_8_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_8_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_8_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_8_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_8_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_8_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_4_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_4_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_6_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_6_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_sc_tag :  in  std_logic_vector(0 downto 0);
    Block1_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block1_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block1_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block1_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block1_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block1_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeB;
architecture convTransposeB_arch of convTransposeB is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeB_CP_5119_start: Boolean;
  signal convTransposeB_CP_5119_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal ptr_deref_1888_load_0_ack_1 : boolean;
  signal type_cast_1895_inst_req_1 : boolean;
  signal type_cast_1895_inst_ack_1 : boolean;
  signal LOAD_padding_1891_load_0_ack_0 : boolean;
  signal ptr_deref_1888_load_0_req_1 : boolean;
  signal LOAD_padding_1891_load_0_req_0 : boolean;
  signal type_cast_1909_inst_ack_1 : boolean;
  signal ptr_deref_1933_load_0_req_0 : boolean;
  signal ptr_deref_1933_load_0_ack_0 : boolean;
  signal type_cast_1895_inst_req_0 : boolean;
  signal ptr_deref_1921_load_0_req_1 : boolean;
  signal ptr_deref_1921_load_0_ack_1 : boolean;
  signal LOAD_padding_1891_load_0_req_1 : boolean;
  signal ptr_deref_1921_load_0_req_0 : boolean;
  signal ptr_deref_1921_load_0_ack_0 : boolean;
  signal type_cast_1895_inst_ack_0 : boolean;
  signal LOAD_padding_1891_load_0_ack_1 : boolean;
  signal ptr_deref_1905_load_0_req_0 : boolean;
  signal type_cast_1909_inst_req_0 : boolean;
  signal type_cast_1909_inst_ack_0 : boolean;
  signal ptr_deref_1905_load_0_ack_0 : boolean;
  signal ptr_deref_1905_load_0_req_1 : boolean;
  signal ptr_deref_1905_load_0_ack_1 : boolean;
  signal type_cast_1909_inst_req_1 : boolean;
  signal ptr_deref_1933_load_0_req_1 : boolean;
  signal ptr_deref_1933_load_0_ack_1 : boolean;
  signal RPIPE_Block1_start_1827_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1827_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1827_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1827_inst_ack_1 : boolean;
  signal ptr_deref_1840_load_0_req_0 : boolean;
  signal ptr_deref_1840_load_0_ack_0 : boolean;
  signal ptr_deref_1840_load_0_req_1 : boolean;
  signal ptr_deref_1840_load_0_ack_1 : boolean;
  signal type_cast_1850_inst_req_0 : boolean;
  signal type_cast_1850_inst_ack_0 : boolean;
  signal type_cast_1850_inst_req_1 : boolean;
  signal type_cast_1850_inst_ack_1 : boolean;
  signal ptr_deref_1862_load_0_req_0 : boolean;
  signal ptr_deref_1862_load_0_ack_0 : boolean;
  signal ptr_deref_1862_load_0_req_1 : boolean;
  signal ptr_deref_1862_load_0_ack_1 : boolean;
  signal ptr_deref_1872_load_0_req_0 : boolean;
  signal ptr_deref_1872_load_0_ack_0 : boolean;
  signal ptr_deref_1872_load_0_req_1 : boolean;
  signal ptr_deref_1872_load_0_ack_1 : boolean;
  signal type_cast_1876_inst_req_0 : boolean;
  signal type_cast_1876_inst_ack_0 : boolean;
  signal type_cast_1876_inst_req_1 : boolean;
  signal type_cast_1876_inst_ack_1 : boolean;
  signal ptr_deref_1888_load_0_req_0 : boolean;
  signal ptr_deref_1888_load_0_ack_0 : boolean;
  signal ptr_deref_1945_load_0_req_0 : boolean;
  signal ptr_deref_1945_load_0_ack_0 : boolean;
  signal ptr_deref_1945_load_0_req_1 : boolean;
  signal ptr_deref_1945_load_0_ack_1 : boolean;
  signal ptr_deref_1957_load_0_req_0 : boolean;
  signal ptr_deref_1957_load_0_ack_0 : boolean;
  signal ptr_deref_1957_load_0_req_1 : boolean;
  signal ptr_deref_1957_load_0_ack_1 : boolean;
  signal type_cast_1984_inst_req_0 : boolean;
  signal type_cast_1984_inst_ack_0 : boolean;
  signal type_cast_1984_inst_req_1 : boolean;
  signal type_cast_1984_inst_ack_1 : boolean;
  signal type_cast_1989_inst_req_0 : boolean;
  signal type_cast_1989_inst_ack_0 : boolean;
  signal type_cast_1989_inst_req_1 : boolean;
  signal type_cast_1989_inst_ack_1 : boolean;
  signal type_cast_2111_inst_req_0 : boolean;
  signal type_cast_2111_inst_ack_0 : boolean;
  signal type_cast_2111_inst_req_1 : boolean;
  signal type_cast_2111_inst_ack_1 : boolean;
  signal type_cast_2141_inst_req_0 : boolean;
  signal type_cast_2141_inst_ack_0 : boolean;
  signal type_cast_2141_inst_req_1 : boolean;
  signal type_cast_2141_inst_ack_1 : boolean;
  signal array_obj_ref_2147_index_offset_req_0 : boolean;
  signal array_obj_ref_2147_index_offset_ack_0 : boolean;
  signal array_obj_ref_2147_index_offset_req_1 : boolean;
  signal array_obj_ref_2147_index_offset_ack_1 : boolean;
  signal addr_of_2148_final_reg_req_0 : boolean;
  signal addr_of_2148_final_reg_ack_0 : boolean;
  signal addr_of_2148_final_reg_req_1 : boolean;
  signal addr_of_2148_final_reg_ack_1 : boolean;
  signal ptr_deref_2152_load_0_req_0 : boolean;
  signal ptr_deref_2152_load_0_ack_0 : boolean;
  signal ptr_deref_2152_load_0_req_1 : boolean;
  signal ptr_deref_2152_load_0_ack_1 : boolean;
  signal type_cast_2172_inst_req_0 : boolean;
  signal type_cast_2172_inst_ack_0 : boolean;
  signal type_cast_2172_inst_req_1 : boolean;
  signal type_cast_2172_inst_ack_1 : boolean;
  signal array_obj_ref_2178_index_offset_req_0 : boolean;
  signal array_obj_ref_2178_index_offset_ack_0 : boolean;
  signal array_obj_ref_2178_index_offset_req_1 : boolean;
  signal array_obj_ref_2178_index_offset_ack_1 : boolean;
  signal addr_of_2179_final_reg_req_0 : boolean;
  signal addr_of_2179_final_reg_ack_0 : boolean;
  signal addr_of_2179_final_reg_req_1 : boolean;
  signal addr_of_2179_final_reg_ack_1 : boolean;
  signal ptr_deref_2182_store_0_req_0 : boolean;
  signal ptr_deref_2182_store_0_ack_0 : boolean;
  signal ptr_deref_2182_store_0_req_1 : boolean;
  signal ptr_deref_2182_store_0_ack_1 : boolean;
  signal type_cast_2188_inst_req_0 : boolean;
  signal type_cast_2188_inst_ack_0 : boolean;
  signal type_cast_2188_inst_req_1 : boolean;
  signal type_cast_2188_inst_ack_1 : boolean;
  signal if_stmt_2201_branch_req_0 : boolean;
  signal if_stmt_2201_branch_ack_1 : boolean;
  signal if_stmt_2201_branch_ack_0 : boolean;
  signal type_cast_2225_inst_req_0 : boolean;
  signal type_cast_2225_inst_ack_0 : boolean;
  signal type_cast_2225_inst_req_1 : boolean;
  signal type_cast_2225_inst_ack_1 : boolean;
  signal if_stmt_2232_branch_req_0 : boolean;
  signal if_stmt_2232_branch_ack_1 : boolean;
  signal if_stmt_2232_branch_ack_0 : boolean;
  signal type_cast_2253_inst_req_0 : boolean;
  signal type_cast_2253_inst_ack_0 : boolean;
  signal type_cast_2253_inst_req_1 : boolean;
  signal type_cast_2253_inst_ack_1 : boolean;
  signal type_cast_2273_inst_req_0 : boolean;
  signal type_cast_2273_inst_ack_0 : boolean;
  signal type_cast_2273_inst_req_1 : boolean;
  signal type_cast_2273_inst_ack_1 : boolean;
  signal if_stmt_2280_branch_req_0 : boolean;
  signal if_stmt_2280_branch_ack_1 : boolean;
  signal if_stmt_2280_branch_ack_0 : boolean;
  signal WPIPE_Block1_done_2288_inst_req_0 : boolean;
  signal WPIPE_Block1_done_2288_inst_ack_0 : boolean;
  signal WPIPE_Block1_done_2288_inst_req_1 : boolean;
  signal WPIPE_Block1_done_2288_inst_ack_1 : boolean;
  signal phi_stmt_1973_req_0 : boolean;
  signal type_cast_1970_inst_req_0 : boolean;
  signal type_cast_1970_inst_ack_0 : boolean;
  signal type_cast_1970_inst_req_1 : boolean;
  signal type_cast_1970_inst_ack_1 : boolean;
  signal phi_stmt_1967_req_0 : boolean;
  signal type_cast_1979_inst_req_0 : boolean;
  signal type_cast_1979_inst_ack_0 : boolean;
  signal type_cast_1979_inst_req_1 : boolean;
  signal type_cast_1979_inst_ack_1 : boolean;
  signal phi_stmt_1973_req_1 : boolean;
  signal type_cast_1972_inst_req_0 : boolean;
  signal type_cast_1972_inst_ack_0 : boolean;
  signal type_cast_1972_inst_req_1 : boolean;
  signal type_cast_1972_inst_ack_1 : boolean;
  signal phi_stmt_1967_req_1 : boolean;
  signal phi_stmt_1967_ack_0 : boolean;
  signal phi_stmt_1973_ack_0 : boolean;
  signal type_cast_2101_inst_req_0 : boolean;
  signal type_cast_2101_inst_ack_0 : boolean;
  signal type_cast_2101_inst_req_1 : boolean;
  signal type_cast_2101_inst_ack_1 : boolean;
  signal phi_stmt_2095_req_1 : boolean;
  signal phi_stmt_2095_req_0 : boolean;
  signal phi_stmt_2095_ack_0 : boolean;
  signal type_cast_2262_inst_req_0 : boolean;
  signal type_cast_2262_inst_ack_0 : boolean;
  signal type_cast_2262_inst_req_1 : boolean;
  signal type_cast_2262_inst_ack_1 : boolean;
  signal phi_stmt_2257_req_1 : boolean;
  signal type_cast_2268_inst_req_0 : boolean;
  signal type_cast_2268_inst_ack_0 : boolean;
  signal type_cast_2268_inst_req_1 : boolean;
  signal type_cast_2268_inst_ack_1 : boolean;
  signal phi_stmt_2263_req_1 : boolean;
  signal type_cast_2260_inst_req_0 : boolean;
  signal type_cast_2260_inst_ack_0 : boolean;
  signal type_cast_2260_inst_req_1 : boolean;
  signal type_cast_2260_inst_ack_1 : boolean;
  signal phi_stmt_2257_req_0 : boolean;
  signal type_cast_2266_inst_req_0 : boolean;
  signal type_cast_2266_inst_ack_0 : boolean;
  signal type_cast_2266_inst_req_1 : boolean;
  signal type_cast_2266_inst_ack_1 : boolean;
  signal phi_stmt_2263_req_0 : boolean;
  signal phi_stmt_2257_ack_0 : boolean;
  signal phi_stmt_2263_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeB_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeB_CP_5119_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeB_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeB_CP_5119_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeB_CP_5119_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeB_CP_5119_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeB_CP_5119: Block -- control-path 
    signal convTransposeB_CP_5119_elements: BooleanArray(112 downto 0);
    -- 
  begin -- 
    convTransposeB_CP_5119_elements(0) <= convTransposeB_CP_5119_start;
    convTransposeB_CP_5119_symbol <= convTransposeB_CP_5119_elements(72);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1825/$entry
      -- CP-element group 0: 	 branch_block_stmt_1825/branch_block_stmt_1825__entry__
      -- CP-element group 0: 	 branch_block_stmt_1825/assign_stmt_1828__entry__
      -- CP-element group 0: 	 branch_block_stmt_1825/assign_stmt_1828/$entry
      -- CP-element group 0: 	 branch_block_stmt_1825/assign_stmt_1828/RPIPE_Block1_start_1827_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1825/assign_stmt_1828/RPIPE_Block1_start_1827_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1825/assign_stmt_1828/RPIPE_Block1_start_1827_Sample/rr
      -- 
    rr_5177_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5177_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(0), ack => RPIPE_Block1_start_1827_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_1825/assign_stmt_1828/RPIPE_Block1_start_1827_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_1825/assign_stmt_1828/RPIPE_Block1_start_1827_update_start_
      -- CP-element group 1: 	 branch_block_stmt_1825/assign_stmt_1828/RPIPE_Block1_start_1827_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_1825/assign_stmt_1828/RPIPE_Block1_start_1827_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_1825/assign_stmt_1828/RPIPE_Block1_start_1827_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1825/assign_stmt_1828/RPIPE_Block1_start_1827_Update/cr
      -- 
    ra_5178_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1827_inst_ack_0, ack => convTransposeB_CP_5119_elements(1)); -- 
    cr_5182_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5182_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(1), ack => RPIPE_Block1_start_1827_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  place  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	20 
    -- CP-element group 2: 	22 
    -- CP-element group 2: 	26 
    -- CP-element group 2: 	15 
    -- CP-element group 2: 	16 
    -- CP-element group 2: 	18 
    -- CP-element group 2: 	19 
    -- CP-element group 2: 	13 
    -- CP-element group 2: 	12 
    -- CP-element group 2: 	27 
    -- CP-element group 2: 	30 
    -- CP-element group 2: 	14 
    -- CP-element group 2: 	28 
    -- CP-element group 2: 	29 
    -- CP-element group 2: 	23 
    -- CP-element group 2: 	24 
    -- CP-element group 2: 	25 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	4 
    -- CP-element group 2: 	6 
    -- CP-element group 2: 	7 
    -- CP-element group 2: 	8 
    -- CP-element group 2: 	9 
    -- CP-element group 2: 	10 
    -- CP-element group 2:  members (265) 
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1905_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1888_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/type_cast_1895_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/LOAD_padding_1891_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1905_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1905_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/LOAD_padding_1891_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1905_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1905_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1905_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1888_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1905_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1905_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/LOAD_padding_1891_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1905_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1921_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1921_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/type_cast_1909_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1905_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/LOAD_padding_1891_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1921_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1921_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1933_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1933_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1888_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1933_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1933_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1921_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/LOAD_padding_1891_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1921_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1921_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1905_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1933_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1933_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1933_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1921_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1921_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/LOAD_padding_1891_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1905_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1905_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1921_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1888_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/LOAD_padding_1891_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1905_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1921_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1933_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1921_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/LOAD_padding_1891_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/LOAD_padding_1891_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1933_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1933_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1921_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/LOAD_padding_1891_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1933_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1933_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1921_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1921_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1905_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1933_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1905_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1905_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1933_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1933_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1921_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1921_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1933_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1945_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1921_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/LOAD_padding_1891_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1921_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1921_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1933_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1933_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1933_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1905_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1905_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1933_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1933_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1905_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1921_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1933_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1933_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1905_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1905_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1921_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/type_cast_1909_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/type_cast_1895_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1921_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1905_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1905_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/LOAD_padding_1891_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1921_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1921_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1921_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/type_cast_1909_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/type_cast_1895_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1905_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1933_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1933_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1933_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1828__exit__
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964__entry__
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1828/$exit
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1828/RPIPE_Block1_start_1827_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1828/RPIPE_Block1_start_1827_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1828/RPIPE_Block1_start_1827_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1840_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1840_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1840_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1840_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1840_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1840_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1840_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1840_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1840_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1840_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1840_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1840_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1840_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1840_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1840_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1840_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1840_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1840_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1840_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1840_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1840_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1840_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1840_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1840_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1840_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1840_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/type_cast_1850_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/type_cast_1850_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/type_cast_1850_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1862_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1862_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1862_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1862_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1862_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1862_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1862_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1862_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1862_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1862_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1862_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1862_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1862_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1862_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1862_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1862_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1862_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1862_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1862_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1862_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1862_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1862_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1862_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1862_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1862_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1862_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1872_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1905_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1872_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1872_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1872_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1872_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1872_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1872_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1872_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1872_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1872_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1872_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1872_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1872_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1872_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1872_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1872_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1872_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1872_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1872_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1872_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1872_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1872_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1872_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1872_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1872_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1872_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/type_cast_1876_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/type_cast_1876_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/type_cast_1876_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1888_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1888_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1888_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1888_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1888_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1888_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1888_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1888_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1888_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1888_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1888_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1888_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1888_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1888_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1888_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1888_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1888_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1888_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1888_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1888_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1888_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1888_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1945_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1945_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1945_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1945_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1945_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1945_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1945_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1945_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1945_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1945_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1945_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1945_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1945_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1945_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1945_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1945_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1945_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1945_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1945_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1945_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1945_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1945_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1945_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1945_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1945_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1957_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1957_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1957_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1957_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1957_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1957_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1957_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1957_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1957_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1957_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1957_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1957_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1957_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1957_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1957_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1957_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1957_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1957_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1957_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1957_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1957_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1957_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1957_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1957_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1957_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1957_Update/word_access_complete/word_0/cr
      -- 
    ca_5183_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1827_inst_ack_1, ack => convTransposeB_CP_5119_elements(2)); -- 
    cr_5460_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5460_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(2), ack => type_cast_1895_inst_req_1); -- 
    cr_5408_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5408_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(2), ack => ptr_deref_1888_load_0_req_1); -- 
    rr_5430_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5430_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(2), ack => LOAD_padding_1891_load_0_req_0); -- 
    rr_5608_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5608_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(2), ack => ptr_deref_1933_load_0_req_0); -- 
    cr_5569_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5569_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(2), ack => ptr_deref_1921_load_0_req_1); -- 
    cr_5441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(2), ack => LOAD_padding_1891_load_0_req_1); -- 
    rr_5558_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5558_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(2), ack => ptr_deref_1921_load_0_req_0); -- 
    rr_5494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(2), ack => ptr_deref_1905_load_0_req_0); -- 
    cr_5505_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5505_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(2), ack => ptr_deref_1905_load_0_req_1); -- 
    cr_5524_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5524_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(2), ack => type_cast_1909_inst_req_1); -- 
    cr_5619_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5619_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(2), ack => ptr_deref_1933_load_0_req_1); -- 
    rr_5219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(2), ack => ptr_deref_1840_load_0_req_0); -- 
    cr_5230_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5230_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(2), ack => ptr_deref_1840_load_0_req_1); -- 
    cr_5249_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5249_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(2), ack => type_cast_1850_inst_req_1); -- 
    rr_5283_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5283_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(2), ack => ptr_deref_1862_load_0_req_0); -- 
    cr_5294_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5294_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(2), ack => ptr_deref_1862_load_0_req_1); -- 
    rr_5333_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5333_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(2), ack => ptr_deref_1872_load_0_req_0); -- 
    cr_5344_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5344_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(2), ack => ptr_deref_1872_load_0_req_1); -- 
    cr_5363_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5363_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(2), ack => type_cast_1876_inst_req_1); -- 
    rr_5397_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5397_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(2), ack => ptr_deref_1888_load_0_req_0); -- 
    rr_5658_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5658_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(2), ack => ptr_deref_1945_load_0_req_0); -- 
    cr_5669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(2), ack => ptr_deref_1945_load_0_req_1); -- 
    rr_5708_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5708_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(2), ack => ptr_deref_1957_load_0_req_0); -- 
    cr_5719_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5719_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(2), ack => ptr_deref_1957_load_0_req_1); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (5) 
      -- CP-element group 3: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1840_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1840_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1840_Sample/word_access_start/$exit
      -- CP-element group 3: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1840_Sample/word_access_start/word_0/$exit
      -- CP-element group 3: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1840_Sample/word_access_start/word_0/ra
      -- 
    ra_5220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1840_load_0_ack_0, ack => convTransposeB_CP_5119_elements(3)); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	2 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (12) 
      -- CP-element group 4: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1840_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1840_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1840_Update/word_access_complete/$exit
      -- CP-element group 4: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1840_Update/word_access_complete/word_0/$exit
      -- CP-element group 4: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1840_Update/word_access_complete/word_0/ca
      -- CP-element group 4: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1840_Update/ptr_deref_1840_Merge/$entry
      -- CP-element group 4: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1840_Update/ptr_deref_1840_Merge/$exit
      -- CP-element group 4: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1840_Update/ptr_deref_1840_Merge/merge_req
      -- CP-element group 4: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1840_Update/ptr_deref_1840_Merge/merge_ack
      -- CP-element group 4: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/type_cast_1850_sample_start_
      -- CP-element group 4: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/type_cast_1850_Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/type_cast_1850_Sample/rr
      -- 
    ca_5231_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1840_load_0_ack_1, ack => convTransposeB_CP_5119_elements(4)); -- 
    rr_5244_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5244_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(4), ack => type_cast_1850_inst_req_0); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/type_cast_1850_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/type_cast_1850_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/type_cast_1850_Sample/ra
      -- 
    ra_5245_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1850_inst_ack_0, ack => convTransposeB_CP_5119_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	2 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	31 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/type_cast_1850_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/type_cast_1850_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/type_cast_1850_Update/ca
      -- 
    ca_5250_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1850_inst_ack_1, ack => convTransposeB_CP_5119_elements(6)); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	2 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (5) 
      -- CP-element group 7: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1862_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1862_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1862_Sample/word_access_start/$exit
      -- CP-element group 7: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1862_Sample/word_access_start/word_0/$exit
      -- CP-element group 7: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1862_Sample/word_access_start/word_0/ra
      -- 
    ra_5284_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1862_load_0_ack_0, ack => convTransposeB_CP_5119_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	31 
    -- CP-element group 8:  members (9) 
      -- CP-element group 8: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1862_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1862_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1862_Update/word_access_complete/$exit
      -- CP-element group 8: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1862_Update/word_access_complete/word_0/$exit
      -- CP-element group 8: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1862_Update/word_access_complete/word_0/ca
      -- CP-element group 8: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1862_Update/ptr_deref_1862_Merge/$entry
      -- CP-element group 8: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1862_Update/ptr_deref_1862_Merge/$exit
      -- CP-element group 8: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1862_Update/ptr_deref_1862_Merge/merge_req
      -- CP-element group 8: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1862_Update/ptr_deref_1862_Merge/merge_ack
      -- 
    ca_5295_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1862_load_0_ack_1, ack => convTransposeB_CP_5119_elements(8)); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	2 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (5) 
      -- CP-element group 9: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1872_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1872_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1872_Sample/word_access_start/$exit
      -- CP-element group 9: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1872_Sample/word_access_start/word_0/$exit
      -- CP-element group 9: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1872_Sample/word_access_start/word_0/ra
      -- 
    ra_5334_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1872_load_0_ack_0, ack => convTransposeB_CP_5119_elements(9)); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	2 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (12) 
      -- CP-element group 10: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1872_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1872_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1872_Update/word_access_complete/$exit
      -- CP-element group 10: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1872_Update/word_access_complete/word_0/$exit
      -- CP-element group 10: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1872_Update/word_access_complete/word_0/ca
      -- CP-element group 10: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1872_Update/ptr_deref_1872_Merge/$entry
      -- CP-element group 10: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1872_Update/ptr_deref_1872_Merge/$exit
      -- CP-element group 10: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1872_Update/ptr_deref_1872_Merge/merge_req
      -- CP-element group 10: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1872_Update/ptr_deref_1872_Merge/merge_ack
      -- CP-element group 10: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/type_cast_1876_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/type_cast_1876_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/type_cast_1876_Sample/rr
      -- 
    ca_5345_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1872_load_0_ack_1, ack => convTransposeB_CP_5119_elements(10)); -- 
    rr_5358_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5358_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(10), ack => type_cast_1876_inst_req_0); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/type_cast_1876_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/type_cast_1876_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/type_cast_1876_Sample/ra
      -- 
    ra_5359_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1876_inst_ack_0, ack => convTransposeB_CP_5119_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	2 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	31 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/type_cast_1876_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/type_cast_1876_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/type_cast_1876_Update/ca
      -- 
    ca_5364_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1876_inst_ack_1, ack => convTransposeB_CP_5119_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	2 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (5) 
      -- CP-element group 13: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1888_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1888_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1888_Sample/word_access_start/$exit
      -- CP-element group 13: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1888_Sample/word_access_start/word_0/$exit
      -- CP-element group 13: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1888_Sample/word_access_start/word_0/ra
      -- 
    ra_5398_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1888_load_0_ack_0, ack => convTransposeB_CP_5119_elements(13)); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	2 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	31 
    -- CP-element group 14:  members (9) 
      -- CP-element group 14: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1888_Update/word_access_complete/word_0/ca
      -- CP-element group 14: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1888_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1888_Update/ptr_deref_1888_Merge/$exit
      -- CP-element group 14: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1888_Update/ptr_deref_1888_Merge/$entry
      -- CP-element group 14: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1888_Update/ptr_deref_1888_Merge/merge_ack
      -- CP-element group 14: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1888_Update/word_access_complete/word_0/$exit
      -- CP-element group 14: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1888_Update/ptr_deref_1888_Merge/merge_req
      -- CP-element group 14: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1888_Update/word_access_complete/$exit
      -- CP-element group 14: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1888_update_completed_
      -- 
    ca_5409_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1888_load_0_ack_1, ack => convTransposeB_CP_5119_elements(14)); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	2 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (5) 
      -- CP-element group 15: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/LOAD_padding_1891_Sample/word_access_start/word_0/ra
      -- CP-element group 15: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/LOAD_padding_1891_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/LOAD_padding_1891_Sample/word_access_start/$exit
      -- CP-element group 15: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/LOAD_padding_1891_Sample/word_access_start/word_0/$exit
      -- CP-element group 15: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/LOAD_padding_1891_Sample/$exit
      -- 
    ra_5431_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_padding_1891_load_0_ack_0, ack => convTransposeB_CP_5119_elements(15)); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	2 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (12) 
      -- CP-element group 16: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/LOAD_padding_1891_Update/word_access_complete/$exit
      -- CP-element group 16: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/LOAD_padding_1891_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/type_cast_1895_Sample/$entry
      -- CP-element group 16: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/LOAD_padding_1891_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/type_cast_1895_Sample/rr
      -- CP-element group 16: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/LOAD_padding_1891_Update/word_access_complete/word_0/$exit
      -- CP-element group 16: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/LOAD_padding_1891_Update/word_access_complete/word_0/ca
      -- CP-element group 16: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/LOAD_padding_1891_Update/LOAD_padding_1891_Merge/$entry
      -- CP-element group 16: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/LOAD_padding_1891_Update/LOAD_padding_1891_Merge/$exit
      -- CP-element group 16: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/LOAD_padding_1891_Update/LOAD_padding_1891_Merge/merge_req
      -- CP-element group 16: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/LOAD_padding_1891_Update/LOAD_padding_1891_Merge/merge_ack
      -- CP-element group 16: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/type_cast_1895_sample_start_
      -- 
    ca_5442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_padding_1891_load_0_ack_1, ack => convTransposeB_CP_5119_elements(16)); -- 
    rr_5455_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5455_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(16), ack => type_cast_1895_inst_req_0); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/type_cast_1895_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/type_cast_1895_Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/type_cast_1895_sample_completed_
      -- 
    ra_5456_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1895_inst_ack_0, ack => convTransposeB_CP_5119_elements(17)); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	2 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	31 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/type_cast_1895_Update/ca
      -- CP-element group 18: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/type_cast_1895_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/type_cast_1895_update_completed_
      -- 
    ca_5461_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1895_inst_ack_1, ack => convTransposeB_CP_5119_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	2 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (5) 
      -- CP-element group 19: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1905_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1905_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1905_Sample/word_access_start/word_0/$exit
      -- CP-element group 19: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1905_Sample/word_access_start/word_0/ra
      -- CP-element group 19: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1905_Sample/word_access_start/$exit
      -- 
    ra_5495_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1905_load_0_ack_0, ack => convTransposeB_CP_5119_elements(19)); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	2 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (12) 
      -- CP-element group 20: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1905_Update/word_access_complete/$exit
      -- CP-element group 20: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/type_cast_1909_Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/type_cast_1909_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1905_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/type_cast_1909_Sample/rr
      -- CP-element group 20: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1905_Update/word_access_complete/word_0/$exit
      -- CP-element group 20: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1905_Update/word_access_complete/word_0/ca
      -- CP-element group 20: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1905_Update/ptr_deref_1905_Merge/$entry
      -- CP-element group 20: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1905_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1905_Update/ptr_deref_1905_Merge/$exit
      -- CP-element group 20: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1905_Update/ptr_deref_1905_Merge/merge_req
      -- CP-element group 20: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1905_Update/ptr_deref_1905_Merge/merge_ack
      -- 
    ca_5506_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1905_load_0_ack_1, ack => convTransposeB_CP_5119_elements(20)); -- 
    rr_5519_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5519_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(20), ack => type_cast_1909_inst_req_0); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/type_cast_1909_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/type_cast_1909_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/type_cast_1909_Sample/ra
      -- 
    ra_5520_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1909_inst_ack_0, ack => convTransposeB_CP_5119_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	2 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	31 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/type_cast_1909_Update/ca
      -- CP-element group 22: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/type_cast_1909_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/type_cast_1909_update_completed_
      -- 
    ca_5525_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1909_inst_ack_1, ack => convTransposeB_CP_5119_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	2 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (5) 
      -- CP-element group 23: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1921_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1921_Sample/word_access_start/word_0/$exit
      -- CP-element group 23: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1921_Sample/word_access_start/word_0/ra
      -- CP-element group 23: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1921_Sample/word_access_start/$exit
      -- CP-element group 23: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1921_Sample/$exit
      -- 
    ra_5559_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1921_load_0_ack_0, ack => convTransposeB_CP_5119_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	2 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	31 
    -- CP-element group 24:  members (9) 
      -- CP-element group 24: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1921_Update/word_access_complete/word_0/ca
      -- CP-element group 24: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1921_Update/ptr_deref_1921_Merge/$entry
      -- CP-element group 24: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1921_Update/ptr_deref_1921_Merge/$exit
      -- CP-element group 24: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1921_Update/ptr_deref_1921_Merge/merge_req
      -- CP-element group 24: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1921_Update/ptr_deref_1921_Merge/merge_ack
      -- CP-element group 24: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1921_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1921_Update/word_access_complete/$exit
      -- CP-element group 24: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1921_Update/word_access_complete/word_0/$exit
      -- CP-element group 24: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1921_update_completed_
      -- 
    ca_5570_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1921_load_0_ack_1, ack => convTransposeB_CP_5119_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	2 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (5) 
      -- CP-element group 25: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1933_Sample/word_access_start/$exit
      -- CP-element group 25: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1933_Sample/word_access_start/word_0/ra
      -- CP-element group 25: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1933_Sample/word_access_start/word_0/$exit
      -- CP-element group 25: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1933_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1933_sample_completed_
      -- 
    ra_5609_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1933_load_0_ack_0, ack => convTransposeB_CP_5119_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	2 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	31 
    -- CP-element group 26:  members (9) 
      -- CP-element group 26: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1933_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1933_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1933_Update/ptr_deref_1933_Merge/merge_req
      -- CP-element group 26: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1933_Update/ptr_deref_1933_Merge/merge_ack
      -- CP-element group 26: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1933_Update/word_access_complete/word_0/ca
      -- CP-element group 26: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1933_Update/ptr_deref_1933_Merge/$entry
      -- CP-element group 26: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1933_Update/ptr_deref_1933_Merge/$exit
      -- CP-element group 26: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1933_Update/word_access_complete/$exit
      -- CP-element group 26: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1933_Update/word_access_complete/word_0/$exit
      -- 
    ca_5620_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1933_load_0_ack_1, ack => convTransposeB_CP_5119_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	2 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (5) 
      -- CP-element group 27: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1945_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1945_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1945_Sample/word_access_start/$exit
      -- CP-element group 27: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1945_Sample/word_access_start/word_0/$exit
      -- CP-element group 27: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1945_Sample/word_access_start/word_0/ra
      -- 
    ra_5659_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1945_load_0_ack_0, ack => convTransposeB_CP_5119_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	2 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	31 
    -- CP-element group 28:  members (9) 
      -- CP-element group 28: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1945_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1945_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1945_Update/word_access_complete/$exit
      -- CP-element group 28: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1945_Update/word_access_complete/word_0/$exit
      -- CP-element group 28: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1945_Update/word_access_complete/word_0/ca
      -- CP-element group 28: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1945_Update/ptr_deref_1945_Merge/$entry
      -- CP-element group 28: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1945_Update/ptr_deref_1945_Merge/$exit
      -- CP-element group 28: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1945_Update/ptr_deref_1945_Merge/merge_req
      -- CP-element group 28: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1945_Update/ptr_deref_1945_Merge/merge_ack
      -- 
    ca_5670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1945_load_0_ack_1, ack => convTransposeB_CP_5119_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	2 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (5) 
      -- CP-element group 29: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1957_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1957_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1957_Sample/word_access_start/$exit
      -- CP-element group 29: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1957_Sample/word_access_start/word_0/$exit
      -- CP-element group 29: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1957_Sample/word_access_start/word_0/ra
      -- 
    ra_5709_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1957_load_0_ack_0, ack => convTransposeB_CP_5119_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	2 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (9) 
      -- CP-element group 30: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1957_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1957_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1957_Update/word_access_complete/$exit
      -- CP-element group 30: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1957_Update/word_access_complete/word_0/$exit
      -- CP-element group 30: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1957_Update/word_access_complete/word_0/ca
      -- CP-element group 30: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1957_Update/ptr_deref_1957_Merge/$entry
      -- CP-element group 30: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1957_Update/ptr_deref_1957_Merge/$exit
      -- CP-element group 30: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1957_Update/ptr_deref_1957_Merge/merge_req
      -- CP-element group 30: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/ptr_deref_1957_Update/ptr_deref_1957_Merge/merge_ack
      -- 
    ca_5720_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1957_load_0_ack_1, ack => convTransposeB_CP_5119_elements(30)); -- 
    -- CP-element group 31:  join  fork  transition  place  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	22 
    -- CP-element group 31: 	26 
    -- CP-element group 31: 	18 
    -- CP-element group 31: 	12 
    -- CP-element group 31: 	30 
    -- CP-element group 31: 	14 
    -- CP-element group 31: 	28 
    -- CP-element group 31: 	24 
    -- CP-element group 31: 	6 
    -- CP-element group 31: 	8 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	74 
    -- CP-element group 31: 	75 
    -- CP-element group 31: 	73 
    -- CP-element group 31:  members (14) 
      -- CP-element group 31: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964__exit__
      -- CP-element group 31: 	 branch_block_stmt_1825/entry_whilex_xbodyx_xouter
      -- CP-element group 31: 	 branch_block_stmt_1825/assign_stmt_1837_to_assign_stmt_1964/$exit
      -- CP-element group 31: 	 branch_block_stmt_1825/entry_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 31: 	 branch_block_stmt_1825/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1973/$entry
      -- CP-element group 31: 	 branch_block_stmt_1825/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1973/phi_stmt_1973_sources/$entry
      -- CP-element group 31: 	 branch_block_stmt_1825/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1967/$entry
      -- CP-element group 31: 	 branch_block_stmt_1825/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1967/phi_stmt_1967_sources/$entry
      -- CP-element group 31: 	 branch_block_stmt_1825/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1967/phi_stmt_1967_sources/type_cast_1970/$entry
      -- CP-element group 31: 	 branch_block_stmt_1825/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1967/phi_stmt_1967_sources/type_cast_1970/SplitProtocol/$entry
      -- CP-element group 31: 	 branch_block_stmt_1825/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1967/phi_stmt_1967_sources/type_cast_1970/SplitProtocol/Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_1825/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1967/phi_stmt_1967_sources/type_cast_1970/SplitProtocol/Sample/rr
      -- CP-element group 31: 	 branch_block_stmt_1825/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1967/phi_stmt_1967_sources/type_cast_1970/SplitProtocol/Update/$entry
      -- CP-element group 31: 	 branch_block_stmt_1825/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1967/phi_stmt_1967_sources/type_cast_1970/SplitProtocol/Update/cr
      -- 
    rr_6162_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6162_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(31), ack => type_cast_1970_inst_req_0); -- 
    cr_6167_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6167_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(31), ack => type_cast_1970_inst_req_1); -- 
    convTransposeB_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= convTransposeB_CP_5119_elements(22) & convTransposeB_CP_5119_elements(26) & convTransposeB_CP_5119_elements(18) & convTransposeB_CP_5119_elements(12) & convTransposeB_CP_5119_elements(30) & convTransposeB_CP_5119_elements(14) & convTransposeB_CP_5119_elements(28) & convTransposeB_CP_5119_elements(24) & convTransposeB_CP_5119_elements(6) & convTransposeB_CP_5119_elements(8);
      gj_convTransposeB_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5119_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	88 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_1825/assign_stmt_1985_to_assign_stmt_2092/type_cast_1984_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_1825/assign_stmt_1985_to_assign_stmt_2092/type_cast_1984_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_1825/assign_stmt_1985_to_assign_stmt_2092/type_cast_1984_Sample/ra
      -- 
    ra_5737_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1984_inst_ack_0, ack => convTransposeB_CP_5119_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	88 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	36 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_1825/assign_stmt_1985_to_assign_stmt_2092/type_cast_1984_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_1825/assign_stmt_1985_to_assign_stmt_2092/type_cast_1984_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_1825/assign_stmt_1985_to_assign_stmt_2092/type_cast_1984_Update/ca
      -- 
    ca_5742_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1984_inst_ack_1, ack => convTransposeB_CP_5119_elements(33)); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	88 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_1825/assign_stmt_1985_to_assign_stmt_2092/type_cast_1989_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_1825/assign_stmt_1985_to_assign_stmt_2092/type_cast_1989_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_1825/assign_stmt_1985_to_assign_stmt_2092/type_cast_1989_Sample/ra
      -- 
    ra_5751_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1989_inst_ack_0, ack => convTransposeB_CP_5119_elements(34)); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	88 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_1825/assign_stmt_1985_to_assign_stmt_2092/type_cast_1989_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_1825/assign_stmt_1985_to_assign_stmt_2092/type_cast_1989_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_1825/assign_stmt_1985_to_assign_stmt_2092/type_cast_1989_Update/ca
      -- 
    ca_5756_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1989_inst_ack_1, ack => convTransposeB_CP_5119_elements(35)); -- 
    -- CP-element group 36:  join  transition  place  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	33 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	92 
    -- CP-element group 36:  members (6) 
      -- CP-element group 36: 	 branch_block_stmt_1825/assign_stmt_1985_to_assign_stmt_2092__exit__
      -- CP-element group 36: 	 branch_block_stmt_1825/whilex_xbodyx_xouter_whilex_xbody
      -- CP-element group 36: 	 branch_block_stmt_1825/assign_stmt_1985_to_assign_stmt_2092/$exit
      -- CP-element group 36: 	 branch_block_stmt_1825/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$entry
      -- CP-element group 36: 	 branch_block_stmt_1825/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2095/$entry
      -- CP-element group 36: 	 branch_block_stmt_1825/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2095/phi_stmt_2095_sources/$entry
      -- 
    convTransposeB_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5119_elements(33) & convTransposeB_CP_5119_elements(35);
      gj_convTransposeB_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5119_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	94 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/type_cast_2111_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/type_cast_2111_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/type_cast_2111_Sample/ra
      -- 
    ra_5768_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2111_inst_ack_0, ack => convTransposeB_CP_5119_elements(37)); -- 
    -- CP-element group 38:  fork  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	94 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38: 	47 
    -- CP-element group 38:  members (9) 
      -- CP-element group 38: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/type_cast_2111_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/type_cast_2111_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/type_cast_2111_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/type_cast_2141_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/type_cast_2141_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/type_cast_2141_Sample/rr
      -- CP-element group 38: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/type_cast_2172_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/type_cast_2172_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/type_cast_2172_Sample/rr
      -- 
    ca_5773_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2111_inst_ack_1, ack => convTransposeB_CP_5119_elements(38)); -- 
    rr_5781_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5781_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(38), ack => type_cast_2141_inst_req_0); -- 
    rr_5891_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5891_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(38), ack => type_cast_2172_inst_req_0); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/type_cast_2141_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/type_cast_2141_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/type_cast_2141_Sample/ra
      -- 
    ra_5782_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2141_inst_ack_0, ack => convTransposeB_CP_5119_elements(39)); -- 
    -- CP-element group 40:  transition  input  output  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	94 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (16) 
      -- CP-element group 40: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/type_cast_2141_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/type_cast_2141_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/type_cast_2141_Update/ca
      -- CP-element group 40: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/array_obj_ref_2147_index_resized_1
      -- CP-element group 40: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/array_obj_ref_2147_index_scaled_1
      -- CP-element group 40: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/array_obj_ref_2147_index_computed_1
      -- CP-element group 40: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/array_obj_ref_2147_index_resize_1/$entry
      -- CP-element group 40: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/array_obj_ref_2147_index_resize_1/$exit
      -- CP-element group 40: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/array_obj_ref_2147_index_resize_1/index_resize_req
      -- CP-element group 40: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/array_obj_ref_2147_index_resize_1/index_resize_ack
      -- CP-element group 40: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/array_obj_ref_2147_index_scale_1/$entry
      -- CP-element group 40: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/array_obj_ref_2147_index_scale_1/$exit
      -- CP-element group 40: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/array_obj_ref_2147_index_scale_1/scale_rename_req
      -- CP-element group 40: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/array_obj_ref_2147_index_scale_1/scale_rename_ack
      -- CP-element group 40: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/array_obj_ref_2147_final_index_sum_regn_Sample/$entry
      -- CP-element group 40: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/array_obj_ref_2147_final_index_sum_regn_Sample/req
      -- 
    ca_5787_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2141_inst_ack_1, ack => convTransposeB_CP_5119_elements(40)); -- 
    req_5812_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5812_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(40), ack => array_obj_ref_2147_index_offset_req_0); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	58 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/array_obj_ref_2147_final_index_sum_regn_sample_complete
      -- CP-element group 41: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/array_obj_ref_2147_final_index_sum_regn_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/array_obj_ref_2147_final_index_sum_regn_Sample/ack
      -- 
    ack_5813_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2147_index_offset_ack_0, ack => convTransposeB_CP_5119_elements(41)); -- 
    -- CP-element group 42:  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	94 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (11) 
      -- CP-element group 42: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/addr_of_2148_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/array_obj_ref_2147_root_address_calculated
      -- CP-element group 42: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/array_obj_ref_2147_offset_calculated
      -- CP-element group 42: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/array_obj_ref_2147_final_index_sum_regn_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/array_obj_ref_2147_final_index_sum_regn_Update/ack
      -- CP-element group 42: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/array_obj_ref_2147_base_plus_offset/$entry
      -- CP-element group 42: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/array_obj_ref_2147_base_plus_offset/$exit
      -- CP-element group 42: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/array_obj_ref_2147_base_plus_offset/sum_rename_req
      -- CP-element group 42: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/array_obj_ref_2147_base_plus_offset/sum_rename_ack
      -- CP-element group 42: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/addr_of_2148_request/$entry
      -- CP-element group 42: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/addr_of_2148_request/req
      -- 
    ack_5818_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2147_index_offset_ack_1, ack => convTransposeB_CP_5119_elements(42)); -- 
    req_5827_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5827_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(42), ack => addr_of_2148_final_reg_req_0); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/addr_of_2148_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/addr_of_2148_request/$exit
      -- CP-element group 43: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/addr_of_2148_request/ack
      -- 
    ack_5828_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2148_final_reg_ack_0, ack => convTransposeB_CP_5119_elements(43)); -- 
    -- CP-element group 44:  join  fork  transition  input  output  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	94 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (24) 
      -- CP-element group 44: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/addr_of_2148_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/addr_of_2148_complete/$exit
      -- CP-element group 44: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/addr_of_2148_complete/ack
      -- CP-element group 44: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2152_sample_start_
      -- CP-element group 44: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2152_base_address_calculated
      -- CP-element group 44: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2152_word_address_calculated
      -- CP-element group 44: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2152_root_address_calculated
      -- CP-element group 44: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2152_base_address_resized
      -- CP-element group 44: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2152_base_addr_resize/$entry
      -- CP-element group 44: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2152_base_addr_resize/$exit
      -- CP-element group 44: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2152_base_addr_resize/base_resize_req
      -- CP-element group 44: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2152_base_addr_resize/base_resize_ack
      -- CP-element group 44: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2152_base_plus_offset/$entry
      -- CP-element group 44: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2152_base_plus_offset/$exit
      -- CP-element group 44: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2152_base_plus_offset/sum_rename_req
      -- CP-element group 44: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2152_base_plus_offset/sum_rename_ack
      -- CP-element group 44: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2152_word_addrgen/$entry
      -- CP-element group 44: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2152_word_addrgen/$exit
      -- CP-element group 44: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2152_word_addrgen/root_register_req
      -- CP-element group 44: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2152_word_addrgen/root_register_ack
      -- CP-element group 44: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2152_Sample/$entry
      -- CP-element group 44: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2152_Sample/word_access_start/$entry
      -- CP-element group 44: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2152_Sample/word_access_start/word_0/$entry
      -- CP-element group 44: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2152_Sample/word_access_start/word_0/rr
      -- 
    ack_5833_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2148_final_reg_ack_1, ack => convTransposeB_CP_5119_elements(44)); -- 
    rr_5866_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5866_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(44), ack => ptr_deref_2152_load_0_req_0); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	44 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (5) 
      -- CP-element group 45: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2152_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2152_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2152_Sample/word_access_start/$exit
      -- CP-element group 45: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2152_Sample/word_access_start/word_0/$exit
      -- CP-element group 45: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2152_Sample/word_access_start/word_0/ra
      -- 
    ra_5867_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2152_load_0_ack_0, ack => convTransposeB_CP_5119_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	94 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	53 
    -- CP-element group 46:  members (9) 
      -- CP-element group 46: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2152_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2152_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2152_Update/word_access_complete/$exit
      -- CP-element group 46: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2152_Update/word_access_complete/word_0/$exit
      -- CP-element group 46: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2152_Update/word_access_complete/word_0/ca
      -- CP-element group 46: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2152_Update/ptr_deref_2152_Merge/$entry
      -- CP-element group 46: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2152_Update/ptr_deref_2152_Merge/$exit
      -- CP-element group 46: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2152_Update/ptr_deref_2152_Merge/merge_req
      -- CP-element group 46: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2152_Update/ptr_deref_2152_Merge/merge_ack
      -- 
    ca_5878_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2152_load_0_ack_1, ack => convTransposeB_CP_5119_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	38 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/type_cast_2172_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/type_cast_2172_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/type_cast_2172_Sample/ra
      -- 
    ra_5892_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2172_inst_ack_0, ack => convTransposeB_CP_5119_elements(47)); -- 
    -- CP-element group 48:  transition  input  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	94 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (16) 
      -- CP-element group 48: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/type_cast_2172_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/type_cast_2172_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/type_cast_2172_Update/ca
      -- CP-element group 48: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/array_obj_ref_2178_index_resized_1
      -- CP-element group 48: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/array_obj_ref_2178_index_scaled_1
      -- CP-element group 48: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/array_obj_ref_2178_index_computed_1
      -- CP-element group 48: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/array_obj_ref_2178_index_resize_1/$entry
      -- CP-element group 48: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/array_obj_ref_2178_index_resize_1/$exit
      -- CP-element group 48: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/array_obj_ref_2178_index_resize_1/index_resize_req
      -- CP-element group 48: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/array_obj_ref_2178_index_resize_1/index_resize_ack
      -- CP-element group 48: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/array_obj_ref_2178_index_scale_1/$entry
      -- CP-element group 48: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/array_obj_ref_2178_index_scale_1/$exit
      -- CP-element group 48: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/array_obj_ref_2178_index_scale_1/scale_rename_req
      -- CP-element group 48: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/array_obj_ref_2178_index_scale_1/scale_rename_ack
      -- CP-element group 48: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/array_obj_ref_2178_final_index_sum_regn_Sample/$entry
      -- CP-element group 48: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/array_obj_ref_2178_final_index_sum_regn_Sample/req
      -- 
    ca_5897_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2172_inst_ack_1, ack => convTransposeB_CP_5119_elements(48)); -- 
    req_5922_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5922_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(48), ack => array_obj_ref_2178_index_offset_req_0); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	58 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/array_obj_ref_2178_final_index_sum_regn_sample_complete
      -- CP-element group 49: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/array_obj_ref_2178_final_index_sum_regn_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/array_obj_ref_2178_final_index_sum_regn_Sample/ack
      -- 
    ack_5923_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2178_index_offset_ack_0, ack => convTransposeB_CP_5119_elements(49)); -- 
    -- CP-element group 50:  transition  input  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	94 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (11) 
      -- CP-element group 50: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/addr_of_2179_request/$entry
      -- CP-element group 50: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/addr_of_2179_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/array_obj_ref_2178_root_address_calculated
      -- CP-element group 50: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/array_obj_ref_2178_offset_calculated
      -- CP-element group 50: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/array_obj_ref_2178_final_index_sum_regn_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/array_obj_ref_2178_final_index_sum_regn_Update/ack
      -- CP-element group 50: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/array_obj_ref_2178_base_plus_offset/$entry
      -- CP-element group 50: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/array_obj_ref_2178_base_plus_offset/$exit
      -- CP-element group 50: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/array_obj_ref_2178_base_plus_offset/sum_rename_req
      -- CP-element group 50: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/array_obj_ref_2178_base_plus_offset/sum_rename_ack
      -- CP-element group 50: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/addr_of_2179_request/req
      -- 
    ack_5928_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2178_index_offset_ack_1, ack => convTransposeB_CP_5119_elements(50)); -- 
    req_5937_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5937_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(50), ack => addr_of_2179_final_reg_req_0); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/addr_of_2179_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/addr_of_2179_request/$exit
      -- CP-element group 51: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/addr_of_2179_request/ack
      -- 
    ack_5938_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2179_final_reg_ack_0, ack => convTransposeB_CP_5119_elements(51)); -- 
    -- CP-element group 52:  fork  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	94 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	53 
    -- CP-element group 52:  members (19) 
      -- CP-element group 52: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/addr_of_2179_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/addr_of_2179_complete/$exit
      -- CP-element group 52: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/addr_of_2179_complete/ack
      -- CP-element group 52: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2182_base_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2182_word_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2182_root_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2182_base_address_resized
      -- CP-element group 52: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2182_base_addr_resize/$entry
      -- CP-element group 52: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2182_base_addr_resize/$exit
      -- CP-element group 52: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2182_base_addr_resize/base_resize_req
      -- CP-element group 52: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2182_base_addr_resize/base_resize_ack
      -- CP-element group 52: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2182_base_plus_offset/$entry
      -- CP-element group 52: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2182_base_plus_offset/$exit
      -- CP-element group 52: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2182_base_plus_offset/sum_rename_req
      -- CP-element group 52: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2182_base_plus_offset/sum_rename_ack
      -- CP-element group 52: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2182_word_addrgen/$entry
      -- CP-element group 52: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2182_word_addrgen/$exit
      -- CP-element group 52: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2182_word_addrgen/root_register_req
      -- CP-element group 52: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2182_word_addrgen/root_register_ack
      -- 
    ack_5943_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2179_final_reg_ack_1, ack => convTransposeB_CP_5119_elements(52)); -- 
    -- CP-element group 53:  join  transition  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	46 
    -- CP-element group 53: 	52 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (9) 
      -- CP-element group 53: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2182_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2182_Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2182_Sample/ptr_deref_2182_Split/$entry
      -- CP-element group 53: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2182_Sample/ptr_deref_2182_Split/$exit
      -- CP-element group 53: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2182_Sample/ptr_deref_2182_Split/split_req
      -- CP-element group 53: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2182_Sample/ptr_deref_2182_Split/split_ack
      -- CP-element group 53: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2182_Sample/word_access_start/$entry
      -- CP-element group 53: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2182_Sample/word_access_start/word_0/$entry
      -- CP-element group 53: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2182_Sample/word_access_start/word_0/rr
      -- 
    rr_5981_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5981_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(53), ack => ptr_deref_2182_store_0_req_0); -- 
    convTransposeB_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5119_elements(46) & convTransposeB_CP_5119_elements(52);
      gj_convTransposeB_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5119_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (5) 
      -- CP-element group 54: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2182_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2182_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2182_Sample/word_access_start/$exit
      -- CP-element group 54: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2182_Sample/word_access_start/word_0/$exit
      -- CP-element group 54: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2182_Sample/word_access_start/word_0/ra
      -- 
    ra_5982_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2182_store_0_ack_0, ack => convTransposeB_CP_5119_elements(54)); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	94 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	58 
    -- CP-element group 55:  members (5) 
      -- CP-element group 55: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2182_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2182_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2182_Update/word_access_complete/$exit
      -- CP-element group 55: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2182_Update/word_access_complete/word_0/$exit
      -- CP-element group 55: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2182_Update/word_access_complete/word_0/ca
      -- 
    ca_5993_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2182_store_0_ack_1, ack => convTransposeB_CP_5119_elements(55)); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	94 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/type_cast_2188_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/type_cast_2188_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/type_cast_2188_Sample/ra
      -- 
    ra_6002_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2188_inst_ack_0, ack => convTransposeB_CP_5119_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	94 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/type_cast_2188_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/type_cast_2188_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/type_cast_2188_Update/ca
      -- 
    ca_6007_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2188_inst_ack_1, ack => convTransposeB_CP_5119_elements(57)); -- 
    -- CP-element group 58:  branch  join  transition  place  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	41 
    -- CP-element group 58: 	55 
    -- CP-element group 58: 	57 
    -- CP-element group 58: 	49 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	60 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (10) 
      -- CP-element group 58: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200__exit__
      -- CP-element group 58: 	 branch_block_stmt_1825/if_stmt_2201__entry__
      -- CP-element group 58: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/$exit
      -- CP-element group 58: 	 branch_block_stmt_1825/if_stmt_2201_dead_link/$entry
      -- CP-element group 58: 	 branch_block_stmt_1825/if_stmt_2201_eval_test/$entry
      -- CP-element group 58: 	 branch_block_stmt_1825/if_stmt_2201_eval_test/$exit
      -- CP-element group 58: 	 branch_block_stmt_1825/if_stmt_2201_eval_test/branch_req
      -- CP-element group 58: 	 branch_block_stmt_1825/R_cmp_2202_place
      -- CP-element group 58: 	 branch_block_stmt_1825/if_stmt_2201_if_link/$entry
      -- CP-element group 58: 	 branch_block_stmt_1825/if_stmt_2201_else_link/$entry
      -- 
    branch_req_6015_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6015_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(58), ack => if_stmt_2201_branch_req_0); -- 
    convTransposeB_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_5119_elements(41) & convTransposeB_CP_5119_elements(55) & convTransposeB_CP_5119_elements(57) & convTransposeB_CP_5119_elements(49);
      gj_convTransposeB_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5119_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	90 
    -- CP-element group 59: 	89 
    -- CP-element group 59:  members (24) 
      -- CP-element group 59: 	 branch_block_stmt_1825/merge_stmt_2207__exit__
      -- CP-element group 59: 	 branch_block_stmt_1825/assign_stmt_2213__entry__
      -- CP-element group 59: 	 branch_block_stmt_1825/assign_stmt_2213__exit__
      -- CP-element group 59: 	 branch_block_stmt_1825/ifx_xthen_whilex_xbody
      -- CP-element group 59: 	 branch_block_stmt_1825/if_stmt_2201_if_link/$exit
      -- CP-element group 59: 	 branch_block_stmt_1825/if_stmt_2201_if_link/if_choice_transition
      -- CP-element group 59: 	 branch_block_stmt_1825/whilex_xbody_ifx_xthen
      -- CP-element group 59: 	 branch_block_stmt_1825/assign_stmt_2213/$entry
      -- CP-element group 59: 	 branch_block_stmt_1825/assign_stmt_2213/$exit
      -- CP-element group 59: 	 branch_block_stmt_1825/ifx_xthen_whilex_xbody_PhiReq/$entry
      -- CP-element group 59: 	 branch_block_stmt_1825/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2095/$entry
      -- CP-element group 59: 	 branch_block_stmt_1825/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2095/phi_stmt_2095_sources/$entry
      -- CP-element group 59: 	 branch_block_stmt_1825/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2095/phi_stmt_2095_sources/type_cast_2101/$entry
      -- CP-element group 59: 	 branch_block_stmt_1825/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2095/phi_stmt_2095_sources/type_cast_2101/SplitProtocol/$entry
      -- CP-element group 59: 	 branch_block_stmt_1825/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2095/phi_stmt_2095_sources/type_cast_2101/SplitProtocol/Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_1825/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2095/phi_stmt_2095_sources/type_cast_2101/SplitProtocol/Sample/rr
      -- CP-element group 59: 	 branch_block_stmt_1825/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2095/phi_stmt_2095_sources/type_cast_2101/SplitProtocol/Update/$entry
      -- CP-element group 59: 	 branch_block_stmt_1825/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2095/phi_stmt_2095_sources/type_cast_2101/SplitProtocol/Update/cr
      -- CP-element group 59: 	 branch_block_stmt_1825/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 59: 	 branch_block_stmt_1825/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 59: 	 branch_block_stmt_1825/merge_stmt_2207_PhiReqMerge
      -- CP-element group 59: 	 branch_block_stmt_1825/merge_stmt_2207_PhiAck/$entry
      -- CP-element group 59: 	 branch_block_stmt_1825/merge_stmt_2207_PhiAck/$exit
      -- CP-element group 59: 	 branch_block_stmt_1825/merge_stmt_2207_PhiAck/dummy
      -- 
    if_choice_transition_6020_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2201_branch_ack_1, ack => convTransposeB_CP_5119_elements(59)); -- 
    rr_6243_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6243_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(59), ack => type_cast_2101_inst_req_0); -- 
    cr_6248_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6248_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(59), ack => type_cast_2101_inst_req_1); -- 
    -- CP-element group 60:  fork  transition  place  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	58 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60: 	62 
    -- CP-element group 60:  members (18) 
      -- CP-element group 60: 	 branch_block_stmt_1825/merge_stmt_2215__exit__
      -- CP-element group 60: 	 branch_block_stmt_1825/assign_stmt_2221_to_assign_stmt_2231__entry__
      -- CP-element group 60: 	 branch_block_stmt_1825/if_stmt_2201_else_link/$exit
      -- CP-element group 60: 	 branch_block_stmt_1825/if_stmt_2201_else_link/else_choice_transition
      -- CP-element group 60: 	 branch_block_stmt_1825/whilex_xbody_ifx_xelse
      -- CP-element group 60: 	 branch_block_stmt_1825/assign_stmt_2221_to_assign_stmt_2231/$entry
      -- CP-element group 60: 	 branch_block_stmt_1825/assign_stmt_2221_to_assign_stmt_2231/type_cast_2225_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_1825/assign_stmt_2221_to_assign_stmt_2231/type_cast_2225_update_start_
      -- CP-element group 60: 	 branch_block_stmt_1825/assign_stmt_2221_to_assign_stmt_2231/type_cast_2225_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_1825/assign_stmt_2221_to_assign_stmt_2231/type_cast_2225_Sample/rr
      -- CP-element group 60: 	 branch_block_stmt_1825/assign_stmt_2221_to_assign_stmt_2231/type_cast_2225_Update/$entry
      -- CP-element group 60: 	 branch_block_stmt_1825/assign_stmt_2221_to_assign_stmt_2231/type_cast_2225_Update/cr
      -- CP-element group 60: 	 branch_block_stmt_1825/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 60: 	 branch_block_stmt_1825/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 60: 	 branch_block_stmt_1825/merge_stmt_2215_PhiReqMerge
      -- CP-element group 60: 	 branch_block_stmt_1825/merge_stmt_2215_PhiAck/$entry
      -- CP-element group 60: 	 branch_block_stmt_1825/merge_stmt_2215_PhiAck/$exit
      -- CP-element group 60: 	 branch_block_stmt_1825/merge_stmt_2215_PhiAck/dummy
      -- 
    else_choice_transition_6024_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2201_branch_ack_0, ack => convTransposeB_CP_5119_elements(60)); -- 
    rr_6040_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6040_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(60), ack => type_cast_2225_inst_req_0); -- 
    cr_6045_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6045_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(60), ack => type_cast_2225_inst_req_1); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_1825/assign_stmt_2221_to_assign_stmt_2231/type_cast_2225_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_1825/assign_stmt_2221_to_assign_stmt_2231/type_cast_2225_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_1825/assign_stmt_2221_to_assign_stmt_2231/type_cast_2225_Sample/ra
      -- 
    ra_6041_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2225_inst_ack_0, ack => convTransposeB_CP_5119_elements(61)); -- 
    -- CP-element group 62:  branch  transition  place  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	60 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62: 	64 
    -- CP-element group 62:  members (13) 
      -- CP-element group 62: 	 branch_block_stmt_1825/assign_stmt_2221_to_assign_stmt_2231__exit__
      -- CP-element group 62: 	 branch_block_stmt_1825/if_stmt_2232__entry__
      -- CP-element group 62: 	 branch_block_stmt_1825/assign_stmt_2221_to_assign_stmt_2231/$exit
      -- CP-element group 62: 	 branch_block_stmt_1825/assign_stmt_2221_to_assign_stmt_2231/type_cast_2225_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_1825/assign_stmt_2221_to_assign_stmt_2231/type_cast_2225_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_1825/assign_stmt_2221_to_assign_stmt_2231/type_cast_2225_Update/ca
      -- CP-element group 62: 	 branch_block_stmt_1825/if_stmt_2232_dead_link/$entry
      -- CP-element group 62: 	 branch_block_stmt_1825/if_stmt_2232_eval_test/$entry
      -- CP-element group 62: 	 branch_block_stmt_1825/if_stmt_2232_eval_test/$exit
      -- CP-element group 62: 	 branch_block_stmt_1825/if_stmt_2232_eval_test/branch_req
      -- CP-element group 62: 	 branch_block_stmt_1825/R_cmp77_2233_place
      -- CP-element group 62: 	 branch_block_stmt_1825/if_stmt_2232_if_link/$entry
      -- CP-element group 62: 	 branch_block_stmt_1825/if_stmt_2232_else_link/$entry
      -- 
    ca_6046_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2225_inst_ack_1, ack => convTransposeB_CP_5119_elements(62)); -- 
    branch_req_6054_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6054_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(62), ack => if_stmt_2232_branch_req_0); -- 
    -- CP-element group 63:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	65 
    -- CP-element group 63: 	66 
    -- CP-element group 63:  members (18) 
      -- CP-element group 63: 	 branch_block_stmt_1825/merge_stmt_2238__exit__
      -- CP-element group 63: 	 branch_block_stmt_1825/assign_stmt_2244_to_assign_stmt_2254__entry__
      -- CP-element group 63: 	 branch_block_stmt_1825/if_stmt_2232_if_link/$exit
      -- CP-element group 63: 	 branch_block_stmt_1825/if_stmt_2232_if_link/if_choice_transition
      -- CP-element group 63: 	 branch_block_stmt_1825/ifx_xelse_ifx_xthen79
      -- CP-element group 63: 	 branch_block_stmt_1825/assign_stmt_2244_to_assign_stmt_2254/$entry
      -- CP-element group 63: 	 branch_block_stmt_1825/assign_stmt_2244_to_assign_stmt_2254/type_cast_2253_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_1825/assign_stmt_2244_to_assign_stmt_2254/type_cast_2253_update_start_
      -- CP-element group 63: 	 branch_block_stmt_1825/assign_stmt_2244_to_assign_stmt_2254/type_cast_2253_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_1825/assign_stmt_2244_to_assign_stmt_2254/type_cast_2253_Sample/rr
      -- CP-element group 63: 	 branch_block_stmt_1825/assign_stmt_2244_to_assign_stmt_2254/type_cast_2253_Update/$entry
      -- CP-element group 63: 	 branch_block_stmt_1825/assign_stmt_2244_to_assign_stmt_2254/type_cast_2253_Update/cr
      -- CP-element group 63: 	 branch_block_stmt_1825/ifx_xelse_ifx_xthen79_PhiReq/$entry
      -- CP-element group 63: 	 branch_block_stmt_1825/ifx_xelse_ifx_xthen79_PhiReq/$exit
      -- CP-element group 63: 	 branch_block_stmt_1825/merge_stmt_2238_PhiReqMerge
      -- CP-element group 63: 	 branch_block_stmt_1825/merge_stmt_2238_PhiAck/$entry
      -- CP-element group 63: 	 branch_block_stmt_1825/merge_stmt_2238_PhiAck/$exit
      -- CP-element group 63: 	 branch_block_stmt_1825/merge_stmt_2238_PhiAck/dummy
      -- 
    if_choice_transition_6059_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2232_branch_ack_1, ack => convTransposeB_CP_5119_elements(63)); -- 
    rr_6076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(63), ack => type_cast_2253_inst_req_0); -- 
    cr_6081_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6081_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(63), ack => type_cast_2253_inst_req_1); -- 
    -- CP-element group 64:  fork  transition  place  input  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	62 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	96 
    -- CP-element group 64: 	98 
    -- CP-element group 64: 	99 
    -- CP-element group 64: 	95 
    -- CP-element group 64:  members (20) 
      -- CP-element group 64: 	 branch_block_stmt_1825/if_stmt_2232_else_link/$exit
      -- CP-element group 64: 	 branch_block_stmt_1825/if_stmt_2232_else_link/else_choice_transition
      -- CP-element group 64: 	 branch_block_stmt_1825/ifx_xelse_ifx_xend
      -- CP-element group 64: 	 branch_block_stmt_1825/ifx_xelse_ifx_xend_PhiReq/$entry
      -- CP-element group 64: 	 branch_block_stmt_1825/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2257/$entry
      -- CP-element group 64: 	 branch_block_stmt_1825/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2257/phi_stmt_2257_sources/$entry
      -- CP-element group 64: 	 branch_block_stmt_1825/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2257/phi_stmt_2257_sources/type_cast_2262/$entry
      -- CP-element group 64: 	 branch_block_stmt_1825/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2257/phi_stmt_2257_sources/type_cast_2262/SplitProtocol/$entry
      -- CP-element group 64: 	 branch_block_stmt_1825/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2257/phi_stmt_2257_sources/type_cast_2262/SplitProtocol/Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_1825/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2257/phi_stmt_2257_sources/type_cast_2262/SplitProtocol/Sample/rr
      -- CP-element group 64: 	 branch_block_stmt_1825/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2257/phi_stmt_2257_sources/type_cast_2262/SplitProtocol/Update/$entry
      -- CP-element group 64: 	 branch_block_stmt_1825/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2257/phi_stmt_2257_sources/type_cast_2262/SplitProtocol/Update/cr
      -- CP-element group 64: 	 branch_block_stmt_1825/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2263/$entry
      -- CP-element group 64: 	 branch_block_stmt_1825/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2263/phi_stmt_2263_sources/$entry
      -- CP-element group 64: 	 branch_block_stmt_1825/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2263/phi_stmt_2263_sources/type_cast_2268/$entry
      -- CP-element group 64: 	 branch_block_stmt_1825/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2263/phi_stmt_2263_sources/type_cast_2268/SplitProtocol/$entry
      -- CP-element group 64: 	 branch_block_stmt_1825/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2263/phi_stmt_2263_sources/type_cast_2268/SplitProtocol/Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_1825/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2263/phi_stmt_2263_sources/type_cast_2268/SplitProtocol/Sample/rr
      -- CP-element group 64: 	 branch_block_stmt_1825/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2263/phi_stmt_2263_sources/type_cast_2268/SplitProtocol/Update/$entry
      -- CP-element group 64: 	 branch_block_stmt_1825/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2263/phi_stmt_2263_sources/type_cast_2268/SplitProtocol/Update/cr
      -- 
    else_choice_transition_6063_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2232_branch_ack_0, ack => convTransposeB_CP_5119_elements(64)); -- 
    rr_6317_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6317_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(64), ack => type_cast_2262_inst_req_0); -- 
    cr_6322_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6322_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(64), ack => type_cast_2262_inst_req_1); -- 
    rr_6340_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6340_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(64), ack => type_cast_2268_inst_req_0); -- 
    cr_6345_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6345_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(64), ack => type_cast_2268_inst_req_1); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_1825/assign_stmt_2244_to_assign_stmt_2254/type_cast_2253_sample_completed_
      -- CP-element group 65: 	 branch_block_stmt_1825/assign_stmt_2244_to_assign_stmt_2254/type_cast_2253_Sample/$exit
      -- CP-element group 65: 	 branch_block_stmt_1825/assign_stmt_2244_to_assign_stmt_2254/type_cast_2253_Sample/ra
      -- 
    ra_6077_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2253_inst_ack_0, ack => convTransposeB_CP_5119_elements(65)); -- 
    -- CP-element group 66:  fork  transition  place  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	63 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	102 
    -- CP-element group 66: 	105 
    -- CP-element group 66: 	106 
    -- CP-element group 66: 	103 
    -- CP-element group 66:  members (23) 
      -- CP-element group 66: 	 branch_block_stmt_1825/assign_stmt_2244_to_assign_stmt_2254__exit__
      -- CP-element group 66: 	 branch_block_stmt_1825/ifx_xthen79_ifx_xend
      -- CP-element group 66: 	 branch_block_stmt_1825/assign_stmt_2244_to_assign_stmt_2254/$exit
      -- CP-element group 66: 	 branch_block_stmt_1825/assign_stmt_2244_to_assign_stmt_2254/type_cast_2253_update_completed_
      -- CP-element group 66: 	 branch_block_stmt_1825/assign_stmt_2244_to_assign_stmt_2254/type_cast_2253_Update/$exit
      -- CP-element group 66: 	 branch_block_stmt_1825/assign_stmt_2244_to_assign_stmt_2254/type_cast_2253_Update/ca
      -- CP-element group 66: 	 branch_block_stmt_1825/ifx_xthen79_ifx_xend_PhiReq/$entry
      -- CP-element group 66: 	 branch_block_stmt_1825/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2257/$entry
      -- CP-element group 66: 	 branch_block_stmt_1825/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2257/phi_stmt_2257_sources/$entry
      -- CP-element group 66: 	 branch_block_stmt_1825/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2257/phi_stmt_2257_sources/type_cast_2260/$entry
      -- CP-element group 66: 	 branch_block_stmt_1825/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2257/phi_stmt_2257_sources/type_cast_2260/SplitProtocol/$entry
      -- CP-element group 66: 	 branch_block_stmt_1825/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2257/phi_stmt_2257_sources/type_cast_2260/SplitProtocol/Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_1825/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2257/phi_stmt_2257_sources/type_cast_2260/SplitProtocol/Sample/rr
      -- CP-element group 66: 	 branch_block_stmt_1825/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2257/phi_stmt_2257_sources/type_cast_2260/SplitProtocol/Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_1825/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2257/phi_stmt_2257_sources/type_cast_2260/SplitProtocol/Update/cr
      -- CP-element group 66: 	 branch_block_stmt_1825/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2263/$entry
      -- CP-element group 66: 	 branch_block_stmt_1825/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2263/phi_stmt_2263_sources/$entry
      -- CP-element group 66: 	 branch_block_stmt_1825/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2263/phi_stmt_2263_sources/type_cast_2266/$entry
      -- CP-element group 66: 	 branch_block_stmt_1825/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2263/phi_stmt_2263_sources/type_cast_2266/SplitProtocol/$entry
      -- CP-element group 66: 	 branch_block_stmt_1825/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2263/phi_stmt_2263_sources/type_cast_2266/SplitProtocol/Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_1825/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2263/phi_stmt_2263_sources/type_cast_2266/SplitProtocol/Sample/rr
      -- CP-element group 66: 	 branch_block_stmt_1825/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2263/phi_stmt_2263_sources/type_cast_2266/SplitProtocol/Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_1825/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2263/phi_stmt_2263_sources/type_cast_2266/SplitProtocol/Update/cr
      -- 
    ca_6082_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2253_inst_ack_1, ack => convTransposeB_CP_5119_elements(66)); -- 
    rr_6366_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6366_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(66), ack => type_cast_2260_inst_req_0); -- 
    cr_6371_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6371_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(66), ack => type_cast_2260_inst_req_1); -- 
    rr_6389_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6389_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(66), ack => type_cast_2266_inst_req_0); -- 
    cr_6394_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6394_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(66), ack => type_cast_2266_inst_req_1); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	112 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_1825/assign_stmt_2274_to_assign_stmt_2279/type_cast_2273_sample_completed_
      -- CP-element group 67: 	 branch_block_stmt_1825/assign_stmt_2274_to_assign_stmt_2279/type_cast_2273_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_1825/assign_stmt_2274_to_assign_stmt_2279/type_cast_2273_Sample/ra
      -- 
    ra_6094_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2273_inst_ack_0, ack => convTransposeB_CP_5119_elements(67)); -- 
    -- CP-element group 68:  branch  transition  place  input  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	112 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (13) 
      -- CP-element group 68: 	 branch_block_stmt_1825/assign_stmt_2274_to_assign_stmt_2279__exit__
      -- CP-element group 68: 	 branch_block_stmt_1825/if_stmt_2280__entry__
      -- CP-element group 68: 	 branch_block_stmt_1825/assign_stmt_2274_to_assign_stmt_2279/$exit
      -- CP-element group 68: 	 branch_block_stmt_1825/assign_stmt_2274_to_assign_stmt_2279/type_cast_2273_update_completed_
      -- CP-element group 68: 	 branch_block_stmt_1825/assign_stmt_2274_to_assign_stmt_2279/type_cast_2273_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_1825/assign_stmt_2274_to_assign_stmt_2279/type_cast_2273_Update/ca
      -- CP-element group 68: 	 branch_block_stmt_1825/if_stmt_2280_dead_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_1825/if_stmt_2280_eval_test/$entry
      -- CP-element group 68: 	 branch_block_stmt_1825/if_stmt_2280_eval_test/$exit
      -- CP-element group 68: 	 branch_block_stmt_1825/if_stmt_2280_eval_test/branch_req
      -- CP-element group 68: 	 branch_block_stmt_1825/R_cmp89_2281_place
      -- CP-element group 68: 	 branch_block_stmt_1825/if_stmt_2280_if_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_1825/if_stmt_2280_else_link/$entry
      -- 
    ca_6099_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2273_inst_ack_1, ack => convTransposeB_CP_5119_elements(68)); -- 
    branch_req_6107_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6107_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(68), ack => if_stmt_2280_branch_req_0); -- 
    -- CP-element group 69:  merge  transition  place  input  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	71 
    -- CP-element group 69:  members (15) 
      -- CP-element group 69: 	 branch_block_stmt_1825/merge_stmt_2286__exit__
      -- CP-element group 69: 	 branch_block_stmt_1825/assign_stmt_2290__entry__
      -- CP-element group 69: 	 branch_block_stmt_1825/if_stmt_2280_if_link/$exit
      -- CP-element group 69: 	 branch_block_stmt_1825/if_stmt_2280_if_link/if_choice_transition
      -- CP-element group 69: 	 branch_block_stmt_1825/ifx_xend_whilex_xend
      -- CP-element group 69: 	 branch_block_stmt_1825/assign_stmt_2290/$entry
      -- CP-element group 69: 	 branch_block_stmt_1825/assign_stmt_2290/WPIPE_Block1_done_2288_sample_start_
      -- CP-element group 69: 	 branch_block_stmt_1825/assign_stmt_2290/WPIPE_Block1_done_2288_Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_1825/assign_stmt_2290/WPIPE_Block1_done_2288_Sample/req
      -- CP-element group 69: 	 branch_block_stmt_1825/ifx_xend_whilex_xend_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_1825/ifx_xend_whilex_xend_PhiReq/$exit
      -- CP-element group 69: 	 branch_block_stmt_1825/merge_stmt_2286_PhiReqMerge
      -- CP-element group 69: 	 branch_block_stmt_1825/merge_stmt_2286_PhiAck/$entry
      -- CP-element group 69: 	 branch_block_stmt_1825/merge_stmt_2286_PhiAck/$exit
      -- CP-element group 69: 	 branch_block_stmt_1825/merge_stmt_2286_PhiAck/dummy
      -- 
    if_choice_transition_6112_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2280_branch_ack_1, ack => convTransposeB_CP_5119_elements(69)); -- 
    req_6129_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6129_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(69), ack => WPIPE_Block1_done_2288_inst_req_0); -- 
    -- CP-element group 70:  fork  transition  place  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	78 
    -- CP-element group 70: 	79 
    -- CP-element group 70: 	81 
    -- CP-element group 70: 	82 
    -- CP-element group 70:  members (20) 
      -- CP-element group 70: 	 branch_block_stmt_1825/if_stmt_2280_else_link/$exit
      -- CP-element group 70: 	 branch_block_stmt_1825/if_stmt_2280_else_link/else_choice_transition
      -- CP-element group 70: 	 branch_block_stmt_1825/ifx_xend_whilex_xbodyx_xouter
      -- CP-element group 70: 	 branch_block_stmt_1825/ifx_xend_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 70: 	 branch_block_stmt_1825/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1973/$entry
      -- CP-element group 70: 	 branch_block_stmt_1825/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1973/phi_stmt_1973_sources/$entry
      -- CP-element group 70: 	 branch_block_stmt_1825/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1973/phi_stmt_1973_sources/type_cast_1979/$entry
      -- CP-element group 70: 	 branch_block_stmt_1825/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1973/phi_stmt_1973_sources/type_cast_1979/SplitProtocol/$entry
      -- CP-element group 70: 	 branch_block_stmt_1825/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1973/phi_stmt_1973_sources/type_cast_1979/SplitProtocol/Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_1825/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1973/phi_stmt_1973_sources/type_cast_1979/SplitProtocol/Sample/rr
      -- CP-element group 70: 	 branch_block_stmt_1825/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1973/phi_stmt_1973_sources/type_cast_1979/SplitProtocol/Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_1825/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1973/phi_stmt_1973_sources/type_cast_1979/SplitProtocol/Update/cr
      -- CP-element group 70: 	 branch_block_stmt_1825/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1967/$entry
      -- CP-element group 70: 	 branch_block_stmt_1825/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1967/phi_stmt_1967_sources/$entry
      -- CP-element group 70: 	 branch_block_stmt_1825/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1967/phi_stmt_1967_sources/type_cast_1972/$entry
      -- CP-element group 70: 	 branch_block_stmt_1825/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1967/phi_stmt_1967_sources/type_cast_1972/SplitProtocol/$entry
      -- CP-element group 70: 	 branch_block_stmt_1825/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1967/phi_stmt_1967_sources/type_cast_1972/SplitProtocol/Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_1825/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1967/phi_stmt_1967_sources/type_cast_1972/SplitProtocol/Sample/rr
      -- CP-element group 70: 	 branch_block_stmt_1825/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1967/phi_stmt_1967_sources/type_cast_1972/SplitProtocol/Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_1825/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1967/phi_stmt_1967_sources/type_cast_1972/SplitProtocol/Update/cr
      -- 
    else_choice_transition_6116_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2280_branch_ack_0, ack => convTransposeB_CP_5119_elements(70)); -- 
    rr_6188_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6188_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(70), ack => type_cast_1979_inst_req_0); -- 
    cr_6193_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6193_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(70), ack => type_cast_1979_inst_req_1); -- 
    rr_6211_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6211_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(70), ack => type_cast_1972_inst_req_0); -- 
    cr_6216_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6216_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(70), ack => type_cast_1972_inst_req_1); -- 
    -- CP-element group 71:  transition  input  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	69 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	72 
    -- CP-element group 71:  members (6) 
      -- CP-element group 71: 	 branch_block_stmt_1825/assign_stmt_2290/WPIPE_Block1_done_2288_sample_completed_
      -- CP-element group 71: 	 branch_block_stmt_1825/assign_stmt_2290/WPIPE_Block1_done_2288_update_start_
      -- CP-element group 71: 	 branch_block_stmt_1825/assign_stmt_2290/WPIPE_Block1_done_2288_Sample/$exit
      -- CP-element group 71: 	 branch_block_stmt_1825/assign_stmt_2290/WPIPE_Block1_done_2288_Sample/ack
      -- CP-element group 71: 	 branch_block_stmt_1825/assign_stmt_2290/WPIPE_Block1_done_2288_Update/$entry
      -- CP-element group 71: 	 branch_block_stmt_1825/assign_stmt_2290/WPIPE_Block1_done_2288_Update/req
      -- 
    ack_6130_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_done_2288_inst_ack_0, ack => convTransposeB_CP_5119_elements(71)); -- 
    req_6134_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6134_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(71), ack => WPIPE_Block1_done_2288_inst_req_1); -- 
    -- CP-element group 72:  transition  place  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	71 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (16) 
      -- CP-element group 72: 	 $exit
      -- CP-element group 72: 	 branch_block_stmt_1825/$exit
      -- CP-element group 72: 	 branch_block_stmt_1825/branch_block_stmt_1825__exit__
      -- CP-element group 72: 	 branch_block_stmt_1825/assign_stmt_2290__exit__
      -- CP-element group 72: 	 branch_block_stmt_1825/return__
      -- CP-element group 72: 	 branch_block_stmt_1825/merge_stmt_2292__exit__
      -- CP-element group 72: 	 branch_block_stmt_1825/assign_stmt_2290/$exit
      -- CP-element group 72: 	 branch_block_stmt_1825/assign_stmt_2290/WPIPE_Block1_done_2288_update_completed_
      -- CP-element group 72: 	 branch_block_stmt_1825/assign_stmt_2290/WPIPE_Block1_done_2288_Update/$exit
      -- CP-element group 72: 	 branch_block_stmt_1825/assign_stmt_2290/WPIPE_Block1_done_2288_Update/ack
      -- CP-element group 72: 	 branch_block_stmt_1825/return___PhiReq/$entry
      -- CP-element group 72: 	 branch_block_stmt_1825/return___PhiReq/$exit
      -- CP-element group 72: 	 branch_block_stmt_1825/merge_stmt_2292_PhiReqMerge
      -- CP-element group 72: 	 branch_block_stmt_1825/merge_stmt_2292_PhiAck/$entry
      -- CP-element group 72: 	 branch_block_stmt_1825/merge_stmt_2292_PhiAck/$exit
      -- CP-element group 72: 	 branch_block_stmt_1825/merge_stmt_2292_PhiAck/dummy
      -- 
    ack_6135_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_done_2288_inst_ack_1, ack => convTransposeB_CP_5119_elements(72)); -- 
    -- CP-element group 73:  transition  output  delay-element  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	31 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	77 
    -- CP-element group 73:  members (4) 
      -- CP-element group 73: 	 branch_block_stmt_1825/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1973/$exit
      -- CP-element group 73: 	 branch_block_stmt_1825/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1973/phi_stmt_1973_sources/$exit
      -- CP-element group 73: 	 branch_block_stmt_1825/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1973/phi_stmt_1973_sources/type_cast_1977_konst_delay_trans
      -- CP-element group 73: 	 branch_block_stmt_1825/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1973/phi_stmt_1973_req
      -- 
    phi_stmt_1973_req_6146_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1973_req_6146_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(73), ack => phi_stmt_1973_req_0); -- 
    -- Element group convTransposeB_CP_5119_elements(73) is a control-delay.
    cp_element_73_delay: control_delay_element  generic map(name => " 73_delay", delay_value => 1)  port map(req => convTransposeB_CP_5119_elements(31), ack => convTransposeB_CP_5119_elements(73), clk => clk, reset =>reset);
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	31 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (2) 
      -- CP-element group 74: 	 branch_block_stmt_1825/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1967/phi_stmt_1967_sources/type_cast_1970/SplitProtocol/Sample/$exit
      -- CP-element group 74: 	 branch_block_stmt_1825/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1967/phi_stmt_1967_sources/type_cast_1970/SplitProtocol/Sample/ra
      -- 
    ra_6163_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1970_inst_ack_0, ack => convTransposeB_CP_5119_elements(74)); -- 
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	31 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	76 
    -- CP-element group 75:  members (2) 
      -- CP-element group 75: 	 branch_block_stmt_1825/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1967/phi_stmt_1967_sources/type_cast_1970/SplitProtocol/Update/$exit
      -- CP-element group 75: 	 branch_block_stmt_1825/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1967/phi_stmt_1967_sources/type_cast_1970/SplitProtocol/Update/ca
      -- 
    ca_6168_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1970_inst_ack_1, ack => convTransposeB_CP_5119_elements(75)); -- 
    -- CP-element group 76:  join  transition  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: 	75 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76:  members (5) 
      -- CP-element group 76: 	 branch_block_stmt_1825/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1967/$exit
      -- CP-element group 76: 	 branch_block_stmt_1825/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1967/phi_stmt_1967_sources/$exit
      -- CP-element group 76: 	 branch_block_stmt_1825/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1967/phi_stmt_1967_sources/type_cast_1970/$exit
      -- CP-element group 76: 	 branch_block_stmt_1825/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1967/phi_stmt_1967_sources/type_cast_1970/SplitProtocol/$exit
      -- CP-element group 76: 	 branch_block_stmt_1825/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1967/phi_stmt_1967_req
      -- 
    phi_stmt_1967_req_6169_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1967_req_6169_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(76), ack => phi_stmt_1967_req_0); -- 
    convTransposeB_cp_element_group_76: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_76"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5119_elements(74) & convTransposeB_CP_5119_elements(75);
      gj_convTransposeB_cp_element_group_76 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5119_elements(76), clk => clk, reset => reset); --
    end block;
    -- CP-element group 77:  join  transition  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	76 
    -- CP-element group 77: 	73 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	85 
    -- CP-element group 77:  members (1) 
      -- CP-element group 77: 	 branch_block_stmt_1825/entry_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5119_elements(76) & convTransposeB_CP_5119_elements(73);
      gj_convTransposeB_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5119_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	70 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	80 
    -- CP-element group 78:  members (2) 
      -- CP-element group 78: 	 branch_block_stmt_1825/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1973/phi_stmt_1973_sources/type_cast_1979/SplitProtocol/Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_1825/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1973/phi_stmt_1973_sources/type_cast_1979/SplitProtocol/Sample/ra
      -- 
    ra_6189_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1979_inst_ack_0, ack => convTransposeB_CP_5119_elements(78)); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	70 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_1825/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1973/phi_stmt_1973_sources/type_cast_1979/SplitProtocol/Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_1825/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1973/phi_stmt_1973_sources/type_cast_1979/SplitProtocol/Update/ca
      -- 
    ca_6194_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1979_inst_ack_1, ack => convTransposeB_CP_5119_elements(79)); -- 
    -- CP-element group 80:  join  transition  output  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	84 
    -- CP-element group 80:  members (5) 
      -- CP-element group 80: 	 branch_block_stmt_1825/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1973/$exit
      -- CP-element group 80: 	 branch_block_stmt_1825/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1973/phi_stmt_1973_sources/$exit
      -- CP-element group 80: 	 branch_block_stmt_1825/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1973/phi_stmt_1973_sources/type_cast_1979/$exit
      -- CP-element group 80: 	 branch_block_stmt_1825/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1973/phi_stmt_1973_sources/type_cast_1979/SplitProtocol/$exit
      -- CP-element group 80: 	 branch_block_stmt_1825/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1973/phi_stmt_1973_req
      -- 
    phi_stmt_1973_req_6195_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1973_req_6195_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(80), ack => phi_stmt_1973_req_1); -- 
    convTransposeB_cp_element_group_80: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_80"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5119_elements(78) & convTransposeB_CP_5119_elements(79);
      gj_convTransposeB_cp_element_group_80 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5119_elements(80), clk => clk, reset => reset); --
    end block;
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	70 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	83 
    -- CP-element group 81:  members (2) 
      -- CP-element group 81: 	 branch_block_stmt_1825/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1967/phi_stmt_1967_sources/type_cast_1972/SplitProtocol/Sample/$exit
      -- CP-element group 81: 	 branch_block_stmt_1825/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1967/phi_stmt_1967_sources/type_cast_1972/SplitProtocol/Sample/ra
      -- 
    ra_6212_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1972_inst_ack_0, ack => convTransposeB_CP_5119_elements(81)); -- 
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	70 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (2) 
      -- CP-element group 82: 	 branch_block_stmt_1825/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1967/phi_stmt_1967_sources/type_cast_1972/SplitProtocol/Update/$exit
      -- CP-element group 82: 	 branch_block_stmt_1825/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1967/phi_stmt_1967_sources/type_cast_1972/SplitProtocol/Update/ca
      -- 
    ca_6217_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1972_inst_ack_1, ack => convTransposeB_CP_5119_elements(82)); -- 
    -- CP-element group 83:  join  transition  output  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	81 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (5) 
      -- CP-element group 83: 	 branch_block_stmt_1825/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1967/$exit
      -- CP-element group 83: 	 branch_block_stmt_1825/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1967/phi_stmt_1967_sources/$exit
      -- CP-element group 83: 	 branch_block_stmt_1825/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1967/phi_stmt_1967_sources/type_cast_1972/$exit
      -- CP-element group 83: 	 branch_block_stmt_1825/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1967/phi_stmt_1967_sources/type_cast_1972/SplitProtocol/$exit
      -- CP-element group 83: 	 branch_block_stmt_1825/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1967/phi_stmt_1967_req
      -- 
    phi_stmt_1967_req_6218_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1967_req_6218_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(83), ack => phi_stmt_1967_req_1); -- 
    convTransposeB_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5119_elements(81) & convTransposeB_CP_5119_elements(82);
      gj_convTransposeB_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5119_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  join  transition  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	80 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84:  members (1) 
      -- CP-element group 84: 	 branch_block_stmt_1825/ifx_xend_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5119_elements(80) & convTransposeB_CP_5119_elements(83);
      gj_convTransposeB_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5119_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  merge  fork  transition  place  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	77 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85: 	86 
    -- CP-element group 85:  members (2) 
      -- CP-element group 85: 	 branch_block_stmt_1825/merge_stmt_1966_PhiReqMerge
      -- CP-element group 85: 	 branch_block_stmt_1825/merge_stmt_1966_PhiAck/$entry
      -- 
    convTransposeB_CP_5119_elements(85) <= OrReduce(convTransposeB_CP_5119_elements(77) & convTransposeB_CP_5119_elements(84));
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	88 
    -- CP-element group 86:  members (1) 
      -- CP-element group 86: 	 branch_block_stmt_1825/merge_stmt_1966_PhiAck/phi_stmt_1967_ack
      -- 
    phi_stmt_1967_ack_6223_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1967_ack_0, ack => convTransposeB_CP_5119_elements(86)); -- 
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (1) 
      -- CP-element group 87: 	 branch_block_stmt_1825/merge_stmt_1966_PhiAck/phi_stmt_1973_ack
      -- 
    phi_stmt_1973_ack_6224_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1973_ack_0, ack => convTransposeB_CP_5119_elements(87)); -- 
    -- CP-element group 88:  join  fork  transition  place  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: 	86 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	33 
    -- CP-element group 88: 	34 
    -- CP-element group 88: 	35 
    -- CP-element group 88: 	32 
    -- CP-element group 88:  members (16) 
      -- CP-element group 88: 	 branch_block_stmt_1825/merge_stmt_1966__exit__
      -- CP-element group 88: 	 branch_block_stmt_1825/assign_stmt_1985_to_assign_stmt_2092__entry__
      -- CP-element group 88: 	 branch_block_stmt_1825/assign_stmt_1985_to_assign_stmt_2092/$entry
      -- CP-element group 88: 	 branch_block_stmt_1825/assign_stmt_1985_to_assign_stmt_2092/type_cast_1984_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_1825/assign_stmt_1985_to_assign_stmt_2092/type_cast_1984_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1825/assign_stmt_1985_to_assign_stmt_2092/type_cast_1984_Sample/$entry
      -- CP-element group 88: 	 branch_block_stmt_1825/assign_stmt_1985_to_assign_stmt_2092/type_cast_1984_Sample/rr
      -- CP-element group 88: 	 branch_block_stmt_1825/assign_stmt_1985_to_assign_stmt_2092/type_cast_1984_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_1825/assign_stmt_1985_to_assign_stmt_2092/type_cast_1984_Update/cr
      -- CP-element group 88: 	 branch_block_stmt_1825/assign_stmt_1985_to_assign_stmt_2092/type_cast_1989_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_1825/assign_stmt_1985_to_assign_stmt_2092/type_cast_1989_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1825/assign_stmt_1985_to_assign_stmt_2092/type_cast_1989_Sample/$entry
      -- CP-element group 88: 	 branch_block_stmt_1825/assign_stmt_1985_to_assign_stmt_2092/type_cast_1989_Sample/rr
      -- CP-element group 88: 	 branch_block_stmt_1825/assign_stmt_1985_to_assign_stmt_2092/type_cast_1989_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_1825/assign_stmt_1985_to_assign_stmt_2092/type_cast_1989_Update/cr
      -- CP-element group 88: 	 branch_block_stmt_1825/merge_stmt_1966_PhiAck/$exit
      -- 
    rr_5736_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5736_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(88), ack => type_cast_1984_inst_req_0); -- 
    cr_5741_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5741_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(88), ack => type_cast_1984_inst_req_1); -- 
    rr_5750_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5750_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(88), ack => type_cast_1989_inst_req_0); -- 
    cr_5755_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5755_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(88), ack => type_cast_1989_inst_req_1); -- 
    convTransposeB_cp_element_group_88: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_88"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5119_elements(87) & convTransposeB_CP_5119_elements(86);
      gj_convTransposeB_cp_element_group_88 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5119_elements(88), clk => clk, reset => reset); --
    end block;
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	59 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (2) 
      -- CP-element group 89: 	 branch_block_stmt_1825/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2095/phi_stmt_2095_sources/type_cast_2101/SplitProtocol/Sample/$exit
      -- CP-element group 89: 	 branch_block_stmt_1825/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2095/phi_stmt_2095_sources/type_cast_2101/SplitProtocol/Sample/ra
      -- 
    ra_6244_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2101_inst_ack_0, ack => convTransposeB_CP_5119_elements(89)); -- 
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	59 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (2) 
      -- CP-element group 90: 	 branch_block_stmt_1825/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2095/phi_stmt_2095_sources/type_cast_2101/SplitProtocol/Update/$exit
      -- CP-element group 90: 	 branch_block_stmt_1825/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2095/phi_stmt_2095_sources/type_cast_2101/SplitProtocol/Update/ca
      -- 
    ca_6249_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2101_inst_ack_1, ack => convTransposeB_CP_5119_elements(90)); -- 
    -- CP-element group 91:  join  transition  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	90 
    -- CP-element group 91: 	89 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	93 
    -- CP-element group 91:  members (6) 
      -- CP-element group 91: 	 branch_block_stmt_1825/ifx_xthen_whilex_xbody_PhiReq/$exit
      -- CP-element group 91: 	 branch_block_stmt_1825/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2095/$exit
      -- CP-element group 91: 	 branch_block_stmt_1825/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2095/phi_stmt_2095_sources/$exit
      -- CP-element group 91: 	 branch_block_stmt_1825/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2095/phi_stmt_2095_sources/type_cast_2101/$exit
      -- CP-element group 91: 	 branch_block_stmt_1825/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2095/phi_stmt_2095_sources/type_cast_2101/SplitProtocol/$exit
      -- CP-element group 91: 	 branch_block_stmt_1825/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2095/phi_stmt_2095_req
      -- 
    phi_stmt_2095_req_6250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2095_req_6250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(91), ack => phi_stmt_2095_req_1); -- 
    convTransposeB_cp_element_group_91: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_91"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5119_elements(90) & convTransposeB_CP_5119_elements(89);
      gj_convTransposeB_cp_element_group_91 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5119_elements(91), clk => clk, reset => reset); --
    end block;
    -- CP-element group 92:  transition  output  delay-element  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	36 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	93 
    -- CP-element group 92:  members (5) 
      -- CP-element group 92: 	 branch_block_stmt_1825/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$exit
      -- CP-element group 92: 	 branch_block_stmt_1825/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2095/$exit
      -- CP-element group 92: 	 branch_block_stmt_1825/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2095/phi_stmt_2095_sources/$exit
      -- CP-element group 92: 	 branch_block_stmt_1825/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2095/phi_stmt_2095_sources/type_cast_2099_konst_delay_trans
      -- CP-element group 92: 	 branch_block_stmt_1825/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2095/phi_stmt_2095_req
      -- 
    phi_stmt_2095_req_6261_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2095_req_6261_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(92), ack => phi_stmt_2095_req_0); -- 
    -- Element group convTransposeB_CP_5119_elements(92) is a control-delay.
    cp_element_92_delay: control_delay_element  generic map(name => " 92_delay", delay_value => 1)  port map(req => convTransposeB_CP_5119_elements(36), ack => convTransposeB_CP_5119_elements(92), clk => clk, reset =>reset);
    -- CP-element group 93:  merge  transition  place  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	91 
    -- CP-element group 93: 	92 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93:  members (2) 
      -- CP-element group 93: 	 branch_block_stmt_1825/merge_stmt_2094_PhiReqMerge
      -- CP-element group 93: 	 branch_block_stmt_1825/merge_stmt_2094_PhiAck/$entry
      -- 
    convTransposeB_CP_5119_elements(93) <= OrReduce(convTransposeB_CP_5119_elements(91) & convTransposeB_CP_5119_elements(92));
    -- CP-element group 94:  fork  transition  place  input  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	37 
    -- CP-element group 94: 	38 
    -- CP-element group 94: 	40 
    -- CP-element group 94: 	55 
    -- CP-element group 94: 	56 
    -- CP-element group 94: 	57 
    -- CP-element group 94: 	42 
    -- CP-element group 94: 	44 
    -- CP-element group 94: 	46 
    -- CP-element group 94: 	48 
    -- CP-element group 94: 	50 
    -- CP-element group 94: 	52 
    -- CP-element group 94:  members (45) 
      -- CP-element group 94: 	 branch_block_stmt_1825/merge_stmt_2094__exit__
      -- CP-element group 94: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200__entry__
      -- CP-element group 94: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/$entry
      -- CP-element group 94: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/type_cast_2111_sample_start_
      -- CP-element group 94: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/type_cast_2111_update_start_
      -- CP-element group 94: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/type_cast_2111_Sample/$entry
      -- CP-element group 94: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/type_cast_2111_Sample/rr
      -- CP-element group 94: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/type_cast_2111_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/type_cast_2111_Update/cr
      -- CP-element group 94: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/type_cast_2141_update_start_
      -- CP-element group 94: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/type_cast_2141_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/type_cast_2141_Update/cr
      -- CP-element group 94: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/addr_of_2148_update_start_
      -- CP-element group 94: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/array_obj_ref_2147_final_index_sum_regn_update_start
      -- CP-element group 94: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/array_obj_ref_2147_final_index_sum_regn_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/array_obj_ref_2147_final_index_sum_regn_Update/req
      -- CP-element group 94: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/addr_of_2148_complete/$entry
      -- CP-element group 94: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/addr_of_2148_complete/req
      -- CP-element group 94: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2152_update_start_
      -- CP-element group 94: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2152_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2152_Update/word_access_complete/$entry
      -- CP-element group 94: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2152_Update/word_access_complete/word_0/$entry
      -- CP-element group 94: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2152_Update/word_access_complete/word_0/cr
      -- CP-element group 94: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/type_cast_2172_update_start_
      -- CP-element group 94: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/type_cast_2172_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/type_cast_2172_Update/cr
      -- CP-element group 94: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/addr_of_2179_update_start_
      -- CP-element group 94: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/array_obj_ref_2178_final_index_sum_regn_update_start
      -- CP-element group 94: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/array_obj_ref_2178_final_index_sum_regn_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/array_obj_ref_2178_final_index_sum_regn_Update/req
      -- CP-element group 94: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/addr_of_2179_complete/$entry
      -- CP-element group 94: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/addr_of_2179_complete/req
      -- CP-element group 94: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2182_update_start_
      -- CP-element group 94: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2182_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2182_Update/word_access_complete/$entry
      -- CP-element group 94: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2182_Update/word_access_complete/word_0/$entry
      -- CP-element group 94: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/ptr_deref_2182_Update/word_access_complete/word_0/cr
      -- CP-element group 94: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/type_cast_2188_sample_start_
      -- CP-element group 94: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/type_cast_2188_update_start_
      -- CP-element group 94: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/type_cast_2188_Sample/$entry
      -- CP-element group 94: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/type_cast_2188_Sample/rr
      -- CP-element group 94: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/type_cast_2188_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_1825/assign_stmt_2108_to_assign_stmt_2200/type_cast_2188_Update/cr
      -- CP-element group 94: 	 branch_block_stmt_1825/merge_stmt_2094_PhiAck/$exit
      -- CP-element group 94: 	 branch_block_stmt_1825/merge_stmt_2094_PhiAck/phi_stmt_2095_ack
      -- 
    phi_stmt_2095_ack_6266_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2095_ack_0, ack => convTransposeB_CP_5119_elements(94)); -- 
    rr_5767_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5767_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(94), ack => type_cast_2111_inst_req_0); -- 
    cr_5772_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5772_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(94), ack => type_cast_2111_inst_req_1); -- 
    cr_5786_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5786_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(94), ack => type_cast_2141_inst_req_1); -- 
    req_5817_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5817_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(94), ack => array_obj_ref_2147_index_offset_req_1); -- 
    req_5832_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5832_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(94), ack => addr_of_2148_final_reg_req_1); -- 
    cr_5877_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5877_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(94), ack => ptr_deref_2152_load_0_req_1); -- 
    cr_5896_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5896_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(94), ack => type_cast_2172_inst_req_1); -- 
    req_5927_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5927_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(94), ack => array_obj_ref_2178_index_offset_req_1); -- 
    req_5942_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5942_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(94), ack => addr_of_2179_final_reg_req_1); -- 
    cr_5992_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5992_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(94), ack => ptr_deref_2182_store_0_req_1); -- 
    rr_6001_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6001_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(94), ack => type_cast_2188_inst_req_0); -- 
    cr_6006_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6006_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(94), ack => type_cast_2188_inst_req_1); -- 
    -- CP-element group 95:  transition  input  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	64 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	97 
    -- CP-element group 95:  members (2) 
      -- CP-element group 95: 	 branch_block_stmt_1825/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2257/phi_stmt_2257_sources/type_cast_2262/SplitProtocol/Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_1825/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2257/phi_stmt_2257_sources/type_cast_2262/SplitProtocol/Sample/ra
      -- 
    ra_6318_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2262_inst_ack_0, ack => convTransposeB_CP_5119_elements(95)); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	64 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (2) 
      -- CP-element group 96: 	 branch_block_stmt_1825/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2257/phi_stmt_2257_sources/type_cast_2262/SplitProtocol/Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_1825/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2257/phi_stmt_2257_sources/type_cast_2262/SplitProtocol/Update/ca
      -- 
    ca_6323_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2262_inst_ack_1, ack => convTransposeB_CP_5119_elements(96)); -- 
    -- CP-element group 97:  join  transition  output  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	96 
    -- CP-element group 97: 	95 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	101 
    -- CP-element group 97:  members (5) 
      -- CP-element group 97: 	 branch_block_stmt_1825/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2257/$exit
      -- CP-element group 97: 	 branch_block_stmt_1825/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2257/phi_stmt_2257_sources/$exit
      -- CP-element group 97: 	 branch_block_stmt_1825/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2257/phi_stmt_2257_sources/type_cast_2262/$exit
      -- CP-element group 97: 	 branch_block_stmt_1825/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2257/phi_stmt_2257_sources/type_cast_2262/SplitProtocol/$exit
      -- CP-element group 97: 	 branch_block_stmt_1825/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2257/phi_stmt_2257_req
      -- 
    phi_stmt_2257_req_6324_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2257_req_6324_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(97), ack => phi_stmt_2257_req_1); -- 
    convTransposeB_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5119_elements(96) & convTransposeB_CP_5119_elements(95);
      gj_convTransposeB_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5119_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	64 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	100 
    -- CP-element group 98:  members (2) 
      -- CP-element group 98: 	 branch_block_stmt_1825/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2263/phi_stmt_2263_sources/type_cast_2268/SplitProtocol/Sample/$exit
      -- CP-element group 98: 	 branch_block_stmt_1825/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2263/phi_stmt_2263_sources/type_cast_2268/SplitProtocol/Sample/ra
      -- 
    ra_6341_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2268_inst_ack_0, ack => convTransposeB_CP_5119_elements(98)); -- 
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	64 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99:  members (2) 
      -- CP-element group 99: 	 branch_block_stmt_1825/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2263/phi_stmt_2263_sources/type_cast_2268/SplitProtocol/Update/$exit
      -- CP-element group 99: 	 branch_block_stmt_1825/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2263/phi_stmt_2263_sources/type_cast_2268/SplitProtocol/Update/ca
      -- 
    ca_6346_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2268_inst_ack_1, ack => convTransposeB_CP_5119_elements(99)); -- 
    -- CP-element group 100:  join  transition  output  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	98 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	101 
    -- CP-element group 100:  members (5) 
      -- CP-element group 100: 	 branch_block_stmt_1825/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2263/$exit
      -- CP-element group 100: 	 branch_block_stmt_1825/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2263/phi_stmt_2263_sources/$exit
      -- CP-element group 100: 	 branch_block_stmt_1825/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2263/phi_stmt_2263_sources/type_cast_2268/$exit
      -- CP-element group 100: 	 branch_block_stmt_1825/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2263/phi_stmt_2263_sources/type_cast_2268/SplitProtocol/$exit
      -- CP-element group 100: 	 branch_block_stmt_1825/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2263/phi_stmt_2263_req
      -- 
    phi_stmt_2263_req_6347_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2263_req_6347_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(100), ack => phi_stmt_2263_req_1); -- 
    convTransposeB_cp_element_group_100: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_100"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5119_elements(98) & convTransposeB_CP_5119_elements(99);
      gj_convTransposeB_cp_element_group_100 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5119_elements(100), clk => clk, reset => reset); --
    end block;
    -- CP-element group 101:  join  transition  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	97 
    -- CP-element group 101: 	100 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	109 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_1825/ifx_xelse_ifx_xend_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_101: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_101"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5119_elements(97) & convTransposeB_CP_5119_elements(100);
      gj_convTransposeB_cp_element_group_101 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5119_elements(101), clk => clk, reset => reset); --
    end block;
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	66 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	104 
    -- CP-element group 102:  members (2) 
      -- CP-element group 102: 	 branch_block_stmt_1825/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2257/phi_stmt_2257_sources/type_cast_2260/SplitProtocol/Sample/$exit
      -- CP-element group 102: 	 branch_block_stmt_1825/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2257/phi_stmt_2257_sources/type_cast_2260/SplitProtocol/Sample/ra
      -- 
    ra_6367_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2260_inst_ack_0, ack => convTransposeB_CP_5119_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	66 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (2) 
      -- CP-element group 103: 	 branch_block_stmt_1825/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2257/phi_stmt_2257_sources/type_cast_2260/SplitProtocol/Update/$exit
      -- CP-element group 103: 	 branch_block_stmt_1825/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2257/phi_stmt_2257_sources/type_cast_2260/SplitProtocol/Update/ca
      -- 
    ca_6372_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2260_inst_ack_1, ack => convTransposeB_CP_5119_elements(103)); -- 
    -- CP-element group 104:  join  transition  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	102 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	108 
    -- CP-element group 104:  members (5) 
      -- CP-element group 104: 	 branch_block_stmt_1825/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2257/$exit
      -- CP-element group 104: 	 branch_block_stmt_1825/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2257/phi_stmt_2257_sources/$exit
      -- CP-element group 104: 	 branch_block_stmt_1825/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2257/phi_stmt_2257_sources/type_cast_2260/$exit
      -- CP-element group 104: 	 branch_block_stmt_1825/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2257/phi_stmt_2257_sources/type_cast_2260/SplitProtocol/$exit
      -- CP-element group 104: 	 branch_block_stmt_1825/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2257/phi_stmt_2257_req
      -- 
    phi_stmt_2257_req_6373_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2257_req_6373_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(104), ack => phi_stmt_2257_req_0); -- 
    convTransposeB_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5119_elements(102) & convTransposeB_CP_5119_elements(103);
      gj_convTransposeB_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5119_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	66 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	107 
    -- CP-element group 105:  members (2) 
      -- CP-element group 105: 	 branch_block_stmt_1825/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2263/phi_stmt_2263_sources/type_cast_2266/SplitProtocol/Sample/$exit
      -- CP-element group 105: 	 branch_block_stmt_1825/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2263/phi_stmt_2263_sources/type_cast_2266/SplitProtocol/Sample/ra
      -- 
    ra_6390_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2266_inst_ack_0, ack => convTransposeB_CP_5119_elements(105)); -- 
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	66 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_1825/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2263/phi_stmt_2263_sources/type_cast_2266/SplitProtocol/Update/$exit
      -- CP-element group 106: 	 branch_block_stmt_1825/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2263/phi_stmt_2263_sources/type_cast_2266/SplitProtocol/Update/ca
      -- 
    ca_6395_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2266_inst_ack_1, ack => convTransposeB_CP_5119_elements(106)); -- 
    -- CP-element group 107:  join  transition  output  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	105 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107:  members (5) 
      -- CP-element group 107: 	 branch_block_stmt_1825/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2263/$exit
      -- CP-element group 107: 	 branch_block_stmt_1825/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2263/phi_stmt_2263_sources/$exit
      -- CP-element group 107: 	 branch_block_stmt_1825/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2263/phi_stmt_2263_sources/type_cast_2266/$exit
      -- CP-element group 107: 	 branch_block_stmt_1825/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2263/phi_stmt_2263_sources/type_cast_2266/SplitProtocol/$exit
      -- CP-element group 107: 	 branch_block_stmt_1825/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2263/phi_stmt_2263_req
      -- 
    phi_stmt_2263_req_6396_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2263_req_6396_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(107), ack => phi_stmt_2263_req_0); -- 
    convTransposeB_cp_element_group_107: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_107"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5119_elements(105) & convTransposeB_CP_5119_elements(106);
      gj_convTransposeB_cp_element_group_107 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5119_elements(107), clk => clk, reset => reset); --
    end block;
    -- CP-element group 108:  join  transition  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	107 
    -- CP-element group 108: 	104 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	109 
    -- CP-element group 108:  members (1) 
      -- CP-element group 108: 	 branch_block_stmt_1825/ifx_xthen79_ifx_xend_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5119_elements(107) & convTransposeB_CP_5119_elements(104);
      gj_convTransposeB_cp_element_group_108 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5119_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  merge  fork  transition  place  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	101 
    -- CP-element group 109: 	108 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	110 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (2) 
      -- CP-element group 109: 	 branch_block_stmt_1825/merge_stmt_2256_PhiReqMerge
      -- CP-element group 109: 	 branch_block_stmt_1825/merge_stmt_2256_PhiAck/$entry
      -- 
    convTransposeB_CP_5119_elements(109) <= OrReduce(convTransposeB_CP_5119_elements(101) & convTransposeB_CP_5119_elements(108));
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	109 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	112 
    -- CP-element group 110:  members (1) 
      -- CP-element group 110: 	 branch_block_stmt_1825/merge_stmt_2256_PhiAck/phi_stmt_2257_ack
      -- 
    phi_stmt_2257_ack_6401_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2257_ack_0, ack => convTransposeB_CP_5119_elements(110)); -- 
    -- CP-element group 111:  transition  input  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111:  members (1) 
      -- CP-element group 111: 	 branch_block_stmt_1825/merge_stmt_2256_PhiAck/phi_stmt_2263_ack
      -- 
    phi_stmt_2263_ack_6402_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2263_ack_0, ack => convTransposeB_CP_5119_elements(111)); -- 
    -- CP-element group 112:  join  fork  transition  place  output  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	110 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	67 
    -- CP-element group 112: 	68 
    -- CP-element group 112:  members (10) 
      -- CP-element group 112: 	 branch_block_stmt_1825/merge_stmt_2256__exit__
      -- CP-element group 112: 	 branch_block_stmt_1825/assign_stmt_2274_to_assign_stmt_2279__entry__
      -- CP-element group 112: 	 branch_block_stmt_1825/assign_stmt_2274_to_assign_stmt_2279/$entry
      -- CP-element group 112: 	 branch_block_stmt_1825/assign_stmt_2274_to_assign_stmt_2279/type_cast_2273_sample_start_
      -- CP-element group 112: 	 branch_block_stmt_1825/assign_stmt_2274_to_assign_stmt_2279/type_cast_2273_update_start_
      -- CP-element group 112: 	 branch_block_stmt_1825/assign_stmt_2274_to_assign_stmt_2279/type_cast_2273_Sample/$entry
      -- CP-element group 112: 	 branch_block_stmt_1825/assign_stmt_2274_to_assign_stmt_2279/type_cast_2273_Sample/rr
      -- CP-element group 112: 	 branch_block_stmt_1825/assign_stmt_2274_to_assign_stmt_2279/type_cast_2273_Update/$entry
      -- CP-element group 112: 	 branch_block_stmt_1825/assign_stmt_2274_to_assign_stmt_2279/type_cast_2273_Update/cr
      -- CP-element group 112: 	 branch_block_stmt_1825/merge_stmt_2256_PhiAck/$exit
      -- 
    rr_6093_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6093_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(112), ack => type_cast_2273_inst_req_0); -- 
    cr_6098_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6098_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5119_elements(112), ack => type_cast_2273_inst_req_1); -- 
    convTransposeB_cp_element_group_112: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_112"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5119_elements(110) & convTransposeB_CP_5119_elements(111);
      gj_convTransposeB_cp_element_group_112 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5119_elements(112), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i32_i32_2054_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2075_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2135_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2166_wire : std_logic_vector(31 downto 0);
    signal LOAD_padding_1891_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_padding_1891_word_address_0 : std_logic_vector(0 downto 0);
    signal R_idxprom61_2177_resized : std_logic_vector(13 downto 0);
    signal R_idxprom61_2177_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_2146_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_2146_scaled : std_logic_vector(13 downto 0);
    signal add17_2117 : std_logic_vector(31 downto 0);
    signal add25_2015 : std_logic_vector(31 downto 0);
    signal add36_2030 : std_logic_vector(31 downto 0);
    signal add51_2087 : std_logic_vector(31 downto 0);
    signal add53_2122 : std_logic_vector(31 downto 0);
    signal add66_2195 : std_logic_vector(31 downto 0);
    signal add_2000 : std_logic_vector(31 downto 0);
    signal array_obj_ref_2147_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2147_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2147_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2147_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2147_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2147_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2178_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2178_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2178_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2178_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2178_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2178_root_address : std_logic_vector(13 downto 0);
    signal arrayidx62_2180 : std_logic_vector(31 downto 0);
    signal arrayidx_2149 : std_logic_vector(31 downto 0);
    signal call_1828 : std_logic_vector(15 downto 0);
    signal cmp77_2231 : std_logic_vector(0 downto 0);
    signal cmp89_2279 : std_logic_vector(0 downto 0);
    signal cmp_2200 : std_logic_vector(0 downto 0);
    signal conv12_1985 : std_logic_vector(31 downto 0);
    signal conv15_1990 : std_logic_vector(31 downto 0);
    signal conv22_1877 : std_logic_vector(31 downto 0);
    signal conv27_1896 : std_logic_vector(31 downto 0);
    signal conv33_1910 : std_logic_vector(31 downto 0);
    signal conv46_2056 : std_logic_vector(31 downto 0);
    signal conv49_2077 : std_logic_vector(31 downto 0);
    signal conv65_2189 : std_logic_vector(31 downto 0);
    signal conv75_2226 : std_logic_vector(31 downto 0);
    signal conv84_2254 : std_logic_vector(15 downto 0);
    signal conv86_2274 : std_logic_vector(31 downto 0);
    signal conv9102_2112 : std_logic_vector(31 downto 0);
    signal conv_1851 : std_logic_vector(15 downto 0);
    signal div83_2250 : std_logic_vector(31 downto 0);
    signal div88_1964 : std_logic_vector(31 downto 0);
    signal div_1847 : std_logic_vector(31 downto 0);
    signal iNsTr_10_1954 : std_logic_vector(31 downto 0);
    signal iNsTr_2_1837 : std_logic_vector(31 downto 0);
    signal iNsTr_3_1859 : std_logic_vector(31 downto 0);
    signal iNsTr_4_1869 : std_logic_vector(31 downto 0);
    signal iNsTr_5_1885 : std_logic_vector(31 downto 0);
    signal iNsTr_6_1902 : std_logic_vector(31 downto 0);
    signal iNsTr_7_1918 : std_logic_vector(31 downto 0);
    signal iNsTr_8_1930 : std_logic_vector(31 downto 0);
    signal iNsTr_9_1942 : std_logic_vector(31 downto 0);
    signal idxprom61_2173 : std_logic_vector(63 downto 0);
    signal idxprom_2142 : std_logic_vector(63 downto 0);
    signal inc81_2244 : std_logic_vector(15 downto 0);
    signal inc_2221 : std_logic_vector(15 downto 0);
    signal indvar_2095 : std_logic_vector(15 downto 0);
    signal indvarx_xnext_2213 : std_logic_vector(15 downto 0);
    signal input_dim0x_x0_2263 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2x_xph_1973 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1x_xph_1967 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_2257 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_2108 : std_logic_vector(15 downto 0);
    signal mul16_2005 : std_logic_vector(31 downto 0);
    signal mul23_2010 : std_logic_vector(31 downto 0);
    signal mul34_2025 : std_logic_vector(31 downto 0);
    signal mul50_2082 : std_logic_vector(31 downto 0);
    signal mul52_2092 : std_logic_vector(31 downto 0);
    signal mul_1995 : std_logic_vector(31 downto 0);
    signal ptr_deref_1840_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1840_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1840_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1840_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1840_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1862_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1862_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1862_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1862_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1862_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1872_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1872_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1872_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1872_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1872_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1888_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1888_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1888_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1888_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1888_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1905_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1905_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1905_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1905_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1905_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1921_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1921_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1921_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1921_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1921_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1933_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1933_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1933_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1933_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1933_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1945_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1945_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1945_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1945_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1945_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1957_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1957_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1957_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1957_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1957_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2152_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2152_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2152_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2152_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2152_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2182_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2182_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2182_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2182_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2182_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2182_word_offset_0 : std_logic_vector(13 downto 0);
    signal sext103_2068 : std_logic_vector(31 downto 0);
    signal sext105_2128 : std_logic_vector(31 downto 0);
    signal sext106_2159 : std_logic_vector(31 downto 0);
    signal sext_2047 : std_logic_vector(31 downto 0);
    signal shr60_2168 : std_logic_vector(31 downto 0);
    signal shr_2137 : std_logic_vector(31 downto 0);
    signal sub28_2062 : std_logic_vector(31 downto 0);
    signal sub39_2035 : std_logic_vector(31 downto 0);
    signal sub40_2041 : std_logic_vector(31 downto 0);
    signal sub_2020 : std_logic_vector(31 downto 0);
    signal tmp10_1863 : std_logic_vector(31 downto 0);
    signal tmp21_1873 : std_logic_vector(7 downto 0);
    signal tmp24_1889 : std_logic_vector(31 downto 0);
    signal tmp26_1892 : std_logic_vector(7 downto 0);
    signal tmp32_1906 : std_logic_vector(7 downto 0);
    signal tmp35_1922 : std_logic_vector(31 downto 0);
    signal tmp44_1934 : std_logic_vector(31 downto 0);
    signal tmp47_1946 : std_logic_vector(31 downto 0);
    signal tmp57_2153 : std_logic_vector(63 downto 0);
    signal tmp87_1958 : std_logic_vector(31 downto 0);
    signal tmp_1841 : std_logic_vector(31 downto 0);
    signal type_cast_1845_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1962_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1970_wire : std_logic_vector(15 downto 0);
    signal type_cast_1972_wire : std_logic_vector(15 downto 0);
    signal type_cast_1977_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1979_wire : std_logic_vector(15 downto 0);
    signal type_cast_1983_wire : std_logic_vector(31 downto 0);
    signal type_cast_1988_wire : std_logic_vector(31 downto 0);
    signal type_cast_2039_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2045_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2050_wire : std_logic_vector(31 downto 0);
    signal type_cast_2053_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2060_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2066_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2071_wire : std_logic_vector(31 downto 0);
    signal type_cast_2074_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2099_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2101_wire : std_logic_vector(15 downto 0);
    signal type_cast_2106_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2126_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2131_wire : std_logic_vector(31 downto 0);
    signal type_cast_2134_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2140_wire : std_logic_vector(63 downto 0);
    signal type_cast_2157_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2162_wire : std_logic_vector(31 downto 0);
    signal type_cast_2165_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2171_wire : std_logic_vector(63 downto 0);
    signal type_cast_2187_wire : std_logic_vector(31 downto 0);
    signal type_cast_2193_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2211_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2219_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2224_wire : std_logic_vector(31 downto 0);
    signal type_cast_2242_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2248_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2260_wire : std_logic_vector(15 downto 0);
    signal type_cast_2262_wire : std_logic_vector(15 downto 0);
    signal type_cast_2266_wire : std_logic_vector(15 downto 0);
    signal type_cast_2268_wire : std_logic_vector(15 downto 0);
    signal type_cast_2272_wire : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    LOAD_padding_1891_word_address_0 <= "0";
    array_obj_ref_2147_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2147_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2147_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2147_resized_base_address <= "00000000000000";
    array_obj_ref_2178_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2178_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2178_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2178_resized_base_address <= "00000000000000";
    iNsTr_10_1954 <= "00000000000000000000000000000011";
    iNsTr_2_1837 <= "00000000000000000000000000000100";
    iNsTr_3_1859 <= "00000000000000000000000000000101";
    iNsTr_4_1869 <= "00000000000000000000000000000000";
    iNsTr_5_1885 <= "00000000000000000000000000000100";
    iNsTr_6_1902 <= "00000000000000000000000000000001";
    iNsTr_7_1918 <= "00000000000000000000000000000101";
    iNsTr_8_1930 <= "00000000000000000000000000000101";
    iNsTr_9_1942 <= "00000000000000000000000000000100";
    ptr_deref_1840_word_offset_0 <= "0000000";
    ptr_deref_1862_word_offset_0 <= "0000000";
    ptr_deref_1872_word_offset_0 <= "0";
    ptr_deref_1888_word_offset_0 <= "0000000";
    ptr_deref_1905_word_offset_0 <= "0";
    ptr_deref_1921_word_offset_0 <= "0000000";
    ptr_deref_1933_word_offset_0 <= "0000000";
    ptr_deref_1945_word_offset_0 <= "0000000";
    ptr_deref_1957_word_offset_0 <= "0000000";
    ptr_deref_2152_word_offset_0 <= "00000000000000";
    ptr_deref_2182_word_offset_0 <= "00000000000000";
    type_cast_1845_wire_constant <= "00000000000000000000000000000001";
    type_cast_1962_wire_constant <= "00000000000000000000000000000001";
    type_cast_1977_wire_constant <= "0000000000000000";
    type_cast_2039_wire_constant <= "00000000000000000000000000010000";
    type_cast_2045_wire_constant <= "11111111111111110000000000000000";
    type_cast_2053_wire_constant <= "00000000000000000000000000010000";
    type_cast_2060_wire_constant <= "00000000000000000000000000010000";
    type_cast_2066_wire_constant <= "11111111111111110000000000000000";
    type_cast_2074_wire_constant <= "00000000000000000000000000010000";
    type_cast_2099_wire_constant <= "0000000000000000";
    type_cast_2106_wire_constant <= "0000000000000100";
    type_cast_2126_wire_constant <= "00000000000000000000000000010000";
    type_cast_2134_wire_constant <= "00000000000000000000000000010010";
    type_cast_2157_wire_constant <= "00000000000000000000000000010000";
    type_cast_2165_wire_constant <= "00000000000000000000000000010010";
    type_cast_2193_wire_constant <= "00000000000000000000000000000100";
    type_cast_2211_wire_constant <= "0000000000000001";
    type_cast_2219_wire_constant <= "0000000000000001";
    type_cast_2242_wire_constant <= "0000000000000001";
    type_cast_2248_wire_constant <= "00000000000000000000000000000001";
    phi_stmt_1967: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1970_wire & type_cast_1972_wire;
      req <= phi_stmt_1967_req_0 & phi_stmt_1967_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1967",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1967_ack_0,
          idata => idata,
          odata => input_dim1x_x1x_xph_1967,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1967
    phi_stmt_1973: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1977_wire_constant & type_cast_1979_wire;
      req <= phi_stmt_1973_req_0 & phi_stmt_1973_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1973",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1973_ack_0,
          idata => idata,
          odata => input_dim0x_x2x_xph_1973,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1973
    phi_stmt_2095: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2099_wire_constant & type_cast_2101_wire;
      req <= phi_stmt_2095_req_0 & phi_stmt_2095_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2095",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2095_ack_0,
          idata => idata,
          odata => indvar_2095,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2095
    phi_stmt_2257: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2260_wire & type_cast_2262_wire;
      req <= phi_stmt_2257_req_0 & phi_stmt_2257_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2257",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2257_ack_0,
          idata => idata,
          odata => input_dim1x_x2_2257,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2257
    phi_stmt_2263: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2266_wire & type_cast_2268_wire;
      req <= phi_stmt_2263_req_0 & phi_stmt_2263_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2263",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2263_ack_0,
          idata => idata,
          odata => input_dim0x_x0_2263,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2263
    addr_of_2148_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2148_final_reg_req_0;
      addr_of_2148_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2148_final_reg_req_1;
      addr_of_2148_final_reg_ack_1<= rack(0);
      addr_of_2148_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2148_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2147_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_2149,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2179_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2179_final_reg_req_0;
      addr_of_2179_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2179_final_reg_req_1;
      addr_of_2179_final_reg_ack_1<= rack(0);
      addr_of_2179_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2179_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2178_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx62_2180,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1850_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1850_inst_req_0;
      type_cast_1850_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1850_inst_req_1;
      type_cast_1850_inst_ack_1<= rack(0);
      type_cast_1850_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1850_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div_1847,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_1851,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1876_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1876_inst_req_0;
      type_cast_1876_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1876_inst_req_1;
      type_cast_1876_inst_ack_1<= rack(0);
      type_cast_1876_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1876_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp21_1873,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv22_1877,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1895_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1895_inst_req_0;
      type_cast_1895_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1895_inst_req_1;
      type_cast_1895_inst_ack_1<= rack(0);
      type_cast_1895_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1895_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp26_1892,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv27_1896,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1909_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1909_inst_req_0;
      type_cast_1909_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1909_inst_req_1;
      type_cast_1909_inst_ack_1<= rack(0);
      type_cast_1909_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1909_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp32_1906,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv33_1910,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1970_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1970_inst_req_0;
      type_cast_1970_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1970_inst_req_1;
      type_cast_1970_inst_ack_1<= rack(0);
      type_cast_1970_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1970_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv_1851,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1970_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1972_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1972_inst_req_0;
      type_cast_1972_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1972_inst_req_1;
      type_cast_1972_inst_ack_1<= rack(0);
      type_cast_1972_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1972_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_2257,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1972_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1979_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1979_inst_req_0;
      type_cast_1979_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1979_inst_req_1;
      type_cast_1979_inst_ack_1<= rack(0);
      type_cast_1979_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1979_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x0_2263,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1979_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1984_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1984_inst_req_0;
      type_cast_1984_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1984_inst_req_1;
      type_cast_1984_inst_ack_1<= rack(0);
      type_cast_1984_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1984_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1983_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv12_1985,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1989_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1989_inst_req_0;
      type_cast_1989_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1989_inst_req_1;
      type_cast_1989_inst_ack_1<= rack(0);
      type_cast_1989_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1989_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1988_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv15_1990,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2050_inst
    process(sext_2047) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext_2047(31 downto 0);
      type_cast_2050_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2055_inst
    process(ASHR_i32_i32_2054_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2054_wire(31 downto 0);
      conv46_2056 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2071_inst
    process(sext103_2068) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext103_2068(31 downto 0);
      type_cast_2071_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2076_inst
    process(ASHR_i32_i32_2075_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2075_wire(31 downto 0);
      conv49_2077 <= tmp_var; -- 
    end process;
    type_cast_2101_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2101_inst_req_0;
      type_cast_2101_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2101_inst_req_1;
      type_cast_2101_inst_ack_1<= rack(0);
      type_cast_2101_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2101_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_2213,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2101_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2111_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2111_inst_req_0;
      type_cast_2111_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2111_inst_req_1;
      type_cast_2111_inst_ack_1<= rack(0);
      type_cast_2111_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2111_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_2108,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv9102_2112,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2131_inst
    process(sext105_2128) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext105_2128(31 downto 0);
      type_cast_2131_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2136_inst
    process(ASHR_i32_i32_2135_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2135_wire(31 downto 0);
      shr_2137 <= tmp_var; -- 
    end process;
    type_cast_2141_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2141_inst_req_0;
      type_cast_2141_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2141_inst_req_1;
      type_cast_2141_inst_ack_1<= rack(0);
      type_cast_2141_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2141_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2140_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_2142,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2162_inst
    process(sext106_2159) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext106_2159(31 downto 0);
      type_cast_2162_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2167_inst
    process(ASHR_i32_i32_2166_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2166_wire(31 downto 0);
      shr60_2168 <= tmp_var; -- 
    end process;
    type_cast_2172_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2172_inst_req_0;
      type_cast_2172_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2172_inst_req_1;
      type_cast_2172_inst_ack_1<= rack(0);
      type_cast_2172_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2172_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2171_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom61_2173,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2188_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2188_inst_req_0;
      type_cast_2188_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2188_inst_req_1;
      type_cast_2188_inst_ack_1<= rack(0);
      type_cast_2188_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2188_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2187_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv65_2189,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2225_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2225_inst_req_0;
      type_cast_2225_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2225_inst_req_1;
      type_cast_2225_inst_ack_1<= rack(0);
      type_cast_2225_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2225_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2224_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv75_2226,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2253_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2253_inst_req_0;
      type_cast_2253_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2253_inst_req_1;
      type_cast_2253_inst_ack_1<= rack(0);
      type_cast_2253_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2253_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div83_2250,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv84_2254,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2260_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2260_inst_req_0;
      type_cast_2260_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2260_inst_req_1;
      type_cast_2260_inst_ack_1<= rack(0);
      type_cast_2260_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2260_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv84_2254,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2260_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2262_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2262_inst_req_0;
      type_cast_2262_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2262_inst_req_1;
      type_cast_2262_inst_ack_1<= rack(0);
      type_cast_2262_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2262_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc_2221,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2262_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2266_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2266_inst_req_0;
      type_cast_2266_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2266_inst_req_1;
      type_cast_2266_inst_ack_1<= rack(0);
      type_cast_2266_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2266_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc81_2244,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2266_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2268_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2268_inst_req_0;
      type_cast_2268_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2268_inst_req_1;
      type_cast_2268_inst_ack_1<= rack(0);
      type_cast_2268_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2268_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x2x_xph_1973,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2268_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2273_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2273_inst_req_0;
      type_cast_2273_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2273_inst_req_1;
      type_cast_2273_inst_ack_1<= rack(0);
      type_cast_2273_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2273_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2272_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv86_2274,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence LOAD_padding_1891_gather_scatter
    process(LOAD_padding_1891_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_padding_1891_data_0;
      ov(7 downto 0) := iv;
      tmp26_1892 <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2147_index_1_rename
    process(R_idxprom_2146_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_2146_resized;
      ov(13 downto 0) := iv;
      R_idxprom_2146_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2147_index_1_resize
    process(idxprom_2142) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_2142;
      ov := iv(13 downto 0);
      R_idxprom_2146_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2147_root_address_inst
    process(array_obj_ref_2147_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2147_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2147_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2178_index_1_rename
    process(R_idxprom61_2177_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom61_2177_resized;
      ov(13 downto 0) := iv;
      R_idxprom61_2177_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2178_index_1_resize
    process(idxprom61_2173) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom61_2173;
      ov := iv(13 downto 0);
      R_idxprom61_2177_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2178_root_address_inst
    process(array_obj_ref_2178_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2178_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2178_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1840_addr_0
    process(ptr_deref_1840_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1840_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1840_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1840_base_resize
    process(iNsTr_2_1837) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_2_1837;
      ov := iv(6 downto 0);
      ptr_deref_1840_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1840_gather_scatter
    process(ptr_deref_1840_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1840_data_0;
      ov(31 downto 0) := iv;
      tmp_1841 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1840_root_address_inst
    process(ptr_deref_1840_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1840_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1840_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1862_addr_0
    process(ptr_deref_1862_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1862_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1862_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1862_base_resize
    process(iNsTr_3_1859) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_3_1859;
      ov := iv(6 downto 0);
      ptr_deref_1862_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1862_gather_scatter
    process(ptr_deref_1862_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1862_data_0;
      ov(31 downto 0) := iv;
      tmp10_1863 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1862_root_address_inst
    process(ptr_deref_1862_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1862_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1862_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1872_addr_0
    process(ptr_deref_1872_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1872_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_1872_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1872_base_resize
    process(iNsTr_4_1869) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_4_1869;
      ov := iv(0 downto 0);
      ptr_deref_1872_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1872_gather_scatter
    process(ptr_deref_1872_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1872_data_0;
      ov(7 downto 0) := iv;
      tmp21_1873 <= ov(7 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1872_root_address_inst
    process(ptr_deref_1872_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1872_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_1872_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1888_addr_0
    process(ptr_deref_1888_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1888_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1888_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1888_base_resize
    process(iNsTr_5_1885) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_5_1885;
      ov := iv(6 downto 0);
      ptr_deref_1888_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1888_gather_scatter
    process(ptr_deref_1888_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1888_data_0;
      ov(31 downto 0) := iv;
      tmp24_1889 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1888_root_address_inst
    process(ptr_deref_1888_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1888_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1888_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1905_addr_0
    process(ptr_deref_1905_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1905_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_1905_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1905_base_resize
    process(iNsTr_6_1902) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_6_1902;
      ov := iv(0 downto 0);
      ptr_deref_1905_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1905_gather_scatter
    process(ptr_deref_1905_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1905_data_0;
      ov(7 downto 0) := iv;
      tmp32_1906 <= ov(7 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1905_root_address_inst
    process(ptr_deref_1905_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1905_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_1905_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1921_addr_0
    process(ptr_deref_1921_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1921_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1921_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1921_base_resize
    process(iNsTr_7_1918) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_7_1918;
      ov := iv(6 downto 0);
      ptr_deref_1921_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1921_gather_scatter
    process(ptr_deref_1921_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1921_data_0;
      ov(31 downto 0) := iv;
      tmp35_1922 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1921_root_address_inst
    process(ptr_deref_1921_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1921_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1921_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1933_addr_0
    process(ptr_deref_1933_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1933_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1933_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1933_base_resize
    process(iNsTr_8_1930) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_8_1930;
      ov := iv(6 downto 0);
      ptr_deref_1933_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1933_gather_scatter
    process(ptr_deref_1933_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1933_data_0;
      ov(31 downto 0) := iv;
      tmp44_1934 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1933_root_address_inst
    process(ptr_deref_1933_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1933_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1933_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1945_addr_0
    process(ptr_deref_1945_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1945_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1945_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1945_base_resize
    process(iNsTr_9_1942) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_9_1942;
      ov := iv(6 downto 0);
      ptr_deref_1945_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1945_gather_scatter
    process(ptr_deref_1945_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1945_data_0;
      ov(31 downto 0) := iv;
      tmp47_1946 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1945_root_address_inst
    process(ptr_deref_1945_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1945_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1945_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1957_addr_0
    process(ptr_deref_1957_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1957_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1957_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1957_base_resize
    process(iNsTr_10_1954) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_10_1954;
      ov := iv(6 downto 0);
      ptr_deref_1957_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1957_gather_scatter
    process(ptr_deref_1957_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1957_data_0;
      ov(31 downto 0) := iv;
      tmp87_1958 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1957_root_address_inst
    process(ptr_deref_1957_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1957_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1957_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2152_addr_0
    process(ptr_deref_2152_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2152_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2152_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2152_base_resize
    process(arrayidx_2149) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_2149;
      ov := iv(13 downto 0);
      ptr_deref_2152_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2152_gather_scatter
    process(ptr_deref_2152_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2152_data_0;
      ov(63 downto 0) := iv;
      tmp57_2153 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2152_root_address_inst
    process(ptr_deref_2152_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2152_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2152_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2182_addr_0
    process(ptr_deref_2182_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2182_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2182_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2182_base_resize
    process(arrayidx62_2180) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx62_2180;
      ov := iv(13 downto 0);
      ptr_deref_2182_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2182_gather_scatter
    process(tmp57_2153) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp57_2153;
      ov(63 downto 0) := iv;
      ptr_deref_2182_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2182_root_address_inst
    process(ptr_deref_2182_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2182_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2182_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_2201_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_2200;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2201_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2201_branch_req_0,
          ack0 => if_stmt_2201_branch_ack_0,
          ack1 => if_stmt_2201_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2232_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp77_2231;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2232_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2232_branch_req_0,
          ack0 => if_stmt_2232_branch_ack_0,
          ack1 => if_stmt_2232_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2280_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp89_2279;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2280_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2280_branch_req_0,
          ack0 => if_stmt_2280_branch_ack_0,
          ack1 => if_stmt_2280_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_2212_inst
    process(indvar_2095) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_2095, type_cast_2211_wire_constant, tmp_var);
      indvarx_xnext_2213 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2220_inst
    process(input_dim1x_x1x_xph_1967) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_1967, type_cast_2219_wire_constant, tmp_var);
      inc_2221 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2243_inst
    process(input_dim0x_x2x_xph_1973) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim0x_x2x_xph_1973, type_cast_2242_wire_constant, tmp_var);
      inc81_2244 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1999_inst
    process(mul_1995, conv12_1985) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul_1995, conv12_1985, tmp_var);
      add_2000 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2014_inst
    process(mul23_2010, tmp24_1889) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul23_2010, tmp24_1889, tmp_var);
      add25_2015 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2029_inst
    process(mul34_2025, tmp35_1922) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul34_2025, tmp35_1922, tmp_var);
      add36_2030 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2046_inst
    process(sub40_2041) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub40_2041, type_cast_2045_wire_constant, tmp_var);
      sext_2047 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2067_inst
    process(sub28_2062) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub28_2062, type_cast_2066_wire_constant, tmp_var);
      sext103_2068 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2086_inst
    process(conv46_2056, mul50_2082) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv46_2056, mul50_2082, tmp_var);
      add51_2087 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2116_inst
    process(mul16_2005, conv9102_2112) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul16_2005, conv9102_2112, tmp_var);
      add17_2117 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2121_inst
    process(mul52_2092, conv9102_2112) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul52_2092, conv9102_2112, tmp_var);
      add53_2122 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2194_inst
    process(conv65_2189) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv65_2189, type_cast_2193_wire_constant, tmp_var);
      add66_2195 <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2054_inst
    process(type_cast_2050_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2050_wire, type_cast_2053_wire_constant, tmp_var);
      ASHR_i32_i32_2054_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2075_inst
    process(type_cast_2071_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2071_wire, type_cast_2074_wire_constant, tmp_var);
      ASHR_i32_i32_2075_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2135_inst
    process(type_cast_2131_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2131_wire, type_cast_2134_wire_constant, tmp_var);
      ASHR_i32_i32_2135_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2166_inst
    process(type_cast_2162_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2162_wire, type_cast_2165_wire_constant, tmp_var);
      ASHR_i32_i32_2166_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2230_inst
    process(conv75_2226, tmp_1841) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv75_2226, tmp_1841, tmp_var);
      cmp77_2231 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2278_inst
    process(conv86_2274, div88_1964) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv86_2274, div88_1964, tmp_var);
      cmp89_2279 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1846_inst
    process(tmp_1841) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp_1841, type_cast_1845_wire_constant, tmp_var);
      div_1847 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1963_inst
    process(tmp87_1958) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp87_1958, type_cast_1962_wire_constant, tmp_var);
      div88_1964 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2249_inst
    process(tmp_1841) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp_1841, type_cast_2248_wire_constant, tmp_var);
      div83_2250 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2107_inst
    process(indvar_2095) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_2095, type_cast_2106_wire_constant, tmp_var);
      input_dim2x_x1_2108 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1994_inst
    process(tmp_1841, conv15_1990) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp_1841, conv15_1990, tmp_var);
      mul_1995 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2004_inst
    process(add_2000, tmp10_1863) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add_2000, tmp10_1863, tmp_var);
      mul16_2005 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2009_inst
    process(conv22_1877, conv15_1990) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv22_1877, conv15_1990, tmp_var);
      mul23_2010 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2024_inst
    process(conv33_1910, conv12_1985) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv33_1910, conv12_1985, tmp_var);
      mul34_2025 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2081_inst
    process(tmp47_1946, conv49_2077) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp47_1946, conv49_2077, tmp_var);
      mul50_2082 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2091_inst
    process(add51_2087, tmp44_1934) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add51_2087, tmp44_1934, tmp_var);
      mul52_2092 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2040_inst
    process(sub39_2035) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(sub39_2035, type_cast_2039_wire_constant, tmp_var);
      sub40_2041 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2061_inst
    process(sub_2020) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(sub_2020, type_cast_2060_wire_constant, tmp_var);
      sub28_2062 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2127_inst
    process(add17_2117) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add17_2117, type_cast_2126_wire_constant, tmp_var);
      sext105_2128 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2158_inst
    process(add53_2122) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add53_2122, type_cast_2157_wire_constant, tmp_var);
      sext106_2159 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_2019_inst
    process(add25_2015, conv27_1896) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(add25_2015, conv27_1896, tmp_var);
      sub_2020 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_2034_inst
    process(add36_2030, conv27_1896) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(add36_2030, conv27_1896, tmp_var);
      sub39_2035 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_2199_inst
    process(add66_2195, tmp10_1863) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add66_2195, tmp10_1863, tmp_var);
      cmp_2200 <= tmp_var; --
    end process;
    -- shared split operator group (35) : array_obj_ref_2147_index_offset 
    ApIntAdd_group_35: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_2146_scaled;
      array_obj_ref_2147_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2147_index_offset_req_0;
      array_obj_ref_2147_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2147_index_offset_req_1;
      array_obj_ref_2147_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_35_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_35_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_35",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 35
    -- shared split operator group (36) : array_obj_ref_2178_index_offset 
    ApIntAdd_group_36: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom61_2177_scaled;
      array_obj_ref_2178_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2178_index_offset_req_0;
      array_obj_ref_2178_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2178_index_offset_req_1;
      array_obj_ref_2178_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_36_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_36_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_36",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 36
    -- unary operator type_cast_1983_inst
    process(input_dim1x_x1x_xph_1967) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim1x_x1x_xph_1967, tmp_var);
      type_cast_1983_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1988_inst
    process(input_dim0x_x2x_xph_1973) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim0x_x2x_xph_1973, tmp_var);
      type_cast_1988_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2140_inst
    process(shr_2137) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr_2137, tmp_var);
      type_cast_2140_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2171_inst
    process(shr60_2168) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr60_2168, tmp_var);
      type_cast_2171_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2187_inst
    process(input_dim2x_x1_2108) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim2x_x1_2108, tmp_var);
      type_cast_2187_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2224_inst
    process(inc_2221) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc_2221, tmp_var);
      type_cast_2224_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2272_inst
    process(input_dim0x_x0_2263) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim0x_x0_2263, tmp_var);
      type_cast_2272_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : LOAD_padding_1891_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_padding_1891_load_0_req_0;
      LOAD_padding_1891_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_padding_1891_load_0_req_1;
      LOAD_padding_1891_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_padding_1891_word_address_0;
      LOAD_padding_1891_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_7_lr_req(0),
          mack => memory_space_7_lr_ack(0),
          maddr => memory_space_7_lr_addr(0 downto 0),
          mtag => memory_space_7_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 8,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_7_lc_req(0),
          mack => memory_space_7_lc_ack(0),
          mdata => memory_space_7_lc_data(7 downto 0),
          mtag => memory_space_7_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_1862_load_0 ptr_deref_1840_load_0 ptr_deref_1957_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(20 downto 0);
      signal data_out: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_1862_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_1840_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1957_load_0_req_0;
      ptr_deref_1862_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_1840_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1957_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_1862_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_1840_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1957_load_0_req_1;
      ptr_deref_1862_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_1840_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1957_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      LoadGroup1_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1862_word_address_0 & ptr_deref_1840_word_address_0 & ptr_deref_1957_word_address_0;
      ptr_deref_1862_data_0 <= data_out(95 downto 64);
      ptr_deref_1840_data_0 <= data_out(63 downto 32);
      ptr_deref_1957_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 7,
        num_reqs => 3,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(6 downto 0),
          mtag => memory_space_1_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 32,
        num_reqs => 3,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(31 downto 0),
          mtag => memory_space_1_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : ptr_deref_1905_load_0 ptr_deref_1872_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1905_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1872_load_0_req_0;
      ptr_deref_1905_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1872_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1905_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1872_load_0_req_1;
      ptr_deref_1905_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1872_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup2_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup2_gI: SplitGuardInterface generic map(name => "LoadGroup2_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1905_word_address_0 & ptr_deref_1872_word_address_0;
      ptr_deref_1905_data_0 <= data_out(15 downto 8);
      ptr_deref_1872_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup2", addr_width => 1,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_8_lr_req(0),
          mack => memory_space_8_lr_ack(0),
          maddr => memory_space_8_lr_addr(0 downto 0),
          mtag => memory_space_8_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup2 load-complete ",
        data_width => 8,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_8_lc_req(0),
          mack => memory_space_8_lc_ack(0),
          mdata => memory_space_8_lc_data(7 downto 0),
          mtag => memory_space_8_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared load operator group (3) : ptr_deref_1921_load_0 ptr_deref_1888_load_0 
    LoadGroup3: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1921_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1888_load_0_req_0;
      ptr_deref_1921_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1888_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1921_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1888_load_0_req_1;
      ptr_deref_1921_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1888_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup3_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup3_gI: SplitGuardInterface generic map(name => "LoadGroup3_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1921_word_address_0 & ptr_deref_1888_word_address_0;
      ptr_deref_1921_data_0 <= data_out(63 downto 32);
      ptr_deref_1888_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup3", addr_width => 7,
        num_reqs => 2,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(6 downto 0),
          mtag => memory_space_2_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup3 load-complete ",
        data_width => 32,
        num_reqs => 2,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(31 downto 0),
          mtag => memory_space_2_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 3
    -- shared load operator group (4) : ptr_deref_1933_load_0 ptr_deref_1945_load_0 
    LoadGroup4: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1933_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1945_load_0_req_0;
      ptr_deref_1933_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1945_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1933_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1945_load_0_req_1;
      ptr_deref_1933_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1945_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup4_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup4_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup4_gI: SplitGuardInterface generic map(name => "LoadGroup4_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1933_word_address_0 & ptr_deref_1945_word_address_0;
      ptr_deref_1933_data_0 <= data_out(63 downto 32);
      ptr_deref_1945_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup4", addr_width => 7,
        num_reqs => 2,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(6 downto 0),
          mtag => memory_space_3_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup4 load-complete ",
        data_width => 32,
        num_reqs => 2,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(31 downto 0),
          mtag => memory_space_3_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 4
    -- shared load operator group (5) : ptr_deref_2152_load_0 
    LoadGroup5: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2152_load_0_req_0;
      ptr_deref_2152_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2152_load_0_req_1;
      ptr_deref_2152_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup5_gI: SplitGuardInterface generic map(name => "LoadGroup5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2152_word_address_0;
      ptr_deref_2152_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup5", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_4_lr_req(0),
          mack => memory_space_4_lr_ack(0),
          maddr => memory_space_4_lr_addr(13 downto 0),
          mtag => memory_space_4_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup5 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_4_lc_req(0),
          mack => memory_space_4_lc_ack(0),
          mdata => memory_space_4_lc_data(63 downto 0),
          mtag => memory_space_4_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 5
    -- shared store operator group (0) : ptr_deref_2182_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2182_store_0_req_0;
      ptr_deref_2182_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2182_store_0_req_1;
      ptr_deref_2182_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_2182_word_address_0;
      data_in <= ptr_deref_2182_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_6_sr_req(0),
          mack => memory_space_6_sr_ack(0),
          maddr => memory_space_6_sr_addr(13 downto 0),
          mdata => memory_space_6_sr_data(63 downto 0),
          mtag => memory_space_6_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_6_sc_req(0),
          mack => memory_space_6_sc_ack(0),
          mtag => memory_space_6_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block1_start_1827_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block1_start_1827_inst_req_0;
      RPIPE_Block1_start_1827_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block1_start_1827_inst_req_1;
      RPIPE_Block1_start_1827_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call_1828 <= data_out(15 downto 0);
      Block1_start_read_0_gI: SplitGuardInterface generic map(name => "Block1_start_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block1_start_read_0: InputPortRevised -- 
        generic map ( name => "Block1_start_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block1_start_pipe_read_req(0),
          oack => Block1_start_pipe_read_ack(0),
          odata => Block1_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block1_done_2288_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block1_done_2288_inst_req_0;
      WPIPE_Block1_done_2288_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block1_done_2288_inst_req_1;
      WPIPE_Block1_done_2288_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= call_1828;
      Block1_done_write_0_gI: SplitGuardInterface generic map(name => "Block1_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block1_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block1_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block1_done_pipe_write_req(0),
          oack => Block1_done_pipe_write_ack(0),
          odata => Block1_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeB_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeC is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_7_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_8_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_8_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_8_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_8_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_8_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_8_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_4_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_4_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_6_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_6_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_sc_tag :  in  std_logic_vector(0 downto 0);
    Block2_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block2_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block2_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block2_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block2_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block2_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeC;
architecture convTransposeC_arch of convTransposeC is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeC_CP_6423_start: Boolean;
  signal convTransposeC_CP_6423_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal type_cast_2696_inst_ack_1 : boolean;
  signal type_cast_2696_inst_req_1 : boolean;
  signal type_cast_2450_inst_req_0 : boolean;
  signal type_cast_2659_inst_ack_1 : boolean;
  signal addr_of_2650_final_reg_req_1 : boolean;
  signal WPIPE_Block2_done_2737_inst_ack_1 : boolean;
  signal WPIPE_Block2_done_2737_inst_req_1 : boolean;
  signal type_cast_2659_inst_req_1 : boolean;
  signal addr_of_2650_final_reg_ack_1 : boolean;
  signal ptr_deref_2653_store_0_ack_0 : boolean;
  signal addr_of_2650_final_reg_ack_0 : boolean;
  signal type_cast_2659_inst_ack_0 : boolean;
  signal type_cast_2722_inst_ack_1 : boolean;
  signal ptr_deref_2653_store_0_req_0 : boolean;
  signal addr_of_2650_final_reg_req_0 : boolean;
  signal type_cast_2450_inst_ack_0 : boolean;
  signal type_cast_2659_inst_req_0 : boolean;
  signal type_cast_2722_inst_req_0 : boolean;
  signal if_stmt_2729_branch_ack_0 : boolean;
  signal type_cast_2722_inst_ack_0 : boolean;
  signal if_stmt_2672_branch_req_0 : boolean;
  signal type_cast_2448_inst_req_0 : boolean;
  signal type_cast_2448_inst_ack_0 : boolean;
  signal phi_stmt_2438_req_1 : boolean;
  signal type_cast_2441_inst_ack_0 : boolean;
  signal phi_stmt_2445_req_0 : boolean;
  signal type_cast_2572_inst_req_0 : boolean;
  signal if_stmt_2672_branch_ack_1 : boolean;
  signal if_stmt_2672_branch_ack_0 : boolean;
  signal if_stmt_2729_branch_req_0 : boolean;
  signal type_cast_2448_inst_req_1 : boolean;
  signal type_cast_2448_inst_ack_1 : boolean;
  signal type_cast_2441_inst_req_1 : boolean;
  signal type_cast_2441_inst_req_0 : boolean;
  signal phi_stmt_2445_req_1 : boolean;
  signal type_cast_2572_inst_ack_0 : boolean;
  signal type_cast_2441_inst_ack_1 : boolean;
  signal if_stmt_2729_branch_ack_1 : boolean;
  signal phi_stmt_2438_req_0 : boolean;
  signal type_cast_2722_inst_req_1 : boolean;
  signal phi_stmt_2438_ack_0 : boolean;
  signal phi_stmt_2445_ack_0 : boolean;
  signal type_cast_2450_inst_req_1 : boolean;
  signal type_cast_2705_inst_req_0 : boolean;
  signal type_cast_2705_inst_ack_0 : boolean;
  signal type_cast_2572_inst_ack_1 : boolean;
  signal phi_stmt_2566_req_1 : boolean;
  signal phi_stmt_2566_ack_0 : boolean;
  signal phi_stmt_2566_req_0 : boolean;
  signal type_cast_2572_inst_req_1 : boolean;
  signal type_cast_2450_inst_ack_1 : boolean;
  signal type_cast_2705_inst_req_1 : boolean;
  signal type_cast_2705_inst_ack_1 : boolean;
  signal RPIPE_Block2_start_2298_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2298_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2298_inst_req_1 : boolean;
  signal RPIPE_Block2_start_2298_inst_ack_1 : boolean;
  signal ptr_deref_2311_load_0_req_0 : boolean;
  signal ptr_deref_2311_load_0_ack_0 : boolean;
  signal ptr_deref_2311_load_0_req_1 : boolean;
  signal ptr_deref_2311_load_0_ack_1 : boolean;
  signal type_cast_2321_inst_req_0 : boolean;
  signal type_cast_2321_inst_ack_0 : boolean;
  signal type_cast_2321_inst_req_1 : boolean;
  signal type_cast_2321_inst_ack_1 : boolean;
  signal ptr_deref_2333_load_0_req_0 : boolean;
  signal ptr_deref_2333_load_0_ack_0 : boolean;
  signal ptr_deref_2333_load_0_req_1 : boolean;
  signal ptr_deref_2333_load_0_ack_1 : boolean;
  signal ptr_deref_2345_load_0_req_0 : boolean;
  signal ptr_deref_2345_load_0_ack_0 : boolean;
  signal ptr_deref_2345_load_0_req_1 : boolean;
  signal ptr_deref_2345_load_0_ack_1 : boolean;
  signal ptr_deref_2355_load_0_req_0 : boolean;
  signal ptr_deref_2355_load_0_ack_0 : boolean;
  signal ptr_deref_2355_load_0_req_1 : boolean;
  signal ptr_deref_2355_load_0_ack_1 : boolean;
  signal type_cast_2359_inst_req_0 : boolean;
  signal type_cast_2359_inst_ack_0 : boolean;
  signal type_cast_2359_inst_req_1 : boolean;
  signal type_cast_2359_inst_ack_1 : boolean;
  signal ptr_deref_2371_load_0_req_0 : boolean;
  signal ptr_deref_2371_load_0_ack_0 : boolean;
  signal ptr_deref_2371_load_0_req_1 : boolean;
  signal ptr_deref_2371_load_0_ack_1 : boolean;
  signal LOAD_padding_2374_load_0_req_0 : boolean;
  signal LOAD_padding_2374_load_0_ack_0 : boolean;
  signal LOAD_padding_2374_load_0_req_1 : boolean;
  signal LOAD_padding_2374_load_0_ack_1 : boolean;
  signal type_cast_2378_inst_req_0 : boolean;
  signal type_cast_2378_inst_ack_0 : boolean;
  signal type_cast_2378_inst_req_1 : boolean;
  signal type_cast_2378_inst_ack_1 : boolean;
  signal ptr_deref_2388_load_0_req_0 : boolean;
  signal ptr_deref_2388_load_0_ack_0 : boolean;
  signal ptr_deref_2388_load_0_req_1 : boolean;
  signal ptr_deref_2388_load_0_ack_1 : boolean;
  signal type_cast_2392_inst_req_0 : boolean;
  signal type_cast_2696_inst_ack_0 : boolean;
  signal type_cast_2392_inst_ack_0 : boolean;
  signal WPIPE_Block2_done_2737_inst_ack_0 : boolean;
  signal type_cast_2392_inst_req_1 : boolean;
  signal type_cast_2696_inst_req_0 : boolean;
  signal type_cast_2392_inst_ack_1 : boolean;
  signal ptr_deref_2653_store_0_ack_1 : boolean;
  signal ptr_deref_2653_store_0_req_1 : boolean;
  signal ptr_deref_2404_load_0_req_0 : boolean;
  signal ptr_deref_2404_load_0_ack_0 : boolean;
  signal ptr_deref_2404_load_0_req_1 : boolean;
  signal ptr_deref_2404_load_0_ack_1 : boolean;
  signal ptr_deref_2416_load_0_req_0 : boolean;
  signal ptr_deref_2416_load_0_ack_0 : boolean;
  signal ptr_deref_2416_load_0_req_1 : boolean;
  signal ptr_deref_2416_load_0_ack_1 : boolean;
  signal ptr_deref_2428_load_0_req_0 : boolean;
  signal ptr_deref_2428_load_0_ack_0 : boolean;
  signal ptr_deref_2428_load_0_req_1 : boolean;
  signal ptr_deref_2428_load_0_ack_1 : boolean;
  signal type_cast_2455_inst_req_0 : boolean;
  signal type_cast_2455_inst_ack_0 : boolean;
  signal type_cast_2455_inst_req_1 : boolean;
  signal type_cast_2455_inst_ack_1 : boolean;
  signal type_cast_2460_inst_req_0 : boolean;
  signal type_cast_2460_inst_ack_0 : boolean;
  signal type_cast_2460_inst_req_1 : boolean;
  signal type_cast_2460_inst_ack_1 : boolean;
  signal type_cast_2582_inst_req_0 : boolean;
  signal type_cast_2582_inst_ack_0 : boolean;
  signal type_cast_2582_inst_req_1 : boolean;
  signal type_cast_2582_inst_ack_1 : boolean;
  signal type_cast_2612_inst_req_0 : boolean;
  signal type_cast_2612_inst_ack_0 : boolean;
  signal type_cast_2612_inst_req_1 : boolean;
  signal type_cast_2612_inst_ack_1 : boolean;
  signal array_obj_ref_2618_index_offset_req_0 : boolean;
  signal array_obj_ref_2618_index_offset_ack_0 : boolean;
  signal array_obj_ref_2618_index_offset_req_1 : boolean;
  signal array_obj_ref_2618_index_offset_ack_1 : boolean;
  signal addr_of_2619_final_reg_req_0 : boolean;
  signal addr_of_2619_final_reg_ack_0 : boolean;
  signal addr_of_2619_final_reg_req_1 : boolean;
  signal addr_of_2619_final_reg_ack_1 : boolean;
  signal WPIPE_Block2_done_2737_inst_req_0 : boolean;
  signal ptr_deref_2623_load_0_req_0 : boolean;
  signal ptr_deref_2623_load_0_ack_0 : boolean;
  signal ptr_deref_2623_load_0_req_1 : boolean;
  signal ptr_deref_2623_load_0_ack_1 : boolean;
  signal type_cast_2643_inst_req_0 : boolean;
  signal type_cast_2643_inst_ack_0 : boolean;
  signal type_cast_2643_inst_req_1 : boolean;
  signal type_cast_2643_inst_ack_1 : boolean;
  signal array_obj_ref_2649_index_offset_req_0 : boolean;
  signal array_obj_ref_2649_index_offset_ack_0 : boolean;
  signal array_obj_ref_2649_index_offset_req_1 : boolean;
  signal array_obj_ref_2649_index_offset_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeC_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeC_CP_6423_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeC_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeC_CP_6423_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeC_CP_6423_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeC_CP_6423_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeC_CP_6423: Block -- control-path 
    signal convTransposeC_CP_6423_elements: BooleanArray(92 downto 0);
    -- 
  begin -- 
    convTransposeC_CP_6423_elements(0) <= convTransposeC_CP_6423_start;
    convTransposeC_CP_6423_symbol <= convTransposeC_CP_6423_elements(70);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_2296/$entry
      -- CP-element group 0: 	 branch_block_stmt_2296/branch_block_stmt_2296__entry__
      -- CP-element group 0: 	 branch_block_stmt_2296/assign_stmt_2299__entry__
      -- CP-element group 0: 	 branch_block_stmt_2296/assign_stmt_2299/$entry
      -- CP-element group 0: 	 branch_block_stmt_2296/assign_stmt_2299/RPIPE_Block2_start_2298_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_2296/assign_stmt_2299/RPIPE_Block2_start_2298_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_2296/assign_stmt_2299/RPIPE_Block2_start_2298_Sample/rr
      -- 
    rr_6471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(0), ack => RPIPE_Block2_start_2298_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_2296/assign_stmt_2299/RPIPE_Block2_start_2298_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_2296/assign_stmt_2299/RPIPE_Block2_start_2298_update_start_
      -- CP-element group 1: 	 branch_block_stmt_2296/assign_stmt_2299/RPIPE_Block2_start_2298_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_2296/assign_stmt_2299/RPIPE_Block2_start_2298_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_2296/assign_stmt_2299/RPIPE_Block2_start_2298_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2296/assign_stmt_2299/RPIPE_Block2_start_2298_Update/cr
      -- 
    ra_6472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2298_inst_ack_0, ack => convTransposeC_CP_6423_elements(1)); -- 
    cr_6476_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6476_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(1), ack => RPIPE_Block2_start_2298_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  place  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2: 	22 
    -- CP-element group 2: 	9 
    -- CP-element group 2: 	24 
    -- CP-element group 2: 	25 
    -- CP-element group 2: 	26 
    -- CP-element group 2: 	27 
    -- CP-element group 2: 	28 
    -- CP-element group 2: 	7 
    -- CP-element group 2: 	20 
    -- CP-element group 2: 	10 
    -- CP-element group 2: 	29 
    -- CP-element group 2: 	30 
    -- CP-element group 2: 	21 
    -- CP-element group 2: 	14 
    -- CP-element group 2: 	12 
    -- CP-element group 2: 	11 
    -- CP-element group 2: 	15 
    -- CP-element group 2: 	16 
    -- CP-element group 2: 	17 
    -- CP-element group 2: 	18 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	4 
    -- CP-element group 2: 	6 
    -- CP-element group 2:  members (265) 
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2299__exit__
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435__entry__
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2299/$exit
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2299/RPIPE_Block2_start_2298_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2299/RPIPE_Block2_start_2298_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2299/RPIPE_Block2_start_2298_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2311_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2311_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2311_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2311_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2311_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2311_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2311_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2311_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2311_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2311_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2311_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2311_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2311_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2311_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2311_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2311_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2311_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2311_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2311_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2311_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2311_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2311_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2311_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2311_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2311_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2311_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/type_cast_2321_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/type_cast_2321_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/type_cast_2321_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2333_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2333_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2333_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2333_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2333_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2333_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2333_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2333_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2333_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2333_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2333_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2333_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2333_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2333_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2333_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2333_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2333_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2333_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2333_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2333_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2333_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2333_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2333_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2333_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2333_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2333_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2345_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2345_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2345_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2345_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2345_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2345_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2345_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2345_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2345_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2345_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2345_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2345_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2345_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2345_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2345_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2345_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2345_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2345_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2345_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2345_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2345_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2345_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2345_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2345_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2345_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2345_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2355_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2355_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2355_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2355_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2355_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2355_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2355_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2355_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2355_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2355_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2355_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2355_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2355_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2355_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2355_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2355_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2355_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2355_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2355_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2355_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2355_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2355_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2355_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2355_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2355_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2355_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/type_cast_2359_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/type_cast_2359_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/type_cast_2359_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2371_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2416_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2371_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2371_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2371_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2371_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2371_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2371_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2371_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2371_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2371_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2371_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2371_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2371_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2371_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2371_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2371_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2371_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2371_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2371_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2371_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2371_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2371_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2371_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2371_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2371_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2371_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/LOAD_padding_2374_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/LOAD_padding_2374_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/LOAD_padding_2374_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/LOAD_padding_2374_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/LOAD_padding_2374_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/LOAD_padding_2374_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/LOAD_padding_2374_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/LOAD_padding_2374_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/LOAD_padding_2374_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/LOAD_padding_2374_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/LOAD_padding_2374_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/LOAD_padding_2374_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/type_cast_2378_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/type_cast_2378_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/type_cast_2378_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2388_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2388_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2388_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2388_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2388_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2388_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2388_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2388_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2388_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2388_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2388_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2388_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2388_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2388_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2388_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2388_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2388_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2388_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2388_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2388_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2388_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2388_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2388_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2388_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2388_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2388_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/type_cast_2392_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/type_cast_2392_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/type_cast_2392_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2404_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2404_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2404_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2404_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2404_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2404_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2404_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2404_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2404_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2404_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2404_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2404_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2404_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2404_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2404_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2404_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2404_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2404_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2404_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2404_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2404_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2404_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2404_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2404_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2404_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2404_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2416_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2416_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2416_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2416_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2416_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2416_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2416_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2416_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2416_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2416_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2416_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2416_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2416_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2416_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2416_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2416_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2416_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2416_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2416_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2416_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2416_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2416_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2416_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2416_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2416_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2428_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2428_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2428_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2428_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2428_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2428_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2428_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2428_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2428_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2428_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2428_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2428_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2428_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2428_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2428_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2428_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2428_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2428_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2428_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2428_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2428_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2428_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2428_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2428_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2428_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2428_Update/word_access_complete/word_0/cr
      -- 
    ca_6477_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2298_inst_ack_1, ack => convTransposeC_CP_6423_elements(2)); -- 
    rr_6513_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6513_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(2), ack => ptr_deref_2311_load_0_req_0); -- 
    cr_6524_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6524_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(2), ack => ptr_deref_2311_load_0_req_1); -- 
    cr_6543_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6543_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(2), ack => type_cast_2321_inst_req_1); -- 
    rr_6577_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6577_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(2), ack => ptr_deref_2333_load_0_req_0); -- 
    cr_6588_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6588_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(2), ack => ptr_deref_2333_load_0_req_1); -- 
    rr_6627_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6627_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(2), ack => ptr_deref_2345_load_0_req_0); -- 
    cr_6638_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6638_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(2), ack => ptr_deref_2345_load_0_req_1); -- 
    rr_6677_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6677_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(2), ack => ptr_deref_2355_load_0_req_0); -- 
    cr_6688_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6688_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(2), ack => ptr_deref_2355_load_0_req_1); -- 
    cr_6707_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6707_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(2), ack => type_cast_2359_inst_req_1); -- 
    rr_6741_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6741_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(2), ack => ptr_deref_2371_load_0_req_0); -- 
    cr_6752_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6752_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(2), ack => ptr_deref_2371_load_0_req_1); -- 
    rr_6774_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6774_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(2), ack => LOAD_padding_2374_load_0_req_0); -- 
    cr_6785_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6785_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(2), ack => LOAD_padding_2374_load_0_req_1); -- 
    cr_6804_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6804_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(2), ack => type_cast_2378_inst_req_1); -- 
    rr_6838_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6838_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(2), ack => ptr_deref_2388_load_0_req_0); -- 
    cr_6849_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6849_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(2), ack => ptr_deref_2388_load_0_req_1); -- 
    cr_6868_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6868_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(2), ack => type_cast_2392_inst_req_1); -- 
    rr_6902_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6902_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(2), ack => ptr_deref_2404_load_0_req_0); -- 
    cr_6913_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6913_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(2), ack => ptr_deref_2404_load_0_req_1); -- 
    rr_6952_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6952_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(2), ack => ptr_deref_2416_load_0_req_0); -- 
    cr_6963_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6963_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(2), ack => ptr_deref_2416_load_0_req_1); -- 
    rr_7002_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7002_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(2), ack => ptr_deref_2428_load_0_req_0); -- 
    cr_7013_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7013_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(2), ack => ptr_deref_2428_load_0_req_1); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (5) 
      -- CP-element group 3: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2311_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2311_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2311_Sample/word_access_start/$exit
      -- CP-element group 3: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2311_Sample/word_access_start/word_0/$exit
      -- CP-element group 3: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2311_Sample/word_access_start/word_0/ra
      -- 
    ra_6514_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2311_load_0_ack_0, ack => convTransposeC_CP_6423_elements(3)); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	2 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (12) 
      -- CP-element group 4: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2311_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2311_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2311_Update/word_access_complete/$exit
      -- CP-element group 4: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2311_Update/word_access_complete/word_0/$exit
      -- CP-element group 4: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2311_Update/word_access_complete/word_0/ca
      -- CP-element group 4: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2311_Update/ptr_deref_2311_Merge/$entry
      -- CP-element group 4: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2311_Update/ptr_deref_2311_Merge/$exit
      -- CP-element group 4: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2311_Update/ptr_deref_2311_Merge/merge_req
      -- CP-element group 4: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2311_Update/ptr_deref_2311_Merge/merge_ack
      -- CP-element group 4: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/type_cast_2321_sample_start_
      -- CP-element group 4: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/type_cast_2321_Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/type_cast_2321_Sample/rr
      -- 
    ca_6525_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2311_load_0_ack_1, ack => convTransposeC_CP_6423_elements(4)); -- 
    rr_6538_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6538_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(4), ack => type_cast_2321_inst_req_0); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/type_cast_2321_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/type_cast_2321_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/type_cast_2321_Sample/ra
      -- 
    ra_6539_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2321_inst_ack_0, ack => convTransposeC_CP_6423_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	2 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	31 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/type_cast_2321_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/type_cast_2321_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/type_cast_2321_Update/ca
      -- 
    ca_6544_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2321_inst_ack_1, ack => convTransposeC_CP_6423_elements(6)); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	2 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (5) 
      -- CP-element group 7: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2333_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2333_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2333_Sample/word_access_start/$exit
      -- CP-element group 7: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2333_Sample/word_access_start/word_0/$exit
      -- CP-element group 7: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2333_Sample/word_access_start/word_0/ra
      -- 
    ra_6578_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2333_load_0_ack_0, ack => convTransposeC_CP_6423_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	31 
    -- CP-element group 8:  members (9) 
      -- CP-element group 8: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2333_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2333_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2333_Update/word_access_complete/$exit
      -- CP-element group 8: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2333_Update/word_access_complete/word_0/$exit
      -- CP-element group 8: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2333_Update/word_access_complete/word_0/ca
      -- CP-element group 8: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2333_Update/ptr_deref_2333_Merge/$entry
      -- CP-element group 8: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2333_Update/ptr_deref_2333_Merge/$exit
      -- CP-element group 8: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2333_Update/ptr_deref_2333_Merge/merge_req
      -- CP-element group 8: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2333_Update/ptr_deref_2333_Merge/merge_ack
      -- 
    ca_6589_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2333_load_0_ack_1, ack => convTransposeC_CP_6423_elements(8)); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	2 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (5) 
      -- CP-element group 9: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2345_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2345_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2345_Sample/word_access_start/$exit
      -- CP-element group 9: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2345_Sample/word_access_start/word_0/$exit
      -- CP-element group 9: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2345_Sample/word_access_start/word_0/ra
      -- 
    ra_6628_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2345_load_0_ack_0, ack => convTransposeC_CP_6423_elements(9)); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	2 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	31 
    -- CP-element group 10:  members (9) 
      -- CP-element group 10: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2345_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2345_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2345_Update/word_access_complete/$exit
      -- CP-element group 10: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2345_Update/word_access_complete/word_0/$exit
      -- CP-element group 10: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2345_Update/word_access_complete/word_0/ca
      -- CP-element group 10: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2345_Update/ptr_deref_2345_Merge/$entry
      -- CP-element group 10: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2345_Update/ptr_deref_2345_Merge/$exit
      -- CP-element group 10: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2345_Update/ptr_deref_2345_Merge/merge_req
      -- CP-element group 10: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2345_Update/ptr_deref_2345_Merge/merge_ack
      -- 
    ca_6639_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2345_load_0_ack_1, ack => convTransposeC_CP_6423_elements(10)); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	2 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (5) 
      -- CP-element group 11: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2355_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2355_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2355_Sample/word_access_start/$exit
      -- CP-element group 11: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2355_Sample/word_access_start/word_0/$exit
      -- CP-element group 11: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2355_Sample/word_access_start/word_0/ra
      -- 
    ra_6678_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2355_load_0_ack_0, ack => convTransposeC_CP_6423_elements(11)); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	2 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (12) 
      -- CP-element group 12: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2355_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2355_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2355_Update/word_access_complete/$exit
      -- CP-element group 12: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2355_Update/word_access_complete/word_0/$exit
      -- CP-element group 12: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2355_Update/word_access_complete/word_0/ca
      -- CP-element group 12: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2355_Update/ptr_deref_2355_Merge/$entry
      -- CP-element group 12: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2355_Update/ptr_deref_2355_Merge/$exit
      -- CP-element group 12: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2355_Update/ptr_deref_2355_Merge/merge_req
      -- CP-element group 12: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2355_Update/ptr_deref_2355_Merge/merge_ack
      -- CP-element group 12: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/type_cast_2359_sample_start_
      -- CP-element group 12: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/type_cast_2359_Sample/$entry
      -- CP-element group 12: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/type_cast_2359_Sample/rr
      -- 
    ca_6689_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2355_load_0_ack_1, ack => convTransposeC_CP_6423_elements(12)); -- 
    rr_6702_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6702_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(12), ack => type_cast_2359_inst_req_0); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/type_cast_2359_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/type_cast_2359_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/type_cast_2359_Sample/ra
      -- 
    ra_6703_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2359_inst_ack_0, ack => convTransposeC_CP_6423_elements(13)); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	2 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	31 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/type_cast_2359_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/type_cast_2359_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/type_cast_2359_Update/ca
      -- 
    ca_6708_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2359_inst_ack_1, ack => convTransposeC_CP_6423_elements(14)); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	2 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (5) 
      -- CP-element group 15: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2371_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2371_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2371_Sample/word_access_start/$exit
      -- CP-element group 15: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2371_Sample/word_access_start/word_0/$exit
      -- CP-element group 15: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2371_Sample/word_access_start/word_0/ra
      -- 
    ra_6742_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2371_load_0_ack_0, ack => convTransposeC_CP_6423_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	2 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	31 
    -- CP-element group 16:  members (9) 
      -- CP-element group 16: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2371_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2371_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2371_Update/word_access_complete/$exit
      -- CP-element group 16: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2371_Update/word_access_complete/word_0/$exit
      -- CP-element group 16: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2371_Update/word_access_complete/word_0/ca
      -- CP-element group 16: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2371_Update/ptr_deref_2371_Merge/$entry
      -- CP-element group 16: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2371_Update/ptr_deref_2371_Merge/$exit
      -- CP-element group 16: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2371_Update/ptr_deref_2371_Merge/merge_req
      -- CP-element group 16: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2371_Update/ptr_deref_2371_Merge/merge_ack
      -- 
    ca_6753_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2371_load_0_ack_1, ack => convTransposeC_CP_6423_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	2 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (5) 
      -- CP-element group 17: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/LOAD_padding_2374_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/LOAD_padding_2374_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/LOAD_padding_2374_Sample/word_access_start/$exit
      -- CP-element group 17: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/LOAD_padding_2374_Sample/word_access_start/word_0/$exit
      -- CP-element group 17: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/LOAD_padding_2374_Sample/word_access_start/word_0/ra
      -- 
    ra_6775_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_padding_2374_load_0_ack_0, ack => convTransposeC_CP_6423_elements(17)); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	2 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (12) 
      -- CP-element group 18: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/LOAD_padding_2374_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/LOAD_padding_2374_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/LOAD_padding_2374_Update/word_access_complete/$exit
      -- CP-element group 18: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/LOAD_padding_2374_Update/word_access_complete/word_0/$exit
      -- CP-element group 18: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/LOAD_padding_2374_Update/word_access_complete/word_0/ca
      -- CP-element group 18: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/LOAD_padding_2374_Update/LOAD_padding_2374_Merge/$entry
      -- CP-element group 18: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/LOAD_padding_2374_Update/LOAD_padding_2374_Merge/$exit
      -- CP-element group 18: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/LOAD_padding_2374_Update/LOAD_padding_2374_Merge/merge_req
      -- CP-element group 18: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/LOAD_padding_2374_Update/LOAD_padding_2374_Merge/merge_ack
      -- CP-element group 18: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/type_cast_2378_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/type_cast_2378_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/type_cast_2378_Sample/rr
      -- 
    ca_6786_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_padding_2374_load_0_ack_1, ack => convTransposeC_CP_6423_elements(18)); -- 
    rr_6799_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6799_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(18), ack => type_cast_2378_inst_req_0); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/type_cast_2378_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/type_cast_2378_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/type_cast_2378_Sample/ra
      -- 
    ra_6800_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2378_inst_ack_0, ack => convTransposeC_CP_6423_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	2 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	31 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/type_cast_2378_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/type_cast_2378_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/type_cast_2378_Update/ca
      -- 
    ca_6805_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2378_inst_ack_1, ack => convTransposeC_CP_6423_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	2 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (5) 
      -- CP-element group 21: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2388_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2388_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2388_Sample/word_access_start/$exit
      -- CP-element group 21: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2388_Sample/word_access_start/word_0/$exit
      -- CP-element group 21: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2388_Sample/word_access_start/word_0/ra
      -- 
    ra_6839_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2388_load_0_ack_0, ack => convTransposeC_CP_6423_elements(21)); -- 
    -- CP-element group 22:  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	2 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (12) 
      -- CP-element group 22: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2388_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2388_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2388_Update/word_access_complete/$exit
      -- CP-element group 22: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2388_Update/word_access_complete/word_0/$exit
      -- CP-element group 22: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2388_Update/word_access_complete/word_0/ca
      -- CP-element group 22: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2388_Update/ptr_deref_2388_Merge/$entry
      -- CP-element group 22: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2388_Update/ptr_deref_2388_Merge/$exit
      -- CP-element group 22: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2388_Update/ptr_deref_2388_Merge/merge_req
      -- CP-element group 22: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2388_Update/ptr_deref_2388_Merge/merge_ack
      -- CP-element group 22: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/type_cast_2392_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/type_cast_2392_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/type_cast_2392_Sample/rr
      -- 
    ca_6850_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2388_load_0_ack_1, ack => convTransposeC_CP_6423_elements(22)); -- 
    rr_6863_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6863_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(22), ack => type_cast_2392_inst_req_0); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/type_cast_2392_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/type_cast_2392_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/type_cast_2392_Sample/ra
      -- 
    ra_6864_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2392_inst_ack_0, ack => convTransposeC_CP_6423_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	2 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	31 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/type_cast_2392_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/type_cast_2392_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/type_cast_2392_Update/ca
      -- 
    ca_6869_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2392_inst_ack_1, ack => convTransposeC_CP_6423_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	2 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (5) 
      -- CP-element group 25: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2404_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2404_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2404_Sample/word_access_start/$exit
      -- CP-element group 25: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2404_Sample/word_access_start/word_0/$exit
      -- CP-element group 25: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2404_Sample/word_access_start/word_0/ra
      -- 
    ra_6903_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2404_load_0_ack_0, ack => convTransposeC_CP_6423_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	2 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	31 
    -- CP-element group 26:  members (9) 
      -- CP-element group 26: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2404_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2404_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2404_Update/word_access_complete/$exit
      -- CP-element group 26: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2404_Update/word_access_complete/word_0/$exit
      -- CP-element group 26: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2404_Update/word_access_complete/word_0/ca
      -- CP-element group 26: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2404_Update/ptr_deref_2404_Merge/$entry
      -- CP-element group 26: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2404_Update/ptr_deref_2404_Merge/$exit
      -- CP-element group 26: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2404_Update/ptr_deref_2404_Merge/merge_req
      -- CP-element group 26: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2404_Update/ptr_deref_2404_Merge/merge_ack
      -- 
    ca_6914_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2404_load_0_ack_1, ack => convTransposeC_CP_6423_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	2 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (5) 
      -- CP-element group 27: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2416_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2416_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2416_Sample/word_access_start/$exit
      -- CP-element group 27: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2416_Sample/word_access_start/word_0/$exit
      -- CP-element group 27: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2416_Sample/word_access_start/word_0/ra
      -- 
    ra_6953_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2416_load_0_ack_0, ack => convTransposeC_CP_6423_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	2 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	31 
    -- CP-element group 28:  members (9) 
      -- CP-element group 28: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2416_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2416_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2416_Update/word_access_complete/$exit
      -- CP-element group 28: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2416_Update/word_access_complete/word_0/$exit
      -- CP-element group 28: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2416_Update/word_access_complete/word_0/ca
      -- CP-element group 28: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2416_Update/ptr_deref_2416_Merge/$entry
      -- CP-element group 28: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2416_Update/ptr_deref_2416_Merge/$exit
      -- CP-element group 28: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2416_Update/ptr_deref_2416_Merge/merge_req
      -- CP-element group 28: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2416_Update/ptr_deref_2416_Merge/merge_ack
      -- 
    ca_6964_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2416_load_0_ack_1, ack => convTransposeC_CP_6423_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	2 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (5) 
      -- CP-element group 29: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2428_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2428_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2428_Sample/word_access_start/$exit
      -- CP-element group 29: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2428_Sample/word_access_start/word_0/$exit
      -- CP-element group 29: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2428_Sample/word_access_start/word_0/ra
      -- 
    ra_7003_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2428_load_0_ack_0, ack => convTransposeC_CP_6423_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	2 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (9) 
      -- CP-element group 30: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2428_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2428_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2428_Update/word_access_complete/$exit
      -- CP-element group 30: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2428_Update/word_access_complete/word_0/$exit
      -- CP-element group 30: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2428_Update/word_access_complete/word_0/ca
      -- CP-element group 30: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2428_Update/ptr_deref_2428_Merge/$entry
      -- CP-element group 30: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2428_Update/ptr_deref_2428_Merge/$exit
      -- CP-element group 30: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2428_Update/ptr_deref_2428_Merge/merge_req
      -- CP-element group 30: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/ptr_deref_2428_Update/ptr_deref_2428_Merge/merge_ack
      -- 
    ca_7014_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2428_load_0_ack_1, ack => convTransposeC_CP_6423_elements(30)); -- 
    -- CP-element group 31:  join  fork  transition  place  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	8 
    -- CP-element group 31: 	24 
    -- CP-element group 31: 	26 
    -- CP-element group 31: 	28 
    -- CP-element group 31: 	20 
    -- CP-element group 31: 	10 
    -- CP-element group 31: 	30 
    -- CP-element group 31: 	14 
    -- CP-element group 31: 	16 
    -- CP-element group 31: 	6 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	71 
    -- CP-element group 31: 	72 
    -- CP-element group 31: 	73 
    -- CP-element group 31:  members (14) 
      -- CP-element group 31: 	 branch_block_stmt_2296/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2438/phi_stmt_2438_sources/$entry
      -- CP-element group 31: 	 branch_block_stmt_2296/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2445/phi_stmt_2445_sources/type_cast_2450/SplitProtocol/Sample/rr
      -- CP-element group 31: 	 branch_block_stmt_2296/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2445/phi_stmt_2445_sources/type_cast_2450/SplitProtocol/Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_2296/entry_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 31: 	 branch_block_stmt_2296/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2445/phi_stmt_2445_sources/type_cast_2450/SplitProtocol/Update/$entry
      -- CP-element group 31: 	 branch_block_stmt_2296/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2445/$entry
      -- CP-element group 31: 	 branch_block_stmt_2296/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2445/phi_stmt_2445_sources/$entry
      -- CP-element group 31: 	 branch_block_stmt_2296/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2438/$entry
      -- CP-element group 31: 	 branch_block_stmt_2296/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2445/phi_stmt_2445_sources/type_cast_2450/$entry
      -- CP-element group 31: 	 branch_block_stmt_2296/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2445/phi_stmt_2445_sources/type_cast_2450/SplitProtocol/Update/cr
      -- CP-element group 31: 	 branch_block_stmt_2296/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2445/phi_stmt_2445_sources/type_cast_2450/SplitProtocol/$entry
      -- CP-element group 31: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435__exit__
      -- CP-element group 31: 	 branch_block_stmt_2296/entry_whilex_xbodyx_xouter
      -- CP-element group 31: 	 branch_block_stmt_2296/assign_stmt_2308_to_assign_stmt_2435/$exit
      -- 
    rr_7431_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7431_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(31), ack => type_cast_2450_inst_req_0); -- 
    cr_7436_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7436_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(31), ack => type_cast_2450_inst_req_1); -- 
    convTransposeC_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= convTransposeC_CP_6423_elements(8) & convTransposeC_CP_6423_elements(24) & convTransposeC_CP_6423_elements(26) & convTransposeC_CP_6423_elements(28) & convTransposeC_CP_6423_elements(20) & convTransposeC_CP_6423_elements(10) & convTransposeC_CP_6423_elements(30) & convTransposeC_CP_6423_elements(14) & convTransposeC_CP_6423_elements(16) & convTransposeC_CP_6423_elements(6);
      gj_convTransposeC_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6423_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	86 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_2296/assign_stmt_2456_to_assign_stmt_2563/type_cast_2455_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_2296/assign_stmt_2456_to_assign_stmt_2563/type_cast_2455_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_2296/assign_stmt_2456_to_assign_stmt_2563/type_cast_2455_Sample/ra
      -- 
    ra_7031_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2455_inst_ack_0, ack => convTransposeC_CP_6423_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	86 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	36 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_2296/assign_stmt_2456_to_assign_stmt_2563/type_cast_2455_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_2296/assign_stmt_2456_to_assign_stmt_2563/type_cast_2455_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_2296/assign_stmt_2456_to_assign_stmt_2563/type_cast_2455_Update/ca
      -- 
    ca_7036_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2455_inst_ack_1, ack => convTransposeC_CP_6423_elements(33)); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	86 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_2296/assign_stmt_2456_to_assign_stmt_2563/type_cast_2460_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_2296/assign_stmt_2456_to_assign_stmt_2563/type_cast_2460_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_2296/assign_stmt_2456_to_assign_stmt_2563/type_cast_2460_Sample/ra
      -- 
    ra_7045_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2460_inst_ack_0, ack => convTransposeC_CP_6423_elements(34)); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	86 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_2296/assign_stmt_2456_to_assign_stmt_2563/type_cast_2460_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_2296/assign_stmt_2456_to_assign_stmt_2563/type_cast_2460_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_2296/assign_stmt_2456_to_assign_stmt_2563/type_cast_2460_Update/ca
      -- 
    ca_7050_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2460_inst_ack_1, ack => convTransposeC_CP_6423_elements(35)); -- 
    -- CP-element group 36:  join  transition  place  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	33 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	90 
    -- CP-element group 36:  members (6) 
      -- CP-element group 36: 	 branch_block_stmt_2296/assign_stmt_2456_to_assign_stmt_2563__exit__
      -- CP-element group 36: 	 branch_block_stmt_2296/whilex_xbodyx_xouter_whilex_xbody
      -- CP-element group 36: 	 branch_block_stmt_2296/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$entry
      -- CP-element group 36: 	 branch_block_stmt_2296/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2566/$entry
      -- CP-element group 36: 	 branch_block_stmt_2296/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2566/phi_stmt_2566_sources/$entry
      -- CP-element group 36: 	 branch_block_stmt_2296/assign_stmt_2456_to_assign_stmt_2563/$exit
      -- 
    convTransposeC_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_6423_elements(33) & convTransposeC_CP_6423_elements(35);
      gj_convTransposeC_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6423_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	92 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/type_cast_2582_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/type_cast_2582_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/type_cast_2582_Sample/ra
      -- 
    ra_7062_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2582_inst_ack_0, ack => convTransposeC_CP_6423_elements(37)); -- 
    -- CP-element group 38:  fork  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	92 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38: 	47 
    -- CP-element group 38:  members (9) 
      -- CP-element group 38: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/type_cast_2582_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/type_cast_2582_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/type_cast_2582_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/type_cast_2612_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/type_cast_2612_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/type_cast_2612_Sample/rr
      -- CP-element group 38: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/type_cast_2643_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/type_cast_2643_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/type_cast_2643_Sample/rr
      -- 
    ca_7067_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2582_inst_ack_1, ack => convTransposeC_CP_6423_elements(38)); -- 
    rr_7075_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7075_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(38), ack => type_cast_2612_inst_req_0); -- 
    rr_7185_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7185_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(38), ack => type_cast_2643_inst_req_0); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/type_cast_2612_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/type_cast_2612_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/type_cast_2612_Sample/ra
      -- 
    ra_7076_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2612_inst_ack_0, ack => convTransposeC_CP_6423_elements(39)); -- 
    -- CP-element group 40:  transition  input  output  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	92 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (16) 
      -- CP-element group 40: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/type_cast_2612_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/type_cast_2612_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/type_cast_2612_Update/ca
      -- CP-element group 40: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/array_obj_ref_2618_index_resized_1
      -- CP-element group 40: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/array_obj_ref_2618_index_scaled_1
      -- CP-element group 40: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/array_obj_ref_2618_index_computed_1
      -- CP-element group 40: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/array_obj_ref_2618_index_resize_1/$entry
      -- CP-element group 40: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/array_obj_ref_2618_index_resize_1/$exit
      -- CP-element group 40: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/array_obj_ref_2618_index_resize_1/index_resize_req
      -- CP-element group 40: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/array_obj_ref_2618_index_resize_1/index_resize_ack
      -- CP-element group 40: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/array_obj_ref_2618_index_scale_1/$entry
      -- CP-element group 40: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/array_obj_ref_2618_index_scale_1/$exit
      -- CP-element group 40: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/array_obj_ref_2618_index_scale_1/scale_rename_req
      -- CP-element group 40: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/array_obj_ref_2618_index_scale_1/scale_rename_ack
      -- CP-element group 40: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/array_obj_ref_2618_final_index_sum_regn_Sample/$entry
      -- CP-element group 40: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/array_obj_ref_2618_final_index_sum_regn_Sample/req
      -- 
    ca_7081_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2612_inst_ack_1, ack => convTransposeC_CP_6423_elements(40)); -- 
    req_7106_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7106_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(40), ack => array_obj_ref_2618_index_offset_req_0); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	58 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/array_obj_ref_2618_final_index_sum_regn_sample_complete
      -- CP-element group 41: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/array_obj_ref_2618_final_index_sum_regn_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/array_obj_ref_2618_final_index_sum_regn_Sample/ack
      -- 
    ack_7107_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2618_index_offset_ack_0, ack => convTransposeC_CP_6423_elements(41)); -- 
    -- CP-element group 42:  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	92 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (11) 
      -- CP-element group 42: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/addr_of_2619_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/array_obj_ref_2618_root_address_calculated
      -- CP-element group 42: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/array_obj_ref_2618_offset_calculated
      -- CP-element group 42: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/array_obj_ref_2618_final_index_sum_regn_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/array_obj_ref_2618_final_index_sum_regn_Update/ack
      -- CP-element group 42: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/array_obj_ref_2618_base_plus_offset/$entry
      -- CP-element group 42: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/array_obj_ref_2618_base_plus_offset/$exit
      -- CP-element group 42: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/array_obj_ref_2618_base_plus_offset/sum_rename_req
      -- CP-element group 42: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/array_obj_ref_2618_base_plus_offset/sum_rename_ack
      -- CP-element group 42: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/addr_of_2619_request/$entry
      -- CP-element group 42: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/addr_of_2619_request/req
      -- 
    ack_7112_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2618_index_offset_ack_1, ack => convTransposeC_CP_6423_elements(42)); -- 
    req_7121_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7121_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(42), ack => addr_of_2619_final_reg_req_0); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/addr_of_2619_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/addr_of_2619_request/$exit
      -- CP-element group 43: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/addr_of_2619_request/ack
      -- 
    ack_7122_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2619_final_reg_ack_0, ack => convTransposeC_CP_6423_elements(43)); -- 
    -- CP-element group 44:  join  fork  transition  input  output  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	92 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (24) 
      -- CP-element group 44: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/addr_of_2619_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/addr_of_2619_complete/$exit
      -- CP-element group 44: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/addr_of_2619_complete/ack
      -- CP-element group 44: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2623_sample_start_
      -- CP-element group 44: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2623_base_address_calculated
      -- CP-element group 44: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2623_word_address_calculated
      -- CP-element group 44: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2623_root_address_calculated
      -- CP-element group 44: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2623_base_address_resized
      -- CP-element group 44: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2623_base_addr_resize/$entry
      -- CP-element group 44: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2623_base_addr_resize/$exit
      -- CP-element group 44: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2623_base_addr_resize/base_resize_req
      -- CP-element group 44: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2623_base_addr_resize/base_resize_ack
      -- CP-element group 44: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2623_base_plus_offset/$entry
      -- CP-element group 44: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2623_base_plus_offset/$exit
      -- CP-element group 44: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2623_base_plus_offset/sum_rename_req
      -- CP-element group 44: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2623_base_plus_offset/sum_rename_ack
      -- CP-element group 44: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2623_word_addrgen/$entry
      -- CP-element group 44: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2623_word_addrgen/$exit
      -- CP-element group 44: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2623_word_addrgen/root_register_req
      -- CP-element group 44: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2623_word_addrgen/root_register_ack
      -- CP-element group 44: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2623_Sample/$entry
      -- CP-element group 44: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2623_Sample/word_access_start/$entry
      -- CP-element group 44: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2623_Sample/word_access_start/word_0/$entry
      -- CP-element group 44: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2623_Sample/word_access_start/word_0/rr
      -- 
    ack_7127_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2619_final_reg_ack_1, ack => convTransposeC_CP_6423_elements(44)); -- 
    rr_7160_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7160_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(44), ack => ptr_deref_2623_load_0_req_0); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	44 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (5) 
      -- CP-element group 45: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2623_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2623_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2623_Sample/word_access_start/$exit
      -- CP-element group 45: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2623_Sample/word_access_start/word_0/$exit
      -- CP-element group 45: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2623_Sample/word_access_start/word_0/ra
      -- 
    ra_7161_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2623_load_0_ack_0, ack => convTransposeC_CP_6423_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	92 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	53 
    -- CP-element group 46:  members (9) 
      -- CP-element group 46: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2623_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2623_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2623_Update/word_access_complete/$exit
      -- CP-element group 46: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2623_Update/word_access_complete/word_0/$exit
      -- CP-element group 46: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2623_Update/word_access_complete/word_0/ca
      -- CP-element group 46: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2623_Update/ptr_deref_2623_Merge/$entry
      -- CP-element group 46: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2623_Update/ptr_deref_2623_Merge/$exit
      -- CP-element group 46: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2623_Update/ptr_deref_2623_Merge/merge_req
      -- CP-element group 46: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2623_Update/ptr_deref_2623_Merge/merge_ack
      -- 
    ca_7172_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2623_load_0_ack_1, ack => convTransposeC_CP_6423_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	38 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/type_cast_2643_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/type_cast_2643_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/type_cast_2643_Sample/ra
      -- 
    ra_7186_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2643_inst_ack_0, ack => convTransposeC_CP_6423_elements(47)); -- 
    -- CP-element group 48:  transition  input  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	92 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (16) 
      -- CP-element group 48: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/type_cast_2643_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/type_cast_2643_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/type_cast_2643_Update/ca
      -- CP-element group 48: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/array_obj_ref_2649_index_resized_1
      -- CP-element group 48: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/array_obj_ref_2649_index_scaled_1
      -- CP-element group 48: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/array_obj_ref_2649_index_computed_1
      -- CP-element group 48: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/array_obj_ref_2649_index_resize_1/$entry
      -- CP-element group 48: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/array_obj_ref_2649_index_resize_1/$exit
      -- CP-element group 48: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/array_obj_ref_2649_index_resize_1/index_resize_req
      -- CP-element group 48: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/array_obj_ref_2649_index_resize_1/index_resize_ack
      -- CP-element group 48: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/array_obj_ref_2649_index_scale_1/$entry
      -- CP-element group 48: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/array_obj_ref_2649_index_scale_1/$exit
      -- CP-element group 48: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/array_obj_ref_2649_index_scale_1/scale_rename_req
      -- CP-element group 48: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/array_obj_ref_2649_index_scale_1/scale_rename_ack
      -- CP-element group 48: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/array_obj_ref_2649_final_index_sum_regn_Sample/$entry
      -- CP-element group 48: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/array_obj_ref_2649_final_index_sum_regn_Sample/req
      -- 
    ca_7191_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2643_inst_ack_1, ack => convTransposeC_CP_6423_elements(48)); -- 
    req_7216_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7216_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(48), ack => array_obj_ref_2649_index_offset_req_0); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	58 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/array_obj_ref_2649_final_index_sum_regn_sample_complete
      -- CP-element group 49: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/array_obj_ref_2649_final_index_sum_regn_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/array_obj_ref_2649_final_index_sum_regn_Sample/ack
      -- 
    ack_7217_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2649_index_offset_ack_0, ack => convTransposeC_CP_6423_elements(49)); -- 
    -- CP-element group 50:  transition  input  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	92 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (11) 
      -- CP-element group 50: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/addr_of_2650_request/$entry
      -- CP-element group 50: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/addr_of_2650_request/req
      -- CP-element group 50: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/addr_of_2650_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/array_obj_ref_2649_root_address_calculated
      -- CP-element group 50: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/array_obj_ref_2649_offset_calculated
      -- CP-element group 50: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/array_obj_ref_2649_final_index_sum_regn_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/array_obj_ref_2649_final_index_sum_regn_Update/ack
      -- CP-element group 50: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/array_obj_ref_2649_base_plus_offset/$entry
      -- CP-element group 50: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/array_obj_ref_2649_base_plus_offset/$exit
      -- CP-element group 50: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/array_obj_ref_2649_base_plus_offset/sum_rename_req
      -- CP-element group 50: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/array_obj_ref_2649_base_plus_offset/sum_rename_ack
      -- 
    ack_7222_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2649_index_offset_ack_1, ack => convTransposeC_CP_6423_elements(50)); -- 
    req_7231_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7231_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(50), ack => addr_of_2650_final_reg_req_0); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/addr_of_2650_request/$exit
      -- CP-element group 51: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/addr_of_2650_request/ack
      -- CP-element group 51: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/addr_of_2650_sample_completed_
      -- 
    ack_7232_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2650_final_reg_ack_0, ack => convTransposeC_CP_6423_elements(51)); -- 
    -- CP-element group 52:  fork  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	92 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	53 
    -- CP-element group 52:  members (19) 
      -- CP-element group 52: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2653_base_plus_offset/$entry
      -- CP-element group 52: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2653_base_address_resized
      -- CP-element group 52: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2653_base_addr_resize/$exit
      -- CP-element group 52: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2653_word_addrgen/root_register_ack
      -- CP-element group 52: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/addr_of_2650_complete/ack
      -- CP-element group 52: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/addr_of_2650_complete/$exit
      -- CP-element group 52: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2653_base_addr_resize/$entry
      -- CP-element group 52: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2653_base_addr_resize/base_resize_req
      -- CP-element group 52: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2653_word_addrgen/root_register_req
      -- CP-element group 52: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2653_base_addr_resize/base_resize_ack
      -- CP-element group 52: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2653_base_plus_offset/$exit
      -- CP-element group 52: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2653_base_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2653_word_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2653_base_plus_offset/sum_rename_req
      -- CP-element group 52: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2653_root_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2653_word_addrgen/$exit
      -- CP-element group 52: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2653_word_addrgen/$entry
      -- CP-element group 52: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2653_base_plus_offset/sum_rename_ack
      -- CP-element group 52: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/addr_of_2650_update_completed_
      -- 
    ack_7237_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2650_final_reg_ack_1, ack => convTransposeC_CP_6423_elements(52)); -- 
    -- CP-element group 53:  join  transition  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	46 
    -- CP-element group 53: 	52 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (9) 
      -- CP-element group 53: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2653_Sample/ptr_deref_2653_Split/split_req
      -- CP-element group 53: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2653_Sample/ptr_deref_2653_Split/split_ack
      -- CP-element group 53: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2653_Sample/ptr_deref_2653_Split/$exit
      -- CP-element group 53: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2653_Sample/word_access_start/$entry
      -- CP-element group 53: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2653_Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2653_Sample/ptr_deref_2653_Split/$entry
      -- CP-element group 53: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2653_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2653_Sample/word_access_start/word_0/rr
      -- CP-element group 53: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2653_Sample/word_access_start/word_0/$entry
      -- 
    rr_7275_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7275_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(53), ack => ptr_deref_2653_store_0_req_0); -- 
    convTransposeC_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_6423_elements(46) & convTransposeC_CP_6423_elements(52);
      gj_convTransposeC_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6423_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (5) 
      -- CP-element group 54: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2653_Sample/word_access_start/$exit
      -- CP-element group 54: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2653_Sample/word_access_start/word_0/ra
      -- CP-element group 54: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2653_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2653_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2653_Sample/word_access_start/word_0/$exit
      -- 
    ra_7276_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2653_store_0_ack_0, ack => convTransposeC_CP_6423_elements(54)); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	92 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	58 
    -- CP-element group 55:  members (5) 
      -- CP-element group 55: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2653_Update/word_access_complete/$exit
      -- CP-element group 55: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2653_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2653_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2653_Update/word_access_complete/word_0/ca
      -- CP-element group 55: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2653_Update/word_access_complete/word_0/$exit
      -- 
    ca_7287_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2653_store_0_ack_1, ack => convTransposeC_CP_6423_elements(55)); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	92 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/type_cast_2659_Sample/ra
      -- CP-element group 56: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/type_cast_2659_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/type_cast_2659_sample_completed_
      -- 
    ra_7296_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2659_inst_ack_0, ack => convTransposeC_CP_6423_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	92 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/type_cast_2659_Update/ca
      -- CP-element group 57: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/type_cast_2659_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/type_cast_2659_update_completed_
      -- 
    ca_7301_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2659_inst_ack_1, ack => convTransposeC_CP_6423_elements(57)); -- 
    -- CP-element group 58:  branch  join  transition  place  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	41 
    -- CP-element group 58: 	49 
    -- CP-element group 58: 	55 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58: 	60 
    -- CP-element group 58:  members (10) 
      -- CP-element group 58: 	 branch_block_stmt_2296/if_stmt_2672_eval_test/$entry
      -- CP-element group 58: 	 branch_block_stmt_2296/if_stmt_2672_dead_link/$entry
      -- CP-element group 58: 	 branch_block_stmt_2296/if_stmt_2672__entry__
      -- CP-element group 58: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671__exit__
      -- CP-element group 58: 	 branch_block_stmt_2296/if_stmt_2672_eval_test/$exit
      -- CP-element group 58: 	 branch_block_stmt_2296/if_stmt_2672_eval_test/branch_req
      -- CP-element group 58: 	 branch_block_stmt_2296/if_stmt_2672_if_link/$entry
      -- CP-element group 58: 	 branch_block_stmt_2296/if_stmt_2672_else_link/$entry
      -- CP-element group 58: 	 branch_block_stmt_2296/R_cmp_2673_place
      -- CP-element group 58: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/$exit
      -- 
    branch_req_7309_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_7309_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(58), ack => if_stmt_2672_branch_req_0); -- 
    convTransposeC_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_6423_elements(41) & convTransposeC_CP_6423_elements(49) & convTransposeC_CP_6423_elements(55) & convTransposeC_CP_6423_elements(57);
      gj_convTransposeC_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6423_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	87 
    -- CP-element group 59: 	88 
    -- CP-element group 59:  members (24) 
      -- CP-element group 59: 	 branch_block_stmt_2296/merge_stmt_2678_PhiReqMerge
      -- CP-element group 59: 	 branch_block_stmt_2296/whilex_xbody_ifx_xthen
      -- CP-element group 59: 	 branch_block_stmt_2296/assign_stmt_2684/$exit
      -- CP-element group 59: 	 branch_block_stmt_2296/merge_stmt_2678__exit__
      -- CP-element group 59: 	 branch_block_stmt_2296/ifx_xthen_whilex_xbody
      -- CP-element group 59: 	 branch_block_stmt_2296/assign_stmt_2684__exit__
      -- CP-element group 59: 	 branch_block_stmt_2296/assign_stmt_2684__entry__
      -- CP-element group 59: 	 branch_block_stmt_2296/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2566/phi_stmt_2566_sources/$entry
      -- CP-element group 59: 	 branch_block_stmt_2296/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2566/$entry
      -- CP-element group 59: 	 branch_block_stmt_2296/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2566/phi_stmt_2566_sources/type_cast_2572/SplitProtocol/Sample/rr
      -- CP-element group 59: 	 branch_block_stmt_2296/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2566/phi_stmt_2566_sources/type_cast_2572/$entry
      -- CP-element group 59: 	 branch_block_stmt_2296/if_stmt_2672_if_link/$exit
      -- CP-element group 59: 	 branch_block_stmt_2296/if_stmt_2672_if_link/if_choice_transition
      -- CP-element group 59: 	 branch_block_stmt_2296/assign_stmt_2684/$entry
      -- CP-element group 59: 	 branch_block_stmt_2296/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2566/phi_stmt_2566_sources/type_cast_2572/SplitProtocol/Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_2296/ifx_xthen_whilex_xbody_PhiReq/$entry
      -- CP-element group 59: 	 branch_block_stmt_2296/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2566/phi_stmt_2566_sources/type_cast_2572/SplitProtocol/Update/$entry
      -- CP-element group 59: 	 branch_block_stmt_2296/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2566/phi_stmt_2566_sources/type_cast_2572/SplitProtocol/$entry
      -- CP-element group 59: 	 branch_block_stmt_2296/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2566/phi_stmt_2566_sources/type_cast_2572/SplitProtocol/Update/cr
      -- CP-element group 59: 	 branch_block_stmt_2296/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 59: 	 branch_block_stmt_2296/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 59: 	 branch_block_stmt_2296/merge_stmt_2678_PhiAck/$entry
      -- CP-element group 59: 	 branch_block_stmt_2296/merge_stmt_2678_PhiAck/$exit
      -- CP-element group 59: 	 branch_block_stmt_2296/merge_stmt_2678_PhiAck/dummy
      -- 
    if_choice_transition_7314_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2672_branch_ack_1, ack => convTransposeC_CP_6423_elements(59)); -- 
    rr_7512_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7512_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(59), ack => type_cast_2572_inst_req_0); -- 
    cr_7517_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7517_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(59), ack => type_cast_2572_inst_req_1); -- 
    -- CP-element group 60:  fork  transition  place  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	58 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60: 	62 
    -- CP-element group 60: 	64 
    -- CP-element group 60: 	66 
    -- CP-element group 60:  members (24) 
      -- CP-element group 60: 	 branch_block_stmt_2296/whilex_xbody_ifx_xelse
      -- CP-element group 60: 	 branch_block_stmt_2296/assign_stmt_2692_to_assign_stmt_2728/type_cast_2696_update_start_
      -- CP-element group 60: 	 branch_block_stmt_2296/assign_stmt_2692_to_assign_stmt_2728/type_cast_2696_Update/cr
      -- CP-element group 60: 	 branch_block_stmt_2296/assign_stmt_2692_to_assign_stmt_2728/type_cast_2722_update_start_
      -- CP-element group 60: 	 branch_block_stmt_2296/merge_stmt_2686_PhiReqMerge
      -- CP-element group 60: 	 branch_block_stmt_2296/assign_stmt_2692_to_assign_stmt_2728/type_cast_2722_Update/$entry
      -- CP-element group 60: 	 branch_block_stmt_2296/assign_stmt_2692_to_assign_stmt_2728/type_cast_2696_Update/$entry
      -- CP-element group 60: 	 branch_block_stmt_2296/assign_stmt_2692_to_assign_stmt_2728/type_cast_2696_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_2296/assign_stmt_2692_to_assign_stmt_2728/$entry
      -- CP-element group 60: 	 branch_block_stmt_2296/merge_stmt_2686__exit__
      -- CP-element group 60: 	 branch_block_stmt_2296/assign_stmt_2692_to_assign_stmt_2728__entry__
      -- CP-element group 60: 	 branch_block_stmt_2296/assign_stmt_2692_to_assign_stmt_2728/type_cast_2696_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_2296/if_stmt_2672_else_link/$exit
      -- CP-element group 60: 	 branch_block_stmt_2296/if_stmt_2672_else_link/else_choice_transition
      -- CP-element group 60: 	 branch_block_stmt_2296/assign_stmt_2692_to_assign_stmt_2728/type_cast_2705_update_start_
      -- CP-element group 60: 	 branch_block_stmt_2296/merge_stmt_2686_PhiAck/$entry
      -- CP-element group 60: 	 branch_block_stmt_2296/merge_stmt_2686_PhiAck/$exit
      -- CP-element group 60: 	 branch_block_stmt_2296/merge_stmt_2686_PhiAck/dummy
      -- CP-element group 60: 	 branch_block_stmt_2296/assign_stmt_2692_to_assign_stmt_2728/type_cast_2722_Update/cr
      -- CP-element group 60: 	 branch_block_stmt_2296/assign_stmt_2692_to_assign_stmt_2728/type_cast_2705_Update/$entry
      -- CP-element group 60: 	 branch_block_stmt_2296/assign_stmt_2692_to_assign_stmt_2728/type_cast_2705_Update/cr
      -- CP-element group 60: 	 branch_block_stmt_2296/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 60: 	 branch_block_stmt_2296/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 60: 	 branch_block_stmt_2296/assign_stmt_2692_to_assign_stmt_2728/type_cast_2696_Sample/rr
      -- 
    else_choice_transition_7318_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2672_branch_ack_0, ack => convTransposeC_CP_6423_elements(60)); -- 
    cr_7339_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7339_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(60), ack => type_cast_2696_inst_req_1); -- 
    cr_7367_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7367_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(60), ack => type_cast_2722_inst_req_1); -- 
    cr_7353_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7353_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(60), ack => type_cast_2705_inst_req_1); -- 
    rr_7334_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7334_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(60), ack => type_cast_2696_inst_req_0); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_2296/assign_stmt_2692_to_assign_stmt_2728/type_cast_2696_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_2296/assign_stmt_2692_to_assign_stmt_2728/type_cast_2696_Sample/ra
      -- CP-element group 61: 	 branch_block_stmt_2296/assign_stmt_2692_to_assign_stmt_2728/type_cast_2696_Sample/$exit
      -- 
    ra_7335_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2696_inst_ack_0, ack => convTransposeC_CP_6423_elements(61)); -- 
    -- CP-element group 62:  transition  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	60 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (6) 
      -- CP-element group 62: 	 branch_block_stmt_2296/assign_stmt_2692_to_assign_stmt_2728/type_cast_2696_Update/ca
      -- CP-element group 62: 	 branch_block_stmt_2296/assign_stmt_2692_to_assign_stmt_2728/type_cast_2705_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_2296/assign_stmt_2692_to_assign_stmt_2728/type_cast_2696_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_2296/assign_stmt_2692_to_assign_stmt_2728/type_cast_2696_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_2296/assign_stmt_2692_to_assign_stmt_2728/type_cast_2705_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_2296/assign_stmt_2692_to_assign_stmt_2728/type_cast_2705_Sample/rr
      -- 
    ca_7340_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2696_inst_ack_1, ack => convTransposeC_CP_6423_elements(62)); -- 
    rr_7348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(62), ack => type_cast_2705_inst_req_0); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_2296/assign_stmt_2692_to_assign_stmt_2728/type_cast_2705_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_2296/assign_stmt_2692_to_assign_stmt_2728/type_cast_2705_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_2296/assign_stmt_2692_to_assign_stmt_2728/type_cast_2705_Sample/ra
      -- 
    ra_7349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2705_inst_ack_0, ack => convTransposeC_CP_6423_elements(63)); -- 
    -- CP-element group 64:  transition  input  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	60 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64:  members (6) 
      -- CP-element group 64: 	 branch_block_stmt_2296/assign_stmt_2692_to_assign_stmt_2728/type_cast_2722_Sample/rr
      -- CP-element group 64: 	 branch_block_stmt_2296/assign_stmt_2692_to_assign_stmt_2728/type_cast_2722_Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_2296/assign_stmt_2692_to_assign_stmt_2728/type_cast_2705_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_2296/assign_stmt_2692_to_assign_stmt_2728/type_cast_2705_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_2296/assign_stmt_2692_to_assign_stmt_2728/type_cast_2705_Update/ca
      -- CP-element group 64: 	 branch_block_stmt_2296/assign_stmt_2692_to_assign_stmt_2728/type_cast_2722_sample_start_
      -- 
    ca_7354_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2705_inst_ack_1, ack => convTransposeC_CP_6423_elements(64)); -- 
    rr_7362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(64), ack => type_cast_2722_inst_req_0); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_2296/assign_stmt_2692_to_assign_stmt_2728/type_cast_2722_Sample/$exit
      -- CP-element group 65: 	 branch_block_stmt_2296/assign_stmt_2692_to_assign_stmt_2728/type_cast_2722_Sample/ra
      -- CP-element group 65: 	 branch_block_stmt_2296/assign_stmt_2692_to_assign_stmt_2728/type_cast_2722_sample_completed_
      -- 
    ra_7363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2722_inst_ack_0, ack => convTransposeC_CP_6423_elements(65)); -- 
    -- CP-element group 66:  branch  transition  place  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	60 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66: 	68 
    -- CP-element group 66:  members (13) 
      -- CP-element group 66: 	 branch_block_stmt_2296/if_stmt_2729_eval_test/$exit
      -- CP-element group 66: 	 branch_block_stmt_2296/R_cmp87_2730_place
      -- CP-element group 66: 	 branch_block_stmt_2296/if_stmt_2729_eval_test/$entry
      -- CP-element group 66: 	 branch_block_stmt_2296/assign_stmt_2692_to_assign_stmt_2728/$exit
      -- CP-element group 66: 	 branch_block_stmt_2296/assign_stmt_2692_to_assign_stmt_2728/type_cast_2722_Update/ca
      -- CP-element group 66: 	 branch_block_stmt_2296/if_stmt_2729_dead_link/$entry
      -- CP-element group 66: 	 branch_block_stmt_2296/assign_stmt_2692_to_assign_stmt_2728/type_cast_2722_update_completed_
      -- CP-element group 66: 	 branch_block_stmt_2296/assign_stmt_2692_to_assign_stmt_2728__exit__
      -- CP-element group 66: 	 branch_block_stmt_2296/if_stmt_2729__entry__
      -- CP-element group 66: 	 branch_block_stmt_2296/assign_stmt_2692_to_assign_stmt_2728/type_cast_2722_Update/$exit
      -- CP-element group 66: 	 branch_block_stmt_2296/if_stmt_2729_eval_test/branch_req
      -- CP-element group 66: 	 branch_block_stmt_2296/if_stmt_2729_if_link/$entry
      -- CP-element group 66: 	 branch_block_stmt_2296/if_stmt_2729_else_link/$entry
      -- 
    ca_7368_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2722_inst_ack_1, ack => convTransposeC_CP_6423_elements(66)); -- 
    branch_req_7376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_7376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(66), ack => if_stmt_2729_branch_req_0); -- 
    -- CP-element group 67:  merge  transition  place  input  output  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67:  members (15) 
      -- CP-element group 67: 	 branch_block_stmt_2296/assign_stmt_2739/$entry
      -- CP-element group 67: 	 branch_block_stmt_2296/ifx_xelse_whilex_xend
      -- CP-element group 67: 	 branch_block_stmt_2296/assign_stmt_2739/WPIPE_Block2_done_2737_Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_2296/merge_stmt_2735_PhiReqMerge
      -- CP-element group 67: 	 branch_block_stmt_2296/assign_stmt_2739/WPIPE_Block2_done_2737_sample_start_
      -- CP-element group 67: 	 branch_block_stmt_2296/assign_stmt_2739__entry__
      -- CP-element group 67: 	 branch_block_stmt_2296/merge_stmt_2735__exit__
      -- CP-element group 67: 	 branch_block_stmt_2296/if_stmt_2729_if_link/$exit
      -- CP-element group 67: 	 branch_block_stmt_2296/if_stmt_2729_if_link/if_choice_transition
      -- CP-element group 67: 	 branch_block_stmt_2296/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 67: 	 branch_block_stmt_2296/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 67: 	 branch_block_stmt_2296/merge_stmt_2735_PhiAck/$entry
      -- CP-element group 67: 	 branch_block_stmt_2296/merge_stmt_2735_PhiAck/$exit
      -- CP-element group 67: 	 branch_block_stmt_2296/merge_stmt_2735_PhiAck/dummy
      -- CP-element group 67: 	 branch_block_stmt_2296/assign_stmt_2739/WPIPE_Block2_done_2737_Sample/req
      -- 
    if_choice_transition_7381_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2729_branch_ack_1, ack => convTransposeC_CP_6423_elements(67)); -- 
    req_7398_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7398_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(67), ack => WPIPE_Block2_done_2737_inst_req_0); -- 
    -- CP-element group 68:  fork  transition  place  input  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	80 
    -- CP-element group 68: 	79 
    -- CP-element group 68: 	76 
    -- CP-element group 68: 	77 
    -- CP-element group 68:  members (20) 
      -- CP-element group 68: 	 branch_block_stmt_2296/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2438/$entry
      -- CP-element group 68: 	 branch_block_stmt_2296/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2438/phi_stmt_2438_sources/type_cast_2441/SplitProtocol/$entry
      -- CP-element group 68: 	 branch_block_stmt_2296/ifx_xelse_whilex_xbodyx_xouter
      -- CP-element group 68: 	 branch_block_stmt_2296/if_stmt_2729_else_link/else_choice_transition
      -- CP-element group 68: 	 branch_block_stmt_2296/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2438/phi_stmt_2438_sources/type_cast_2441/$entry
      -- CP-element group 68: 	 branch_block_stmt_2296/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2445/$entry
      -- CP-element group 68: 	 branch_block_stmt_2296/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2445/phi_stmt_2445_sources/type_cast_2448/SplitProtocol/Sample/rr
      -- CP-element group 68: 	 branch_block_stmt_2296/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2445/phi_stmt_2445_sources/$entry
      -- CP-element group 68: 	 branch_block_stmt_2296/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2438/phi_stmt_2438_sources/type_cast_2441/SplitProtocol/Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_2296/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2445/phi_stmt_2445_sources/type_cast_2448/SplitProtocol/Update/cr
      -- CP-element group 68: 	 branch_block_stmt_2296/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2438/phi_stmt_2438_sources/type_cast_2441/SplitProtocol/Update/cr
      -- CP-element group 68: 	 branch_block_stmt_2296/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2445/phi_stmt_2445_sources/type_cast_2448/SplitProtocol/Update/$entry
      -- CP-element group 68: 	 branch_block_stmt_2296/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2445/phi_stmt_2445_sources/type_cast_2448/SplitProtocol/Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_2296/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2438/phi_stmt_2438_sources/$entry
      -- CP-element group 68: 	 branch_block_stmt_2296/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2438/phi_stmt_2438_sources/type_cast_2441/SplitProtocol/Sample/rr
      -- CP-element group 68: 	 branch_block_stmt_2296/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2445/phi_stmt_2445_sources/type_cast_2448/$entry
      -- CP-element group 68: 	 branch_block_stmt_2296/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2438/phi_stmt_2438_sources/type_cast_2441/SplitProtocol/Update/$entry
      -- CP-element group 68: 	 branch_block_stmt_2296/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 68: 	 branch_block_stmt_2296/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2445/phi_stmt_2445_sources/type_cast_2448/SplitProtocol/$entry
      -- CP-element group 68: 	 branch_block_stmt_2296/if_stmt_2729_else_link/$exit
      -- 
    else_choice_transition_7385_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2729_branch_ack_0, ack => convTransposeC_CP_6423_elements(68)); -- 
    rr_7480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(68), ack => type_cast_2448_inst_req_0); -- 
    cr_7485_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7485_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(68), ack => type_cast_2448_inst_req_1); -- 
    cr_7462_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7462_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(68), ack => type_cast_2441_inst_req_1); -- 
    rr_7457_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7457_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(68), ack => type_cast_2441_inst_req_0); -- 
    -- CP-element group 69:  transition  input  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	67 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69:  members (6) 
      -- CP-element group 69: 	 branch_block_stmt_2296/assign_stmt_2739/WPIPE_Block2_done_2737_update_start_
      -- CP-element group 69: 	 branch_block_stmt_2296/assign_stmt_2739/WPIPE_Block2_done_2737_Update/req
      -- CP-element group 69: 	 branch_block_stmt_2296/assign_stmt_2739/WPIPE_Block2_done_2737_sample_completed_
      -- CP-element group 69: 	 branch_block_stmt_2296/assign_stmt_2739/WPIPE_Block2_done_2737_Sample/$exit
      -- CP-element group 69: 	 branch_block_stmt_2296/assign_stmt_2739/WPIPE_Block2_done_2737_Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_2296/assign_stmt_2739/WPIPE_Block2_done_2737_Sample/ack
      -- 
    ack_7399_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_done_2737_inst_ack_0, ack => convTransposeC_CP_6423_elements(69)); -- 
    req_7403_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7403_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(69), ack => WPIPE_Block2_done_2737_inst_req_1); -- 
    -- CP-element group 70:  transition  place  input  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (16) 
      -- CP-element group 70: 	 branch_block_stmt_2296/assign_stmt_2739/$exit
      -- CP-element group 70: 	 branch_block_stmt_2296/assign_stmt_2739/WPIPE_Block2_done_2737_update_completed_
      -- CP-element group 70: 	 branch_block_stmt_2296/assign_stmt_2739/WPIPE_Block2_done_2737_Update/ack
      -- CP-element group 70: 	 branch_block_stmt_2296/assign_stmt_2739/WPIPE_Block2_done_2737_Update/$exit
      -- CP-element group 70: 	 branch_block_stmt_2296/merge_stmt_2741_PhiReqMerge
      -- CP-element group 70: 	 branch_block_stmt_2296/return___PhiReq/$entry
      -- CP-element group 70: 	 $exit
      -- CP-element group 70: 	 branch_block_stmt_2296/$exit
      -- CP-element group 70: 	 branch_block_stmt_2296/branch_block_stmt_2296__exit__
      -- CP-element group 70: 	 branch_block_stmt_2296/assign_stmt_2739__exit__
      -- CP-element group 70: 	 branch_block_stmt_2296/return__
      -- CP-element group 70: 	 branch_block_stmt_2296/merge_stmt_2741__exit__
      -- CP-element group 70: 	 branch_block_stmt_2296/return___PhiReq/$exit
      -- CP-element group 70: 	 branch_block_stmt_2296/merge_stmt_2741_PhiAck/$entry
      -- CP-element group 70: 	 branch_block_stmt_2296/merge_stmt_2741_PhiAck/$exit
      -- CP-element group 70: 	 branch_block_stmt_2296/merge_stmt_2741_PhiAck/dummy
      -- 
    ack_7404_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_done_2737_inst_ack_1, ack => convTransposeC_CP_6423_elements(70)); -- 
    -- CP-element group 71:  transition  output  delay-element  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	31 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	75 
    -- CP-element group 71:  members (4) 
      -- CP-element group 71: 	 branch_block_stmt_2296/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2438/phi_stmt_2438_sources/type_cast_2444_konst_delay_trans
      -- CP-element group 71: 	 branch_block_stmt_2296/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2438/phi_stmt_2438_sources/$exit
      -- CP-element group 71: 	 branch_block_stmt_2296/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2438/$exit
      -- CP-element group 71: 	 branch_block_stmt_2296/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2438/phi_stmt_2438_req
      -- 
    phi_stmt_2438_req_7415_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2438_req_7415_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(71), ack => phi_stmt_2438_req_1); -- 
    -- Element group convTransposeC_CP_6423_elements(71) is a control-delay.
    cp_element_71_delay: control_delay_element  generic map(name => " 71_delay", delay_value => 1)  port map(req => convTransposeC_CP_6423_elements(31), ack => convTransposeC_CP_6423_elements(71), clk => clk, reset =>reset);
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	31 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	74 
    -- CP-element group 72:  members (2) 
      -- CP-element group 72: 	 branch_block_stmt_2296/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2445/phi_stmt_2445_sources/type_cast_2450/SplitProtocol/Sample/$exit
      -- CP-element group 72: 	 branch_block_stmt_2296/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2445/phi_stmt_2445_sources/type_cast_2450/SplitProtocol/Sample/ra
      -- 
    ra_7432_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2450_inst_ack_0, ack => convTransposeC_CP_6423_elements(72)); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	31 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (2) 
      -- CP-element group 73: 	 branch_block_stmt_2296/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2445/phi_stmt_2445_sources/type_cast_2450/SplitProtocol/Update/$exit
      -- CP-element group 73: 	 branch_block_stmt_2296/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2445/phi_stmt_2445_sources/type_cast_2450/SplitProtocol/Update/ca
      -- 
    ca_7437_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2450_inst_ack_1, ack => convTransposeC_CP_6423_elements(73)); -- 
    -- CP-element group 74:  join  transition  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	72 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74:  members (5) 
      -- CP-element group 74: 	 branch_block_stmt_2296/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2445/phi_stmt_2445_sources/type_cast_2450/SplitProtocol/$exit
      -- CP-element group 74: 	 branch_block_stmt_2296/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2445/$exit
      -- CP-element group 74: 	 branch_block_stmt_2296/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2445/phi_stmt_2445_sources/$exit
      -- CP-element group 74: 	 branch_block_stmt_2296/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2445/phi_stmt_2445_req
      -- CP-element group 74: 	 branch_block_stmt_2296/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2445/phi_stmt_2445_sources/type_cast_2450/$exit
      -- 
    phi_stmt_2445_req_7438_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2445_req_7438_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(74), ack => phi_stmt_2445_req_1); -- 
    convTransposeC_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_6423_elements(72) & convTransposeC_CP_6423_elements(73);
      gj_convTransposeC_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6423_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  join  transition  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	71 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	83 
    -- CP-element group 75:  members (1) 
      -- CP-element group 75: 	 branch_block_stmt_2296/entry_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeC_cp_element_group_75: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_75"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_6423_elements(71) & convTransposeC_CP_6423_elements(74);
      gj_convTransposeC_cp_element_group_75 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6423_elements(75), clk => clk, reset => reset); --
    end block;
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	68 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	78 
    -- CP-element group 76:  members (2) 
      -- CP-element group 76: 	 branch_block_stmt_2296/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2438/phi_stmt_2438_sources/type_cast_2441/SplitProtocol/Sample/ra
      -- CP-element group 76: 	 branch_block_stmt_2296/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2438/phi_stmt_2438_sources/type_cast_2441/SplitProtocol/Sample/$exit
      -- 
    ra_7458_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2441_inst_ack_0, ack => convTransposeC_CP_6423_elements(76)); -- 
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	68 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (2) 
      -- CP-element group 77: 	 branch_block_stmt_2296/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2438/phi_stmt_2438_sources/type_cast_2441/SplitProtocol/Update/$exit
      -- CP-element group 77: 	 branch_block_stmt_2296/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2438/phi_stmt_2438_sources/type_cast_2441/SplitProtocol/Update/ca
      -- 
    ca_7463_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2441_inst_ack_1, ack => convTransposeC_CP_6423_elements(77)); -- 
    -- CP-element group 78:  join  transition  output  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	76 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	82 
    -- CP-element group 78:  members (5) 
      -- CP-element group 78: 	 branch_block_stmt_2296/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2438/$exit
      -- CP-element group 78: 	 branch_block_stmt_2296/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2438/phi_stmt_2438_sources/type_cast_2441/SplitProtocol/$exit
      -- CP-element group 78: 	 branch_block_stmt_2296/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2438/phi_stmt_2438_sources/type_cast_2441/$exit
      -- CP-element group 78: 	 branch_block_stmt_2296/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2438/phi_stmt_2438_sources/$exit
      -- CP-element group 78: 	 branch_block_stmt_2296/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2438/phi_stmt_2438_req
      -- 
    phi_stmt_2438_req_7464_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2438_req_7464_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(78), ack => phi_stmt_2438_req_0); -- 
    convTransposeC_cp_element_group_78: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_78"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_6423_elements(76) & convTransposeC_CP_6423_elements(77);
      gj_convTransposeC_cp_element_group_78 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6423_elements(78), clk => clk, reset => reset); --
    end block;
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	68 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	81 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_2296/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2445/phi_stmt_2445_sources/type_cast_2448/SplitProtocol/Sample/ra
      -- CP-element group 79: 	 branch_block_stmt_2296/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2445/phi_stmt_2445_sources/type_cast_2448/SplitProtocol/Sample/$exit
      -- 
    ra_7481_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2448_inst_ack_0, ack => convTransposeC_CP_6423_elements(79)); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	68 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (2) 
      -- CP-element group 80: 	 branch_block_stmt_2296/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2445/phi_stmt_2445_sources/type_cast_2448/SplitProtocol/Update/ca
      -- CP-element group 80: 	 branch_block_stmt_2296/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2445/phi_stmt_2445_sources/type_cast_2448/SplitProtocol/Update/$exit
      -- 
    ca_7486_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2448_inst_ack_1, ack => convTransposeC_CP_6423_elements(80)); -- 
    -- CP-element group 81:  join  transition  output  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	80 
    -- CP-element group 81: 	79 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	82 
    -- CP-element group 81:  members (5) 
      -- CP-element group 81: 	 branch_block_stmt_2296/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2445/phi_stmt_2445_req
      -- CP-element group 81: 	 branch_block_stmt_2296/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2445/$exit
      -- CP-element group 81: 	 branch_block_stmt_2296/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2445/phi_stmt_2445_sources/type_cast_2448/SplitProtocol/$exit
      -- CP-element group 81: 	 branch_block_stmt_2296/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2445/phi_stmt_2445_sources/$exit
      -- CP-element group 81: 	 branch_block_stmt_2296/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2445/phi_stmt_2445_sources/type_cast_2448/$exit
      -- 
    phi_stmt_2445_req_7487_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2445_req_7487_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(81), ack => phi_stmt_2445_req_0); -- 
    convTransposeC_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_6423_elements(80) & convTransposeC_CP_6423_elements(79);
      gj_convTransposeC_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6423_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  join  transition  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	81 
    -- CP-element group 82: 	78 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (1) 
      -- CP-element group 82: 	 branch_block_stmt_2296/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeC_cp_element_group_82: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_82"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_6423_elements(81) & convTransposeC_CP_6423_elements(78);
      gj_convTransposeC_cp_element_group_82 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6423_elements(82), clk => clk, reset => reset); --
    end block;
    -- CP-element group 83:  merge  fork  transition  place  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	82 
    -- CP-element group 83: 	75 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83: 	85 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_2296/merge_stmt_2437_PhiReqMerge
      -- CP-element group 83: 	 branch_block_stmt_2296/merge_stmt_2437_PhiAck/$entry
      -- 
    convTransposeC_CP_6423_elements(83) <= OrReduce(convTransposeC_CP_6423_elements(82) & convTransposeC_CP_6423_elements(75));
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (1) 
      -- CP-element group 84: 	 branch_block_stmt_2296/merge_stmt_2437_PhiAck/phi_stmt_2438_ack
      -- 
    phi_stmt_2438_ack_7492_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2438_ack_0, ack => convTransposeC_CP_6423_elements(84)); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	83 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85:  members (1) 
      -- CP-element group 85: 	 branch_block_stmt_2296/merge_stmt_2437_PhiAck/phi_stmt_2445_ack
      -- 
    phi_stmt_2445_ack_7493_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2445_ack_0, ack => convTransposeC_CP_6423_elements(85)); -- 
    -- CP-element group 86:  join  fork  transition  place  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	32 
    -- CP-element group 86: 	33 
    -- CP-element group 86: 	34 
    -- CP-element group 86: 	35 
    -- CP-element group 86:  members (16) 
      -- CP-element group 86: 	 branch_block_stmt_2296/merge_stmt_2437_PhiAck/$exit
      -- CP-element group 86: 	 branch_block_stmt_2296/merge_stmt_2437__exit__
      -- CP-element group 86: 	 branch_block_stmt_2296/assign_stmt_2456_to_assign_stmt_2563__entry__
      -- CP-element group 86: 	 branch_block_stmt_2296/assign_stmt_2456_to_assign_stmt_2563/$entry
      -- CP-element group 86: 	 branch_block_stmt_2296/assign_stmt_2456_to_assign_stmt_2563/type_cast_2455_sample_start_
      -- CP-element group 86: 	 branch_block_stmt_2296/assign_stmt_2456_to_assign_stmt_2563/type_cast_2455_update_start_
      -- CP-element group 86: 	 branch_block_stmt_2296/assign_stmt_2456_to_assign_stmt_2563/type_cast_2455_Sample/$entry
      -- CP-element group 86: 	 branch_block_stmt_2296/assign_stmt_2456_to_assign_stmt_2563/type_cast_2455_Sample/rr
      -- CP-element group 86: 	 branch_block_stmt_2296/assign_stmt_2456_to_assign_stmt_2563/type_cast_2455_Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_2296/assign_stmt_2456_to_assign_stmt_2563/type_cast_2455_Update/cr
      -- CP-element group 86: 	 branch_block_stmt_2296/assign_stmt_2456_to_assign_stmt_2563/type_cast_2460_sample_start_
      -- CP-element group 86: 	 branch_block_stmt_2296/assign_stmt_2456_to_assign_stmt_2563/type_cast_2460_update_start_
      -- CP-element group 86: 	 branch_block_stmt_2296/assign_stmt_2456_to_assign_stmt_2563/type_cast_2460_Sample/$entry
      -- CP-element group 86: 	 branch_block_stmt_2296/assign_stmt_2456_to_assign_stmt_2563/type_cast_2460_Sample/rr
      -- CP-element group 86: 	 branch_block_stmt_2296/assign_stmt_2456_to_assign_stmt_2563/type_cast_2460_Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_2296/assign_stmt_2456_to_assign_stmt_2563/type_cast_2460_Update/cr
      -- 
    rr_7030_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7030_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(86), ack => type_cast_2455_inst_req_0); -- 
    cr_7035_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7035_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(86), ack => type_cast_2455_inst_req_1); -- 
    rr_7044_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7044_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(86), ack => type_cast_2460_inst_req_0); -- 
    cr_7049_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7049_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(86), ack => type_cast_2460_inst_req_1); -- 
    convTransposeC_cp_element_group_86: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_86"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_6423_elements(84) & convTransposeC_CP_6423_elements(85);
      gj_convTransposeC_cp_element_group_86 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6423_elements(86), clk => clk, reset => reset); --
    end block;
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	59 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	89 
    -- CP-element group 87:  members (2) 
      -- CP-element group 87: 	 branch_block_stmt_2296/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2566/phi_stmt_2566_sources/type_cast_2572/SplitProtocol/Sample/$exit
      -- CP-element group 87: 	 branch_block_stmt_2296/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2566/phi_stmt_2566_sources/type_cast_2572/SplitProtocol/Sample/ra
      -- 
    ra_7513_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2572_inst_ack_0, ack => convTransposeC_CP_6423_elements(87)); -- 
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	59 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	89 
    -- CP-element group 88:  members (2) 
      -- CP-element group 88: 	 branch_block_stmt_2296/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2566/phi_stmt_2566_sources/type_cast_2572/SplitProtocol/Update/ca
      -- CP-element group 88: 	 branch_block_stmt_2296/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2566/phi_stmt_2566_sources/type_cast_2572/SplitProtocol/Update/$exit
      -- 
    ca_7518_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2572_inst_ack_1, ack => convTransposeC_CP_6423_elements(88)); -- 
    -- CP-element group 89:  join  transition  output  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	87 
    -- CP-element group 89: 	88 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (6) 
      -- CP-element group 89: 	 branch_block_stmt_2296/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2566/phi_stmt_2566_sources/$exit
      -- CP-element group 89: 	 branch_block_stmt_2296/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2566/$exit
      -- CP-element group 89: 	 branch_block_stmt_2296/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2566/phi_stmt_2566_sources/type_cast_2572/$exit
      -- CP-element group 89: 	 branch_block_stmt_2296/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2566/phi_stmt_2566_sources/type_cast_2572/SplitProtocol/$exit
      -- CP-element group 89: 	 branch_block_stmt_2296/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2566/phi_stmt_2566_req
      -- CP-element group 89: 	 branch_block_stmt_2296/ifx_xthen_whilex_xbody_PhiReq/$exit
      -- 
    phi_stmt_2566_req_7519_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2566_req_7519_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(89), ack => phi_stmt_2566_req_1); -- 
    convTransposeC_cp_element_group_89: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_89"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_6423_elements(87) & convTransposeC_CP_6423_elements(88);
      gj_convTransposeC_cp_element_group_89 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6423_elements(89), clk => clk, reset => reset); --
    end block;
    -- CP-element group 90:  transition  output  delay-element  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	36 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (5) 
      -- CP-element group 90: 	 branch_block_stmt_2296/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$exit
      -- CP-element group 90: 	 branch_block_stmt_2296/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2566/phi_stmt_2566_sources/$exit
      -- CP-element group 90: 	 branch_block_stmt_2296/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2566/phi_stmt_2566_sources/type_cast_2570_konst_delay_trans
      -- CP-element group 90: 	 branch_block_stmt_2296/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2566/phi_stmt_2566_req
      -- CP-element group 90: 	 branch_block_stmt_2296/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2566/$exit
      -- 
    phi_stmt_2566_req_7530_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2566_req_7530_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(90), ack => phi_stmt_2566_req_0); -- 
    -- Element group convTransposeC_CP_6423_elements(90) is a control-delay.
    cp_element_90_delay: control_delay_element  generic map(name => " 90_delay", delay_value => 1)  port map(req => convTransposeC_CP_6423_elements(36), ack => convTransposeC_CP_6423_elements(90), clk => clk, reset =>reset);
    -- CP-element group 91:  merge  transition  place  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (2) 
      -- CP-element group 91: 	 branch_block_stmt_2296/merge_stmt_2565_PhiReqMerge
      -- CP-element group 91: 	 branch_block_stmt_2296/merge_stmt_2565_PhiAck/$entry
      -- 
    convTransposeC_CP_6423_elements(91) <= OrReduce(convTransposeC_CP_6423_elements(89) & convTransposeC_CP_6423_elements(90));
    -- CP-element group 92:  fork  transition  place  input  output  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	37 
    -- CP-element group 92: 	40 
    -- CP-element group 92: 	38 
    -- CP-element group 92: 	42 
    -- CP-element group 92: 	48 
    -- CP-element group 92: 	50 
    -- CP-element group 92: 	46 
    -- CP-element group 92: 	52 
    -- CP-element group 92: 	55 
    -- CP-element group 92: 	44 
    -- CP-element group 92: 	56 
    -- CP-element group 92: 	57 
    -- CP-element group 92:  members (45) 
      -- CP-element group 92: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/addr_of_2650_complete/$entry
      -- CP-element group 92: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2653_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/type_cast_2659_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2653_Update/word_access_complete/$entry
      -- CP-element group 92: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/addr_of_2650_complete/req
      -- CP-element group 92: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/type_cast_2659_Update/cr
      -- CP-element group 92: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/type_cast_2659_Sample/rr
      -- CP-element group 92: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2653_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2296/merge_stmt_2565__exit__
      -- CP-element group 92: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671__entry__
      -- CP-element group 92: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2653_Update/word_access_complete/word_0/$entry
      -- CP-element group 92: 	 branch_block_stmt_2296/merge_stmt_2565_PhiAck/$exit
      -- CP-element group 92: 	 branch_block_stmt_2296/merge_stmt_2565_PhiAck/phi_stmt_2566_ack
      -- CP-element group 92: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/type_cast_2659_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/type_cast_2659_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/type_cast_2659_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2653_Update/word_access_complete/word_0/cr
      -- CP-element group 92: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/$entry
      -- CP-element group 92: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/type_cast_2582_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/type_cast_2582_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/type_cast_2582_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/type_cast_2582_Sample/rr
      -- CP-element group 92: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/type_cast_2582_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/type_cast_2582_Update/cr
      -- CP-element group 92: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/type_cast_2612_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/type_cast_2612_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/type_cast_2612_Update/cr
      -- CP-element group 92: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/addr_of_2619_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/array_obj_ref_2618_final_index_sum_regn_update_start
      -- CP-element group 92: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/array_obj_ref_2618_final_index_sum_regn_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/array_obj_ref_2618_final_index_sum_regn_Update/req
      -- CP-element group 92: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/addr_of_2619_complete/$entry
      -- CP-element group 92: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/addr_of_2619_complete/req
      -- CP-element group 92: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2623_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2623_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2623_Update/word_access_complete/$entry
      -- CP-element group 92: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2623_Update/word_access_complete/word_0/$entry
      -- CP-element group 92: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/ptr_deref_2623_Update/word_access_complete/word_0/cr
      -- CP-element group 92: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/type_cast_2643_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/type_cast_2643_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/type_cast_2643_Update/cr
      -- CP-element group 92: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/addr_of_2650_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/array_obj_ref_2649_final_index_sum_regn_update_start
      -- CP-element group 92: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/array_obj_ref_2649_final_index_sum_regn_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2296/assign_stmt_2579_to_assign_stmt_2671/array_obj_ref_2649_final_index_sum_regn_Update/req
      -- 
    phi_stmt_2566_ack_7535_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2566_ack_0, ack => convTransposeC_CP_6423_elements(92)); -- 
    req_7236_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7236_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(92), ack => addr_of_2650_final_reg_req_1); -- 
    cr_7300_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7300_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(92), ack => type_cast_2659_inst_req_1); -- 
    rr_7295_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7295_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(92), ack => type_cast_2659_inst_req_0); -- 
    cr_7286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(92), ack => ptr_deref_2653_store_0_req_1); -- 
    rr_7061_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7061_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(92), ack => type_cast_2582_inst_req_0); -- 
    cr_7066_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7066_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(92), ack => type_cast_2582_inst_req_1); -- 
    cr_7080_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7080_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(92), ack => type_cast_2612_inst_req_1); -- 
    req_7111_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7111_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(92), ack => array_obj_ref_2618_index_offset_req_1); -- 
    req_7126_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7126_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(92), ack => addr_of_2619_final_reg_req_1); -- 
    cr_7171_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7171_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(92), ack => ptr_deref_2623_load_0_req_1); -- 
    cr_7190_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7190_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(92), ack => type_cast_2643_inst_req_1); -- 
    req_7221_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7221_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6423_elements(92), ack => array_obj_ref_2649_index_offset_req_1); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i32_i32_2525_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2546_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2606_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2637_wire : std_logic_vector(31 downto 0);
    signal LOAD_padding_2374_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_padding_2374_word_address_0 : std_logic_vector(0 downto 0);
    signal R_idxprom62_2648_resized : std_logic_vector(13 downto 0);
    signal R_idxprom62_2648_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_2617_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_2617_scaled : std_logic_vector(13 downto 0);
    signal add18_2588 : std_logic_vector(31 downto 0);
    signal add26_2486 : std_logic_vector(31 downto 0);
    signal add37_2501 : std_logic_vector(31 downto 0);
    signal add52_2558 : std_logic_vector(31 downto 0);
    signal add54_2593 : std_logic_vector(31 downto 0);
    signal add67_2666 : std_logic_vector(31 downto 0);
    signal add_2471 : std_logic_vector(31 downto 0);
    signal array_obj_ref_2618_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2618_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2618_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2618_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2618_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2618_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2649_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2649_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2649_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2649_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2649_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2649_root_address : std_logic_vector(13 downto 0);
    signal arrayidx63_2651 : std_logic_vector(31 downto 0);
    signal arrayidx_2620 : std_logic_vector(31 downto 0);
    signal call_2299 : std_logic_vector(15 downto 0);
    signal cmp79_2702 : std_logic_vector(0 downto 0);
    signal cmp87_2728 : std_logic_vector(0 downto 0);
    signal cmp_2671 : std_logic_vector(0 downto 0);
    signal conv10100_2583 : std_logic_vector(31 downto 0);
    signal conv13_2456 : std_logic_vector(31 downto 0);
    signal conv16_2461 : std_logic_vector(31 downto 0);
    signal conv23_2360 : std_logic_vector(31 downto 0);
    signal conv28_2379 : std_logic_vector(31 downto 0);
    signal conv34_2393 : std_logic_vector(31 downto 0);
    signal conv47_2527 : std_logic_vector(31 downto 0);
    signal conv50_2548 : std_logic_vector(31 downto 0);
    signal conv66_2660 : std_logic_vector(31 downto 0);
    signal conv76_2697 : std_logic_vector(31 downto 0);
    signal conv85_2723 : std_logic_vector(31 downto 0);
    signal conv_2322 : std_logic_vector(15 downto 0);
    signal div78_2435 : std_logic_vector(31 downto 0);
    signal div_2318 : std_logic_vector(31 downto 0);
    signal iNsTr_10_2425 : std_logic_vector(31 downto 0);
    signal iNsTr_2_2308 : std_logic_vector(31 downto 0);
    signal iNsTr_3_2330 : std_logic_vector(31 downto 0);
    signal iNsTr_4_2342 : std_logic_vector(31 downto 0);
    signal iNsTr_5_2352 : std_logic_vector(31 downto 0);
    signal iNsTr_6_2368 : std_logic_vector(31 downto 0);
    signal iNsTr_7_2385 : std_logic_vector(31 downto 0);
    signal iNsTr_8_2401 : std_logic_vector(31 downto 0);
    signal iNsTr_9_2413 : std_logic_vector(31 downto 0);
    signal idxprom62_2644 : std_logic_vector(63 downto 0);
    signal idxprom_2613 : std_logic_vector(63 downto 0);
    signal inc83_2706 : std_logic_vector(15 downto 0);
    signal inc83x_xinput_dim0x_x2_2711 : std_logic_vector(15 downto 0);
    signal inc_2692 : std_logic_vector(15 downto 0);
    signal indvar_2566 : std_logic_vector(15 downto 0);
    signal indvarx_xnext_2684 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2x_xph_2445 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1x_xph_2438 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_2718 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_2579 : std_logic_vector(15 downto 0);
    signal mul17_2476 : std_logic_vector(31 downto 0);
    signal mul24_2481 : std_logic_vector(31 downto 0);
    signal mul35_2496 : std_logic_vector(31 downto 0);
    signal mul51_2553 : std_logic_vector(31 downto 0);
    signal mul53_2563 : std_logic_vector(31 downto 0);
    signal mul_2466 : std_logic_vector(31 downto 0);
    signal ptr_deref_2311_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2311_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2311_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2311_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2311_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2333_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2333_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2333_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2333_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2333_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2345_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2345_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2345_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2345_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2345_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2355_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2355_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2355_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2355_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2355_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2371_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2371_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2371_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2371_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2371_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2388_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2388_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2388_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2388_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2388_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2404_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2404_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2404_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2404_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2404_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2416_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2416_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2416_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2416_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2416_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2428_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2428_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2428_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2428_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2428_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2623_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2623_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2623_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2623_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2623_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2653_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2653_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2653_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2653_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2653_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2653_word_offset_0 : std_logic_vector(13 downto 0);
    signal sext101_2539 : std_logic_vector(31 downto 0);
    signal sext103_2599 : std_logic_vector(31 downto 0);
    signal sext104_2630 : std_logic_vector(31 downto 0);
    signal sext_2518 : std_logic_vector(31 downto 0);
    signal shr61_2639 : std_logic_vector(31 downto 0);
    signal shr_2608 : std_logic_vector(31 downto 0);
    signal sub29_2533 : std_logic_vector(31 downto 0);
    signal sub40_2506 : std_logic_vector(31 downto 0);
    signal sub41_2512 : std_logic_vector(31 downto 0);
    signal sub_2491 : std_logic_vector(31 downto 0);
    signal tmp11_2334 : std_logic_vector(31 downto 0);
    signal tmp14_2346 : std_logic_vector(31 downto 0);
    signal tmp22_2356 : std_logic_vector(7 downto 0);
    signal tmp25_2372 : std_logic_vector(31 downto 0);
    signal tmp27_2375 : std_logic_vector(7 downto 0);
    signal tmp33_2389 : std_logic_vector(7 downto 0);
    signal tmp36_2405 : std_logic_vector(31 downto 0);
    signal tmp45_2417 : std_logic_vector(31 downto 0);
    signal tmp48_2429 : std_logic_vector(31 downto 0);
    signal tmp58_2624 : std_logic_vector(63 downto 0);
    signal tmp_2312 : std_logic_vector(31 downto 0);
    signal type_cast_2316_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2433_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2441_wire : std_logic_vector(15 downto 0);
    signal type_cast_2444_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2448_wire : std_logic_vector(15 downto 0);
    signal type_cast_2450_wire : std_logic_vector(15 downto 0);
    signal type_cast_2454_wire : std_logic_vector(31 downto 0);
    signal type_cast_2459_wire : std_logic_vector(31 downto 0);
    signal type_cast_2510_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2516_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2521_wire : std_logic_vector(31 downto 0);
    signal type_cast_2524_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2531_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2537_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2542_wire : std_logic_vector(31 downto 0);
    signal type_cast_2545_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2570_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2572_wire : std_logic_vector(15 downto 0);
    signal type_cast_2577_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2597_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2602_wire : std_logic_vector(31 downto 0);
    signal type_cast_2605_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2611_wire : std_logic_vector(63 downto 0);
    signal type_cast_2628_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2633_wire : std_logic_vector(31 downto 0);
    signal type_cast_2636_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2642_wire : std_logic_vector(63 downto 0);
    signal type_cast_2658_wire : std_logic_vector(31 downto 0);
    signal type_cast_2664_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2682_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2690_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2695_wire : std_logic_vector(31 downto 0);
    signal type_cast_2715_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2721_wire : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    LOAD_padding_2374_word_address_0 <= "0";
    array_obj_ref_2618_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2618_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2618_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2618_resized_base_address <= "00000000000000";
    array_obj_ref_2649_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2649_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2649_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2649_resized_base_address <= "00000000000000";
    iNsTr_10_2425 <= "00000000000000000000000000000100";
    iNsTr_2_2308 <= "00000000000000000000000000000011";
    iNsTr_3_2330 <= "00000000000000000000000000000101";
    iNsTr_4_2342 <= "00000000000000000000000000000100";
    iNsTr_5_2352 <= "00000000000000000000000000000000";
    iNsTr_6_2368 <= "00000000000000000000000000000100";
    iNsTr_7_2385 <= "00000000000000000000000000000001";
    iNsTr_8_2401 <= "00000000000000000000000000000101";
    iNsTr_9_2413 <= "00000000000000000000000000000101";
    ptr_deref_2311_word_offset_0 <= "0000000";
    ptr_deref_2333_word_offset_0 <= "0000000";
    ptr_deref_2345_word_offset_0 <= "0000000";
    ptr_deref_2355_word_offset_0 <= "0";
    ptr_deref_2371_word_offset_0 <= "0000000";
    ptr_deref_2388_word_offset_0 <= "0";
    ptr_deref_2404_word_offset_0 <= "0000000";
    ptr_deref_2416_word_offset_0 <= "0000000";
    ptr_deref_2428_word_offset_0 <= "0000000";
    ptr_deref_2623_word_offset_0 <= "00000000000000";
    ptr_deref_2653_word_offset_0 <= "00000000000000";
    type_cast_2316_wire_constant <= "00000000000000000000000000000001";
    type_cast_2433_wire_constant <= "00000000000000000000000000000001";
    type_cast_2444_wire_constant <= "0000000000000000";
    type_cast_2510_wire_constant <= "00000000000000000000000000010000";
    type_cast_2516_wire_constant <= "11111111111111110000000000000000";
    type_cast_2524_wire_constant <= "00000000000000000000000000010000";
    type_cast_2531_wire_constant <= "00000000000000000000000000010000";
    type_cast_2537_wire_constant <= "11111111111111110000000000000000";
    type_cast_2545_wire_constant <= "00000000000000000000000000010000";
    type_cast_2570_wire_constant <= "0000000000000000";
    type_cast_2577_wire_constant <= "0000000000000100";
    type_cast_2597_wire_constant <= "00000000000000000000000000010000";
    type_cast_2605_wire_constant <= "00000000000000000000000000010010";
    type_cast_2628_wire_constant <= "00000000000000000000000000010000";
    type_cast_2636_wire_constant <= "00000000000000000000000000010010";
    type_cast_2664_wire_constant <= "00000000000000000000000000000100";
    type_cast_2682_wire_constant <= "0000000000000001";
    type_cast_2690_wire_constant <= "0000000000000001";
    type_cast_2715_wire_constant <= "0000000000000000";
    phi_stmt_2438: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2441_wire & type_cast_2444_wire_constant;
      req <= phi_stmt_2438_req_0 & phi_stmt_2438_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2438",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2438_ack_0,
          idata => idata,
          odata => input_dim1x_x1x_xph_2438,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2438
    phi_stmt_2445: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2448_wire & type_cast_2450_wire;
      req <= phi_stmt_2445_req_0 & phi_stmt_2445_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2445",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2445_ack_0,
          idata => idata,
          odata => input_dim0x_x2x_xph_2445,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2445
    phi_stmt_2566: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2570_wire_constant & type_cast_2572_wire;
      req <= phi_stmt_2566_req_0 & phi_stmt_2566_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2566",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2566_ack_0,
          idata => idata,
          odata => indvar_2566,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2566
    -- flow-through select operator MUX_2717_inst
    input_dim1x_x2_2718 <= type_cast_2715_wire_constant when (cmp79_2702(0) /=  '0') else inc_2692;
    addr_of_2619_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2619_final_reg_req_0;
      addr_of_2619_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2619_final_reg_req_1;
      addr_of_2619_final_reg_ack_1<= rack(0);
      addr_of_2619_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2619_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2618_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_2620,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2650_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2650_final_reg_req_0;
      addr_of_2650_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2650_final_reg_req_1;
      addr_of_2650_final_reg_ack_1<= rack(0);
      addr_of_2650_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2650_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2649_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx63_2651,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2321_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2321_inst_req_0;
      type_cast_2321_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2321_inst_req_1;
      type_cast_2321_inst_ack_1<= rack(0);
      type_cast_2321_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2321_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div_2318,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_2322,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2359_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2359_inst_req_0;
      type_cast_2359_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2359_inst_req_1;
      type_cast_2359_inst_ack_1<= rack(0);
      type_cast_2359_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2359_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp22_2356,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv23_2360,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2378_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2378_inst_req_0;
      type_cast_2378_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2378_inst_req_1;
      type_cast_2378_inst_ack_1<= rack(0);
      type_cast_2378_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2378_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp27_2375,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv28_2379,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2392_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2392_inst_req_0;
      type_cast_2392_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2392_inst_req_1;
      type_cast_2392_inst_ack_1<= rack(0);
      type_cast_2392_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2392_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp33_2389,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv34_2393,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2441_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2441_inst_req_0;
      type_cast_2441_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2441_inst_req_1;
      type_cast_2441_inst_ack_1<= rack(0);
      type_cast_2441_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2441_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_2718,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2441_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2448_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2448_inst_req_0;
      type_cast_2448_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2448_inst_req_1;
      type_cast_2448_inst_ack_1<= rack(0);
      type_cast_2448_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2448_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc83x_xinput_dim0x_x2_2711,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2448_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2450_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2450_inst_req_0;
      type_cast_2450_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2450_inst_req_1;
      type_cast_2450_inst_ack_1<= rack(0);
      type_cast_2450_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2450_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv_2322,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2450_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2455_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2455_inst_req_0;
      type_cast_2455_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2455_inst_req_1;
      type_cast_2455_inst_ack_1<= rack(0);
      type_cast_2455_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2455_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2454_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv13_2456,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2460_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2460_inst_req_0;
      type_cast_2460_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2460_inst_req_1;
      type_cast_2460_inst_ack_1<= rack(0);
      type_cast_2460_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2460_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2459_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv16_2461,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2521_inst
    process(sext_2518) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext_2518(31 downto 0);
      type_cast_2521_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2526_inst
    process(ASHR_i32_i32_2525_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2525_wire(31 downto 0);
      conv47_2527 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2542_inst
    process(sext101_2539) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext101_2539(31 downto 0);
      type_cast_2542_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2547_inst
    process(ASHR_i32_i32_2546_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2546_wire(31 downto 0);
      conv50_2548 <= tmp_var; -- 
    end process;
    type_cast_2572_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2572_inst_req_0;
      type_cast_2572_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2572_inst_req_1;
      type_cast_2572_inst_ack_1<= rack(0);
      type_cast_2572_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2572_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_2684,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2572_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2582_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2582_inst_req_0;
      type_cast_2582_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2582_inst_req_1;
      type_cast_2582_inst_ack_1<= rack(0);
      type_cast_2582_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2582_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_2579,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv10100_2583,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2602_inst
    process(sext103_2599) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext103_2599(31 downto 0);
      type_cast_2602_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2607_inst
    process(ASHR_i32_i32_2606_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2606_wire(31 downto 0);
      shr_2608 <= tmp_var; -- 
    end process;
    type_cast_2612_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2612_inst_req_0;
      type_cast_2612_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2612_inst_req_1;
      type_cast_2612_inst_ack_1<= rack(0);
      type_cast_2612_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2612_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2611_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_2613,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2633_inst
    process(sext104_2630) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext104_2630(31 downto 0);
      type_cast_2633_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2638_inst
    process(ASHR_i32_i32_2637_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2637_wire(31 downto 0);
      shr61_2639 <= tmp_var; -- 
    end process;
    type_cast_2643_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2643_inst_req_0;
      type_cast_2643_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2643_inst_req_1;
      type_cast_2643_inst_ack_1<= rack(0);
      type_cast_2643_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2643_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2642_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom62_2644,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2659_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2659_inst_req_0;
      type_cast_2659_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2659_inst_req_1;
      type_cast_2659_inst_ack_1<= rack(0);
      type_cast_2659_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2659_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2658_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv66_2660,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2696_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2696_inst_req_0;
      type_cast_2696_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2696_inst_req_1;
      type_cast_2696_inst_ack_1<= rack(0);
      type_cast_2696_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2696_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2695_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv76_2697,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2705_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2705_inst_req_0;
      type_cast_2705_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2705_inst_req_1;
      type_cast_2705_inst_ack_1<= rack(0);
      type_cast_2705_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2705_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp79_2702,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc83_2706,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2722_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2722_inst_req_0;
      type_cast_2722_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2722_inst_req_1;
      type_cast_2722_inst_ack_1<= rack(0);
      type_cast_2722_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2722_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2721_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv85_2723,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence LOAD_padding_2374_gather_scatter
    process(LOAD_padding_2374_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_padding_2374_data_0;
      ov(7 downto 0) := iv;
      tmp27_2375 <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2618_index_1_rename
    process(R_idxprom_2617_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_2617_resized;
      ov(13 downto 0) := iv;
      R_idxprom_2617_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2618_index_1_resize
    process(idxprom_2613) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_2613;
      ov := iv(13 downto 0);
      R_idxprom_2617_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2618_root_address_inst
    process(array_obj_ref_2618_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2618_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2618_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2649_index_1_rename
    process(R_idxprom62_2648_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom62_2648_resized;
      ov(13 downto 0) := iv;
      R_idxprom62_2648_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2649_index_1_resize
    process(idxprom62_2644) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom62_2644;
      ov := iv(13 downto 0);
      R_idxprom62_2648_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2649_root_address_inst
    process(array_obj_ref_2649_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2649_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2649_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2311_addr_0
    process(ptr_deref_2311_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2311_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2311_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2311_base_resize
    process(iNsTr_2_2308) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_2_2308;
      ov := iv(6 downto 0);
      ptr_deref_2311_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2311_gather_scatter
    process(ptr_deref_2311_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2311_data_0;
      ov(31 downto 0) := iv;
      tmp_2312 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2311_root_address_inst
    process(ptr_deref_2311_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2311_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2311_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2333_addr_0
    process(ptr_deref_2333_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2333_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2333_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2333_base_resize
    process(iNsTr_3_2330) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_3_2330;
      ov := iv(6 downto 0);
      ptr_deref_2333_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2333_gather_scatter
    process(ptr_deref_2333_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2333_data_0;
      ov(31 downto 0) := iv;
      tmp11_2334 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2333_root_address_inst
    process(ptr_deref_2333_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2333_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2333_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2345_addr_0
    process(ptr_deref_2345_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2345_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2345_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2345_base_resize
    process(iNsTr_4_2342) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_4_2342;
      ov := iv(6 downto 0);
      ptr_deref_2345_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2345_gather_scatter
    process(ptr_deref_2345_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2345_data_0;
      ov(31 downto 0) := iv;
      tmp14_2346 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2345_root_address_inst
    process(ptr_deref_2345_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2345_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2345_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2355_addr_0
    process(ptr_deref_2355_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2355_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_2355_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2355_base_resize
    process(iNsTr_5_2352) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_5_2352;
      ov := iv(0 downto 0);
      ptr_deref_2355_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2355_gather_scatter
    process(ptr_deref_2355_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2355_data_0;
      ov(7 downto 0) := iv;
      tmp22_2356 <= ov(7 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2355_root_address_inst
    process(ptr_deref_2355_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2355_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_2355_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2371_addr_0
    process(ptr_deref_2371_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2371_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2371_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2371_base_resize
    process(iNsTr_6_2368) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_6_2368;
      ov := iv(6 downto 0);
      ptr_deref_2371_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2371_gather_scatter
    process(ptr_deref_2371_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2371_data_0;
      ov(31 downto 0) := iv;
      tmp25_2372 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2371_root_address_inst
    process(ptr_deref_2371_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2371_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2371_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2388_addr_0
    process(ptr_deref_2388_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2388_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_2388_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2388_base_resize
    process(iNsTr_7_2385) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_7_2385;
      ov := iv(0 downto 0);
      ptr_deref_2388_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2388_gather_scatter
    process(ptr_deref_2388_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2388_data_0;
      ov(7 downto 0) := iv;
      tmp33_2389 <= ov(7 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2388_root_address_inst
    process(ptr_deref_2388_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2388_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_2388_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2404_addr_0
    process(ptr_deref_2404_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2404_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2404_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2404_base_resize
    process(iNsTr_8_2401) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_8_2401;
      ov := iv(6 downto 0);
      ptr_deref_2404_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2404_gather_scatter
    process(ptr_deref_2404_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2404_data_0;
      ov(31 downto 0) := iv;
      tmp36_2405 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2404_root_address_inst
    process(ptr_deref_2404_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2404_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2404_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2416_addr_0
    process(ptr_deref_2416_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2416_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2416_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2416_base_resize
    process(iNsTr_9_2413) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_9_2413;
      ov := iv(6 downto 0);
      ptr_deref_2416_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2416_gather_scatter
    process(ptr_deref_2416_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2416_data_0;
      ov(31 downto 0) := iv;
      tmp45_2417 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2416_root_address_inst
    process(ptr_deref_2416_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2416_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2416_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2428_addr_0
    process(ptr_deref_2428_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2428_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2428_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2428_base_resize
    process(iNsTr_10_2425) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_10_2425;
      ov := iv(6 downto 0);
      ptr_deref_2428_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2428_gather_scatter
    process(ptr_deref_2428_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2428_data_0;
      ov(31 downto 0) := iv;
      tmp48_2429 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2428_root_address_inst
    process(ptr_deref_2428_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2428_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2428_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2623_addr_0
    process(ptr_deref_2623_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2623_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2623_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2623_base_resize
    process(arrayidx_2620) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_2620;
      ov := iv(13 downto 0);
      ptr_deref_2623_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2623_gather_scatter
    process(ptr_deref_2623_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2623_data_0;
      ov(63 downto 0) := iv;
      tmp58_2624 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2623_root_address_inst
    process(ptr_deref_2623_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2623_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2623_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2653_addr_0
    process(ptr_deref_2653_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2653_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2653_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2653_base_resize
    process(arrayidx63_2651) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx63_2651;
      ov := iv(13 downto 0);
      ptr_deref_2653_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2653_gather_scatter
    process(tmp58_2624) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp58_2624;
      ov(63 downto 0) := iv;
      ptr_deref_2653_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2653_root_address_inst
    process(ptr_deref_2653_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2653_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2653_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_2672_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_2671;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2672_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2672_branch_req_0,
          ack0 => if_stmt_2672_branch_ack_0,
          ack1 => if_stmt_2672_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2729_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp87_2728;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2729_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2729_branch_req_0,
          ack0 => if_stmt_2729_branch_ack_0,
          ack1 => if_stmt_2729_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_2683_inst
    process(indvar_2566) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_2566, type_cast_2682_wire_constant, tmp_var);
      indvarx_xnext_2684 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2691_inst
    process(input_dim1x_x1x_xph_2438) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_2438, type_cast_2690_wire_constant, tmp_var);
      inc_2692 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2710_inst
    process(inc83_2706, input_dim0x_x2x_xph_2445) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc83_2706, input_dim0x_x2x_xph_2445, tmp_var);
      inc83x_xinput_dim0x_x2_2711 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2470_inst
    process(mul_2466, conv13_2456) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul_2466, conv13_2456, tmp_var);
      add_2471 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2485_inst
    process(mul24_2481, tmp25_2372) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul24_2481, tmp25_2372, tmp_var);
      add26_2486 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2500_inst
    process(mul35_2496, tmp36_2405) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul35_2496, tmp36_2405, tmp_var);
      add37_2501 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2517_inst
    process(sub41_2512) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub41_2512, type_cast_2516_wire_constant, tmp_var);
      sext_2518 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2538_inst
    process(sub29_2533) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub29_2533, type_cast_2537_wire_constant, tmp_var);
      sext101_2539 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2557_inst
    process(conv47_2527, mul51_2553) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv47_2527, mul51_2553, tmp_var);
      add52_2558 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2587_inst
    process(mul17_2476, conv10100_2583) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul17_2476, conv10100_2583, tmp_var);
      add18_2588 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2592_inst
    process(mul53_2563, conv10100_2583) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul53_2563, conv10100_2583, tmp_var);
      add54_2593 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2665_inst
    process(conv66_2660) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv66_2660, type_cast_2664_wire_constant, tmp_var);
      add67_2666 <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2525_inst
    process(type_cast_2521_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2521_wire, type_cast_2524_wire_constant, tmp_var);
      ASHR_i32_i32_2525_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2546_inst
    process(type_cast_2542_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2542_wire, type_cast_2545_wire_constant, tmp_var);
      ASHR_i32_i32_2546_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2606_inst
    process(type_cast_2602_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2602_wire, type_cast_2605_wire_constant, tmp_var);
      ASHR_i32_i32_2606_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2637_inst
    process(type_cast_2633_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2633_wire, type_cast_2636_wire_constant, tmp_var);
      ASHR_i32_i32_2637_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2701_inst
    process(conv76_2697, div78_2435) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv76_2697, div78_2435, tmp_var);
      cmp79_2702 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2727_inst
    process(conv85_2723, tmp_2312) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv85_2723, tmp_2312, tmp_var);
      cmp87_2728 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2317_inst
    process(tmp_2312) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp_2312, type_cast_2316_wire_constant, tmp_var);
      div_2318 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2434_inst
    process(tmp14_2346) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp14_2346, type_cast_2433_wire_constant, tmp_var);
      div78_2435 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2578_inst
    process(indvar_2566) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_2566, type_cast_2577_wire_constant, tmp_var);
      input_dim2x_x1_2579 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2465_inst
    process(tmp14_2346, conv16_2461) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp14_2346, conv16_2461, tmp_var);
      mul_2466 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2475_inst
    process(add_2471, tmp11_2334) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add_2471, tmp11_2334, tmp_var);
      mul17_2476 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2480_inst
    process(conv23_2360, conv16_2461) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv23_2360, conv16_2461, tmp_var);
      mul24_2481 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2495_inst
    process(conv34_2393, conv13_2456) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv34_2393, conv13_2456, tmp_var);
      mul35_2496 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2552_inst
    process(tmp48_2429, conv50_2548) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp48_2429, conv50_2548, tmp_var);
      mul51_2553 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2562_inst
    process(add52_2558, tmp45_2417) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add52_2558, tmp45_2417, tmp_var);
      mul53_2563 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2511_inst
    process(sub40_2506) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(sub40_2506, type_cast_2510_wire_constant, tmp_var);
      sub41_2512 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2532_inst
    process(sub_2491) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(sub_2491, type_cast_2531_wire_constant, tmp_var);
      sub29_2533 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2598_inst
    process(add18_2588) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add18_2588, type_cast_2597_wire_constant, tmp_var);
      sext103_2599 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2629_inst
    process(add54_2593) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add54_2593, type_cast_2628_wire_constant, tmp_var);
      sext104_2630 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_2490_inst
    process(add26_2486, conv28_2379) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(add26_2486, conv28_2379, tmp_var);
      sub_2491 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_2505_inst
    process(add37_2501, conv28_2379) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(add37_2501, conv28_2379, tmp_var);
      sub40_2506 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_2670_inst
    process(add67_2666, tmp11_2334) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add67_2666, tmp11_2334, tmp_var);
      cmp_2671 <= tmp_var; --
    end process;
    -- shared split operator group (34) : array_obj_ref_2618_index_offset 
    ApIntAdd_group_34: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_2617_scaled;
      array_obj_ref_2618_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2618_index_offset_req_0;
      array_obj_ref_2618_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2618_index_offset_req_1;
      array_obj_ref_2618_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_34_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_34_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_34",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 34
    -- shared split operator group (35) : array_obj_ref_2649_index_offset 
    ApIntAdd_group_35: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom62_2648_scaled;
      array_obj_ref_2649_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2649_index_offset_req_0;
      array_obj_ref_2649_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2649_index_offset_req_1;
      array_obj_ref_2649_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_35_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_35_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_35",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 35
    -- unary operator type_cast_2454_inst
    process(input_dim1x_x1x_xph_2438) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim1x_x1x_xph_2438, tmp_var);
      type_cast_2454_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2459_inst
    process(input_dim0x_x2x_xph_2445) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim0x_x2x_xph_2445, tmp_var);
      type_cast_2459_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2611_inst
    process(shr_2608) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr_2608, tmp_var);
      type_cast_2611_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2642_inst
    process(shr61_2639) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr61_2639, tmp_var);
      type_cast_2642_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2658_inst
    process(input_dim2x_x1_2579) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim2x_x1_2579, tmp_var);
      type_cast_2658_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2695_inst
    process(inc_2692) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc_2692, tmp_var);
      type_cast_2695_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2721_inst
    process(inc83x_xinput_dim0x_x2_2711) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc83x_xinput_dim0x_x2_2711, tmp_var);
      type_cast_2721_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : LOAD_padding_2374_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_padding_2374_load_0_req_0;
      LOAD_padding_2374_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_padding_2374_load_0_req_1;
      LOAD_padding_2374_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_padding_2374_word_address_0;
      LOAD_padding_2374_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_7_lr_req(0),
          mack => memory_space_7_lr_ack(0),
          maddr => memory_space_7_lr_addr(0 downto 0),
          mtag => memory_space_7_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 8,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_7_lc_req(0),
          mack => memory_space_7_lc_ack(0),
          mdata => memory_space_7_lc_data(7 downto 0),
          mtag => memory_space_7_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_2311_load_0 ptr_deref_2333_load_0 ptr_deref_2345_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(20 downto 0);
      signal data_out: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_2311_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_2333_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2345_load_0_req_0;
      ptr_deref_2311_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_2333_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2345_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_2311_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_2333_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2345_load_0_req_1;
      ptr_deref_2311_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_2333_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2345_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      LoadGroup1_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2311_word_address_0 & ptr_deref_2333_word_address_0 & ptr_deref_2345_word_address_0;
      ptr_deref_2311_data_0 <= data_out(95 downto 64);
      ptr_deref_2333_data_0 <= data_out(63 downto 32);
      ptr_deref_2345_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 7,
        num_reqs => 3,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(6 downto 0),
          mtag => memory_space_1_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 32,
        num_reqs => 3,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(31 downto 0),
          mtag => memory_space_1_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : ptr_deref_2355_load_0 ptr_deref_2388_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_2355_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2388_load_0_req_0;
      ptr_deref_2355_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2388_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_2355_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2388_load_0_req_1;
      ptr_deref_2355_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2388_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup2_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup2_gI: SplitGuardInterface generic map(name => "LoadGroup2_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2355_word_address_0 & ptr_deref_2388_word_address_0;
      ptr_deref_2355_data_0 <= data_out(15 downto 8);
      ptr_deref_2388_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup2", addr_width => 1,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_8_lr_req(0),
          mack => memory_space_8_lr_ack(0),
          maddr => memory_space_8_lr_addr(0 downto 0),
          mtag => memory_space_8_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup2 load-complete ",
        data_width => 8,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_8_lc_req(0),
          mack => memory_space_8_lc_ack(0),
          mdata => memory_space_8_lc_data(7 downto 0),
          mtag => memory_space_8_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared load operator group (3) : ptr_deref_2371_load_0 ptr_deref_2404_load_0 
    LoadGroup3: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_2371_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2404_load_0_req_0;
      ptr_deref_2371_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2404_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_2371_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2404_load_0_req_1;
      ptr_deref_2371_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2404_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup3_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup3_gI: SplitGuardInterface generic map(name => "LoadGroup3_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2371_word_address_0 & ptr_deref_2404_word_address_0;
      ptr_deref_2371_data_0 <= data_out(63 downto 32);
      ptr_deref_2404_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup3", addr_width => 7,
        num_reqs => 2,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(6 downto 0),
          mtag => memory_space_2_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup3 load-complete ",
        data_width => 32,
        num_reqs => 2,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(31 downto 0),
          mtag => memory_space_2_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 3
    -- shared load operator group (4) : ptr_deref_2416_load_0 ptr_deref_2428_load_0 
    LoadGroup4: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_2416_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2428_load_0_req_0;
      ptr_deref_2416_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2428_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_2416_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2428_load_0_req_1;
      ptr_deref_2416_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2428_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup4_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup4_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup4_gI: SplitGuardInterface generic map(name => "LoadGroup4_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2416_word_address_0 & ptr_deref_2428_word_address_0;
      ptr_deref_2416_data_0 <= data_out(63 downto 32);
      ptr_deref_2428_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup4", addr_width => 7,
        num_reqs => 2,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(6 downto 0),
          mtag => memory_space_3_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup4 load-complete ",
        data_width => 32,
        num_reqs => 2,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(31 downto 0),
          mtag => memory_space_3_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 4
    -- shared load operator group (5) : ptr_deref_2623_load_0 
    LoadGroup5: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2623_load_0_req_0;
      ptr_deref_2623_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2623_load_0_req_1;
      ptr_deref_2623_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup5_gI: SplitGuardInterface generic map(name => "LoadGroup5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2623_word_address_0;
      ptr_deref_2623_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup5", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_4_lr_req(0),
          mack => memory_space_4_lr_ack(0),
          maddr => memory_space_4_lr_addr(13 downto 0),
          mtag => memory_space_4_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup5 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_4_lc_req(0),
          mack => memory_space_4_lc_ack(0),
          mdata => memory_space_4_lc_data(63 downto 0),
          mtag => memory_space_4_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 5
    -- shared store operator group (0) : ptr_deref_2653_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2653_store_0_req_0;
      ptr_deref_2653_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2653_store_0_req_1;
      ptr_deref_2653_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_2653_word_address_0;
      data_in <= ptr_deref_2653_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_6_sr_req(0),
          mack => memory_space_6_sr_ack(0),
          maddr => memory_space_6_sr_addr(13 downto 0),
          mdata => memory_space_6_sr_data(63 downto 0),
          mtag => memory_space_6_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_6_sc_req(0),
          mack => memory_space_6_sc_ack(0),
          mtag => memory_space_6_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block2_start_2298_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block2_start_2298_inst_req_0;
      RPIPE_Block2_start_2298_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block2_start_2298_inst_req_1;
      RPIPE_Block2_start_2298_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call_2299 <= data_out(15 downto 0);
      Block2_start_read_0_gI: SplitGuardInterface generic map(name => "Block2_start_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block2_start_read_0: InputPortRevised -- 
        generic map ( name => "Block2_start_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block2_start_pipe_read_req(0),
          oack => Block2_start_pipe_read_ack(0),
          odata => Block2_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block2_done_2737_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block2_done_2737_inst_req_0;
      WPIPE_Block2_done_2737_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block2_done_2737_inst_req_1;
      WPIPE_Block2_done_2737_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= call_2299;
      Block2_done_write_0_gI: SplitGuardInterface generic map(name => "Block2_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block2_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block2_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block2_done_pipe_write_req(0),
          oack => Block2_done_pipe_write_ack(0),
          odata => Block2_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeC_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeD is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_7_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_8_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_8_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_8_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_8_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_8_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_8_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_4_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_4_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_6_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_6_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_sc_tag :  in  std_logic_vector(0 downto 0);
    Block3_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block3_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block3_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block3_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block3_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block3_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeD;
architecture convTransposeD_arch of convTransposeD is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeD_CP_7576_start: Boolean;
  signal convTransposeD_CP_7576_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal type_cast_2912_inst_req_0 : boolean;
  signal type_cast_2907_inst_req_1 : boolean;
  signal type_cast_3034_inst_ack_0 : boolean;
  signal type_cast_3034_inst_req_0 : boolean;
  signal ptr_deref_2875_load_0_ack_1 : boolean;
  signal ptr_deref_2875_load_0_req_1 : boolean;
  signal type_cast_3064_inst_ack_0 : boolean;
  signal type_cast_3064_inst_req_0 : boolean;
  signal array_obj_ref_3070_index_offset_ack_0 : boolean;
  signal array_obj_ref_3070_index_offset_req_1 : boolean;
  signal ptr_deref_2887_load_0_req_0 : boolean;
  signal type_cast_2907_inst_req_0 : boolean;
  signal addr_of_3071_final_reg_ack_1 : boolean;
  signal addr_of_3071_final_reg_req_0 : boolean;
  signal addr_of_3071_final_reg_req_1 : boolean;
  signal array_obj_ref_3070_index_offset_ack_1 : boolean;
  signal addr_of_3071_final_reg_ack_0 : boolean;
  signal ptr_deref_2887_load_0_req_1 : boolean;
  signal array_obj_ref_3070_index_offset_req_0 : boolean;
  signal ptr_deref_2887_load_0_ack_0 : boolean;
  signal ptr_deref_2887_load_0_ack_1 : boolean;
  signal type_cast_2912_inst_req_1 : boolean;
  signal type_cast_3034_inst_req_1 : boolean;
  signal type_cast_2912_inst_ack_1 : boolean;
  signal ptr_deref_2875_load_0_req_0 : boolean;
  signal type_cast_3034_inst_ack_1 : boolean;
  signal ptr_deref_2875_load_0_ack_0 : boolean;
  signal type_cast_2912_inst_ack_0 : boolean;
  signal type_cast_2907_inst_ack_1 : boolean;
  signal type_cast_2907_inst_ack_0 : boolean;
  signal type_cast_3064_inst_ack_1 : boolean;
  signal type_cast_3064_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2747_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2747_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2747_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2747_inst_ack_1 : boolean;
  signal ptr_deref_2760_load_0_req_0 : boolean;
  signal ptr_deref_2760_load_0_ack_0 : boolean;
  signal ptr_deref_2760_load_0_req_1 : boolean;
  signal ptr_deref_2760_load_0_ack_1 : boolean;
  signal type_cast_2770_inst_req_0 : boolean;
  signal type_cast_2770_inst_ack_0 : boolean;
  signal type_cast_2770_inst_req_1 : boolean;
  signal type_cast_2770_inst_ack_1 : boolean;
  signal ptr_deref_2782_load_0_req_0 : boolean;
  signal ptr_deref_2782_load_0_ack_0 : boolean;
  signal ptr_deref_2782_load_0_req_1 : boolean;
  signal ptr_deref_2782_load_0_ack_1 : boolean;
  signal type_cast_2792_inst_req_0 : boolean;
  signal type_cast_2792_inst_ack_0 : boolean;
  signal type_cast_2792_inst_req_1 : boolean;
  signal type_cast_2792_inst_ack_1 : boolean;
  signal ptr_deref_2804_load_0_req_0 : boolean;
  signal ptr_deref_2804_load_0_ack_0 : boolean;
  signal ptr_deref_2804_load_0_req_1 : boolean;
  signal ptr_deref_2804_load_0_ack_1 : boolean;
  signal ptr_deref_2814_load_0_req_0 : boolean;
  signal ptr_deref_2814_load_0_ack_0 : boolean;
  signal ptr_deref_2814_load_0_req_1 : boolean;
  signal ptr_deref_2814_load_0_ack_1 : boolean;
  signal type_cast_2818_inst_req_0 : boolean;
  signal type_cast_2818_inst_ack_0 : boolean;
  signal type_cast_2818_inst_req_1 : boolean;
  signal type_cast_2818_inst_ack_1 : boolean;
  signal ptr_deref_2830_load_0_req_0 : boolean;
  signal ptr_deref_2830_load_0_ack_0 : boolean;
  signal ptr_deref_2830_load_0_req_1 : boolean;
  signal ptr_deref_2830_load_0_ack_1 : boolean;
  signal LOAD_padding_2833_load_0_req_0 : boolean;
  signal LOAD_padding_2833_load_0_ack_0 : boolean;
  signal LOAD_padding_2833_load_0_req_1 : boolean;
  signal LOAD_padding_2833_load_0_ack_1 : boolean;
  signal type_cast_2837_inst_req_0 : boolean;
  signal type_cast_2837_inst_ack_0 : boolean;
  signal type_cast_2837_inst_req_1 : boolean;
  signal type_cast_2837_inst_ack_1 : boolean;
  signal ptr_deref_2847_load_0_req_0 : boolean;
  signal ptr_deref_2847_load_0_ack_0 : boolean;
  signal ptr_deref_2847_load_0_req_1 : boolean;
  signal ptr_deref_2847_load_0_ack_1 : boolean;
  signal type_cast_2851_inst_req_0 : boolean;
  signal type_cast_2851_inst_ack_0 : boolean;
  signal type_cast_2851_inst_req_1 : boolean;
  signal type_cast_2851_inst_ack_1 : boolean;
  signal ptr_deref_2863_load_0_req_0 : boolean;
  signal ptr_deref_2863_load_0_ack_0 : boolean;
  signal ptr_deref_2863_load_0_req_1 : boolean;
  signal ptr_deref_2863_load_0_ack_1 : boolean;
  signal ptr_deref_3075_load_0_req_0 : boolean;
  signal ptr_deref_3075_load_0_ack_0 : boolean;
  signal ptr_deref_3075_load_0_req_1 : boolean;
  signal ptr_deref_3075_load_0_ack_1 : boolean;
  signal type_cast_3095_inst_req_0 : boolean;
  signal type_cast_3095_inst_ack_0 : boolean;
  signal type_cast_3095_inst_req_1 : boolean;
  signal type_cast_3095_inst_ack_1 : boolean;
  signal array_obj_ref_3101_index_offset_req_0 : boolean;
  signal array_obj_ref_3101_index_offset_ack_0 : boolean;
  signal array_obj_ref_3101_index_offset_req_1 : boolean;
  signal array_obj_ref_3101_index_offset_ack_1 : boolean;
  signal addr_of_3102_final_reg_req_0 : boolean;
  signal addr_of_3102_final_reg_ack_0 : boolean;
  signal addr_of_3102_final_reg_req_1 : boolean;
  signal addr_of_3102_final_reg_ack_1 : boolean;
  signal ptr_deref_3105_store_0_req_0 : boolean;
  signal ptr_deref_3105_store_0_ack_0 : boolean;
  signal ptr_deref_3105_store_0_req_1 : boolean;
  signal ptr_deref_3105_store_0_ack_1 : boolean;
  signal type_cast_3111_inst_req_0 : boolean;
  signal type_cast_3111_inst_ack_0 : boolean;
  signal type_cast_3111_inst_req_1 : boolean;
  signal type_cast_3111_inst_ack_1 : boolean;
  signal if_stmt_3124_branch_req_0 : boolean;
  signal if_stmt_3124_branch_ack_1 : boolean;
  signal if_stmt_3124_branch_ack_0 : boolean;
  signal type_cast_3148_inst_req_0 : boolean;
  signal type_cast_3148_inst_ack_0 : boolean;
  signal type_cast_3148_inst_req_1 : boolean;
  signal type_cast_3148_inst_ack_1 : boolean;
  signal if_stmt_3155_branch_req_0 : boolean;
  signal if_stmt_3155_branch_ack_1 : boolean;
  signal if_stmt_3155_branch_ack_0 : boolean;
  signal type_cast_3176_inst_req_0 : boolean;
  signal type_cast_3176_inst_ack_0 : boolean;
  signal type_cast_3176_inst_req_1 : boolean;
  signal type_cast_3176_inst_ack_1 : boolean;
  signal type_cast_3196_inst_req_0 : boolean;
  signal type_cast_3196_inst_ack_0 : boolean;
  signal type_cast_3196_inst_req_1 : boolean;
  signal type_cast_3196_inst_ack_1 : boolean;
  signal if_stmt_3203_branch_req_0 : boolean;
  signal if_stmt_3203_branch_ack_1 : boolean;
  signal if_stmt_3203_branch_ack_0 : boolean;
  signal WPIPE_Block3_done_3211_inst_req_0 : boolean;
  signal WPIPE_Block3_done_3211_inst_ack_0 : boolean;
  signal WPIPE_Block3_done_3211_inst_req_1 : boolean;
  signal WPIPE_Block3_done_3211_inst_ack_1 : boolean;
  signal type_cast_2894_inst_req_0 : boolean;
  signal type_cast_2894_inst_ack_0 : boolean;
  signal type_cast_2894_inst_req_1 : boolean;
  signal type_cast_2894_inst_ack_1 : boolean;
  signal phi_stmt_2891_req_0 : boolean;
  signal type_cast_2900_inst_req_0 : boolean;
  signal type_cast_2900_inst_ack_0 : boolean;
  signal type_cast_2900_inst_req_1 : boolean;
  signal type_cast_2900_inst_ack_1 : boolean;
  signal phi_stmt_2897_req_0 : boolean;
  signal type_cast_2896_inst_req_0 : boolean;
  signal type_cast_2896_inst_ack_0 : boolean;
  signal type_cast_2896_inst_req_1 : boolean;
  signal type_cast_2896_inst_ack_1 : boolean;
  signal phi_stmt_2891_req_1 : boolean;
  signal type_cast_2902_inst_req_0 : boolean;
  signal type_cast_2902_inst_ack_0 : boolean;
  signal type_cast_2902_inst_req_1 : boolean;
  signal type_cast_2902_inst_ack_1 : boolean;
  signal phi_stmt_2897_req_1 : boolean;
  signal phi_stmt_2891_ack_0 : boolean;
  signal phi_stmt_2897_ack_0 : boolean;
  signal type_cast_3024_inst_req_0 : boolean;
  signal type_cast_3024_inst_ack_0 : boolean;
  signal type_cast_3024_inst_req_1 : boolean;
  signal type_cast_3024_inst_ack_1 : boolean;
  signal phi_stmt_3018_req_1 : boolean;
  signal phi_stmt_3018_req_0 : boolean;
  signal phi_stmt_3018_ack_0 : boolean;
  signal type_cast_3185_inst_req_0 : boolean;
  signal type_cast_3185_inst_ack_0 : boolean;
  signal type_cast_3185_inst_req_1 : boolean;
  signal type_cast_3185_inst_ack_1 : boolean;
  signal phi_stmt_3180_req_1 : boolean;
  signal type_cast_3191_inst_req_0 : boolean;
  signal type_cast_3191_inst_ack_0 : boolean;
  signal type_cast_3191_inst_req_1 : boolean;
  signal type_cast_3191_inst_ack_1 : boolean;
  signal phi_stmt_3186_req_1 : boolean;
  signal type_cast_3183_inst_req_0 : boolean;
  signal type_cast_3183_inst_ack_0 : boolean;
  signal type_cast_3183_inst_req_1 : boolean;
  signal type_cast_3183_inst_ack_1 : boolean;
  signal phi_stmt_3180_req_0 : boolean;
  signal type_cast_3189_inst_req_0 : boolean;
  signal type_cast_3189_inst_ack_0 : boolean;
  signal type_cast_3189_inst_req_1 : boolean;
  signal type_cast_3189_inst_ack_1 : boolean;
  signal phi_stmt_3186_req_0 : boolean;
  signal phi_stmt_3180_ack_0 : boolean;
  signal phi_stmt_3186_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeD_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeD_CP_7576_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeD_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeD_CP_7576_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeD_CP_7576_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeD_CP_7576_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeD_CP_7576: Block -- control-path 
    signal convTransposeD_CP_7576_elements: BooleanArray(116 downto 0);
    -- 
  begin -- 
    convTransposeD_CP_7576_elements(0) <= convTransposeD_CP_7576_start;
    convTransposeD_CP_7576_symbol <= convTransposeD_CP_7576_elements(74);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 branch_block_stmt_2745/assign_stmt_2748__entry__
      -- CP-element group 0: 	 branch_block_stmt_2745/branch_block_stmt_2745__entry__
      -- CP-element group 0: 	 branch_block_stmt_2745/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_2745/assign_stmt_2748/$entry
      -- CP-element group 0: 	 branch_block_stmt_2745/assign_stmt_2748/RPIPE_Block3_start_2747_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_2745/assign_stmt_2748/RPIPE_Block3_start_2747_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_2745/assign_stmt_2748/RPIPE_Block3_start_2747_Sample/rr
      -- 
    rr_7634_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7634_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(0), ack => RPIPE_Block3_start_2747_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_2745/assign_stmt_2748/RPIPE_Block3_start_2747_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_2745/assign_stmt_2748/RPIPE_Block3_start_2747_update_start_
      -- CP-element group 1: 	 branch_block_stmt_2745/assign_stmt_2748/RPIPE_Block3_start_2747_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_2745/assign_stmt_2748/RPIPE_Block3_start_2747_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_2745/assign_stmt_2748/RPIPE_Block3_start_2747_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2745/assign_stmt_2748/RPIPE_Block3_start_2747_Update/cr
      -- 
    ra_7635_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2747_inst_ack_0, ack => convTransposeD_CP_7576_elements(1)); -- 
    cr_7639_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7639_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(1), ack => RPIPE_Block3_start_2747_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  place  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	29 
    -- CP-element group 2: 	14 
    -- CP-element group 2: 	30 
    -- CP-element group 2: 	20 
    -- CP-element group 2: 	23 
    -- CP-element group 2: 	22 
    -- CP-element group 2: 	13 
    -- CP-element group 2: 	28 
    -- CP-element group 2: 	16 
    -- CP-element group 2: 	27 
    -- CP-element group 2: 	31 
    -- CP-element group 2: 	17 
    -- CP-element group 2: 	24 
    -- CP-element group 2: 	26 
    -- CP-element group 2: 	19 
    -- CP-element group 2: 	32 
    -- CP-element group 2: 	18 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	4 
    -- CP-element group 2: 	6 
    -- CP-element group 2: 	7 
    -- CP-element group 2: 	8 
    -- CP-element group 2: 	10 
    -- CP-element group 2: 	11 
    -- CP-element group 2: 	12 
    -- CP-element group 2:  members (268) 
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2887_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2887_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2875_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2875_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2875_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2887_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2875_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2887_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2875_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2875_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2875_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2875_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2887_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2875_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2875_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2875_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2887_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2875_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2887_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2887_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2875_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2887_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2887_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2875_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2887_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2875_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2887_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2875_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2875_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2875_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2875_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2887_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888__entry__
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2887_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2887_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2748__exit__
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2887_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2887_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2887_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2887_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2887_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2887_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2875_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2875_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2875_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2875_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2887_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2875_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2875_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2887_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2887_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2875_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2887_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2748/$exit
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2887_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2748/RPIPE_Block3_start_2747_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2748/RPIPE_Block3_start_2747_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2748/RPIPE_Block3_start_2747_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2760_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2760_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2760_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2760_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2760_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2760_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2760_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2760_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2760_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2760_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2760_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2760_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2760_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2760_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2760_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2760_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2760_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2760_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2760_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2760_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2760_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2760_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2760_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2760_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2760_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2760_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/type_cast_2770_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/type_cast_2770_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/type_cast_2770_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2782_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2782_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2782_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2782_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2782_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2782_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2782_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2782_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2782_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2782_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2782_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2782_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2782_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2782_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2782_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2782_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2782_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2782_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2782_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2782_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2782_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2782_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2782_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2782_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2782_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2782_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/type_cast_2792_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/type_cast_2792_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/type_cast_2792_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2804_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2804_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2804_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2804_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2804_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2804_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2804_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2804_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2804_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2804_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2804_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2804_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2804_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2804_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2804_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2804_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2804_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2804_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2804_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2804_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2804_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2804_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2804_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2804_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2804_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2804_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2814_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2814_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2814_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2814_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2814_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2814_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2814_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2814_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2814_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2814_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2814_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2814_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2814_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2814_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2814_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2814_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2814_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2814_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2814_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2814_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2814_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2814_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2814_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2814_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2814_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2814_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/type_cast_2818_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/type_cast_2818_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/type_cast_2818_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2830_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2830_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2830_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2830_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2830_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2830_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2830_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2830_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2830_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2830_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2830_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2830_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2830_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2830_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2830_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2830_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2830_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2830_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2830_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2830_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2830_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2830_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2830_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2830_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2830_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2830_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/LOAD_padding_2833_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/LOAD_padding_2833_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/LOAD_padding_2833_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/LOAD_padding_2833_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/LOAD_padding_2833_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/LOAD_padding_2833_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/LOAD_padding_2833_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/LOAD_padding_2833_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/LOAD_padding_2833_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/LOAD_padding_2833_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/LOAD_padding_2833_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/LOAD_padding_2833_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/type_cast_2837_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/type_cast_2837_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/type_cast_2837_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2847_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2847_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2847_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2847_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2847_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2847_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2847_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2847_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2847_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2847_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2847_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2847_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2847_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2847_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2847_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2847_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2847_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2847_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2847_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2847_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2847_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2847_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2847_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2847_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2847_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2847_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/type_cast_2851_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/type_cast_2851_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/type_cast_2851_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2863_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2863_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2863_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2863_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2863_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2863_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2863_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2863_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2863_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2863_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2863_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2863_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2863_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2863_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2863_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2863_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2863_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2863_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2863_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2863_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2863_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2863_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2863_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2863_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2863_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2863_Update/word_access_complete/word_0/cr
      -- 
    ca_7640_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2747_inst_ack_1, ack => convTransposeD_CP_7576_elements(2)); -- 
    cr_8140_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8140_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(2), ack => ptr_deref_2875_load_0_req_1); -- 
    rr_8179_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8179_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(2), ack => ptr_deref_2887_load_0_req_0); -- 
    cr_8190_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8190_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(2), ack => ptr_deref_2887_load_0_req_1); -- 
    rr_8129_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8129_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(2), ack => ptr_deref_2875_load_0_req_0); -- 
    rr_7676_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7676_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(2), ack => ptr_deref_2760_load_0_req_0); -- 
    cr_7687_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7687_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(2), ack => ptr_deref_2760_load_0_req_1); -- 
    cr_7706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(2), ack => type_cast_2770_inst_req_1); -- 
    rr_7740_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7740_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(2), ack => ptr_deref_2782_load_0_req_0); -- 
    cr_7751_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7751_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(2), ack => ptr_deref_2782_load_0_req_1); -- 
    cr_7770_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7770_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(2), ack => type_cast_2792_inst_req_1); -- 
    rr_7804_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7804_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(2), ack => ptr_deref_2804_load_0_req_0); -- 
    cr_7815_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7815_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(2), ack => ptr_deref_2804_load_0_req_1); -- 
    rr_7854_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7854_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(2), ack => ptr_deref_2814_load_0_req_0); -- 
    cr_7865_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7865_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(2), ack => ptr_deref_2814_load_0_req_1); -- 
    cr_7884_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7884_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(2), ack => type_cast_2818_inst_req_1); -- 
    rr_7918_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7918_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(2), ack => ptr_deref_2830_load_0_req_0); -- 
    cr_7929_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7929_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(2), ack => ptr_deref_2830_load_0_req_1); -- 
    rr_7951_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7951_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(2), ack => LOAD_padding_2833_load_0_req_0); -- 
    cr_7962_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7962_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(2), ack => LOAD_padding_2833_load_0_req_1); -- 
    cr_7981_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7981_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(2), ack => type_cast_2837_inst_req_1); -- 
    rr_8015_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8015_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(2), ack => ptr_deref_2847_load_0_req_0); -- 
    cr_8026_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8026_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(2), ack => ptr_deref_2847_load_0_req_1); -- 
    cr_8045_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8045_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(2), ack => type_cast_2851_inst_req_1); -- 
    rr_8079_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8079_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(2), ack => ptr_deref_2863_load_0_req_0); -- 
    cr_8090_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8090_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(2), ack => ptr_deref_2863_load_0_req_1); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (5) 
      -- CP-element group 3: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2760_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2760_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2760_Sample/word_access_start/$exit
      -- CP-element group 3: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2760_Sample/word_access_start/word_0/$exit
      -- CP-element group 3: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2760_Sample/word_access_start/word_0/ra
      -- 
    ra_7677_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2760_load_0_ack_0, ack => convTransposeD_CP_7576_elements(3)); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	2 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (12) 
      -- CP-element group 4: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2760_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2760_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2760_Update/word_access_complete/$exit
      -- CP-element group 4: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2760_Update/word_access_complete/word_0/$exit
      -- CP-element group 4: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2760_Update/word_access_complete/word_0/ca
      -- CP-element group 4: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2760_Update/ptr_deref_2760_Merge/$entry
      -- CP-element group 4: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2760_Update/ptr_deref_2760_Merge/$exit
      -- CP-element group 4: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2760_Update/ptr_deref_2760_Merge/merge_req
      -- CP-element group 4: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2760_Update/ptr_deref_2760_Merge/merge_ack
      -- CP-element group 4: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/type_cast_2770_sample_start_
      -- CP-element group 4: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/type_cast_2770_Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/type_cast_2770_Sample/rr
      -- 
    ca_7688_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2760_load_0_ack_1, ack => convTransposeD_CP_7576_elements(4)); -- 
    rr_7701_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7701_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(4), ack => type_cast_2770_inst_req_0); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/type_cast_2770_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/type_cast_2770_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/type_cast_2770_Sample/ra
      -- 
    ra_7702_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2770_inst_ack_0, ack => convTransposeD_CP_7576_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	2 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	33 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/type_cast_2770_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/type_cast_2770_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/type_cast_2770_Update/ca
      -- 
    ca_7707_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2770_inst_ack_1, ack => convTransposeD_CP_7576_elements(6)); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	2 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (5) 
      -- CP-element group 7: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2782_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2782_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2782_Sample/word_access_start/$exit
      -- CP-element group 7: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2782_Sample/word_access_start/word_0/$exit
      -- CP-element group 7: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2782_Sample/word_access_start/word_0/ra
      -- 
    ra_7741_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2782_load_0_ack_0, ack => convTransposeD_CP_7576_elements(7)); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (12) 
      -- CP-element group 8: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2782_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2782_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2782_Update/word_access_complete/$exit
      -- CP-element group 8: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2782_Update/word_access_complete/word_0/$exit
      -- CP-element group 8: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2782_Update/word_access_complete/word_0/ca
      -- CP-element group 8: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2782_Update/ptr_deref_2782_Merge/$entry
      -- CP-element group 8: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2782_Update/ptr_deref_2782_Merge/$exit
      -- CP-element group 8: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2782_Update/ptr_deref_2782_Merge/merge_req
      -- CP-element group 8: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2782_Update/ptr_deref_2782_Merge/merge_ack
      -- CP-element group 8: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/type_cast_2792_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/type_cast_2792_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/type_cast_2792_Sample/rr
      -- 
    ca_7752_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2782_load_0_ack_1, ack => convTransposeD_CP_7576_elements(8)); -- 
    rr_7765_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7765_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(8), ack => type_cast_2792_inst_req_0); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/type_cast_2792_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/type_cast_2792_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/type_cast_2792_Sample/ra
      -- 
    ra_7766_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2792_inst_ack_0, ack => convTransposeD_CP_7576_elements(9)); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	2 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	33 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/type_cast_2792_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/type_cast_2792_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/type_cast_2792_Update/ca
      -- 
    ca_7771_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2792_inst_ack_1, ack => convTransposeD_CP_7576_elements(10)); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	2 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (5) 
      -- CP-element group 11: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2804_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2804_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2804_Sample/word_access_start/$exit
      -- CP-element group 11: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2804_Sample/word_access_start/word_0/$exit
      -- CP-element group 11: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2804_Sample/word_access_start/word_0/ra
      -- 
    ra_7805_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2804_load_0_ack_0, ack => convTransposeD_CP_7576_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	2 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	33 
    -- CP-element group 12:  members (9) 
      -- CP-element group 12: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2804_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2804_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2804_Update/word_access_complete/$exit
      -- CP-element group 12: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2804_Update/word_access_complete/word_0/$exit
      -- CP-element group 12: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2804_Update/word_access_complete/word_0/ca
      -- CP-element group 12: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2804_Update/ptr_deref_2804_Merge/$entry
      -- CP-element group 12: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2804_Update/ptr_deref_2804_Merge/$exit
      -- CP-element group 12: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2804_Update/ptr_deref_2804_Merge/merge_req
      -- CP-element group 12: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2804_Update/ptr_deref_2804_Merge/merge_ack
      -- 
    ca_7816_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2804_load_0_ack_1, ack => convTransposeD_CP_7576_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	2 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (5) 
      -- CP-element group 13: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2814_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2814_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2814_Sample/word_access_start/$exit
      -- CP-element group 13: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2814_Sample/word_access_start/word_0/$exit
      -- CP-element group 13: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2814_Sample/word_access_start/word_0/ra
      -- 
    ra_7855_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2814_load_0_ack_0, ack => convTransposeD_CP_7576_elements(13)); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	2 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (12) 
      -- CP-element group 14: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2814_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2814_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2814_Update/word_access_complete/$exit
      -- CP-element group 14: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2814_Update/word_access_complete/word_0/$exit
      -- CP-element group 14: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2814_Update/word_access_complete/word_0/ca
      -- CP-element group 14: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2814_Update/ptr_deref_2814_Merge/$entry
      -- CP-element group 14: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2814_Update/ptr_deref_2814_Merge/$exit
      -- CP-element group 14: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2814_Update/ptr_deref_2814_Merge/merge_req
      -- CP-element group 14: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2814_Update/ptr_deref_2814_Merge/merge_ack
      -- CP-element group 14: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/type_cast_2818_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/type_cast_2818_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/type_cast_2818_Sample/rr
      -- 
    ca_7866_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2814_load_0_ack_1, ack => convTransposeD_CP_7576_elements(14)); -- 
    rr_7879_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7879_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(14), ack => type_cast_2818_inst_req_0); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/type_cast_2818_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/type_cast_2818_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/type_cast_2818_Sample/ra
      -- 
    ra_7880_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2818_inst_ack_0, ack => convTransposeD_CP_7576_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	2 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	33 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/type_cast_2818_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/type_cast_2818_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/type_cast_2818_Update/ca
      -- 
    ca_7885_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2818_inst_ack_1, ack => convTransposeD_CP_7576_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	2 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (5) 
      -- CP-element group 17: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2830_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2830_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2830_Sample/word_access_start/$exit
      -- CP-element group 17: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2830_Sample/word_access_start/word_0/$exit
      -- CP-element group 17: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2830_Sample/word_access_start/word_0/ra
      -- 
    ra_7919_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2830_load_0_ack_0, ack => convTransposeD_CP_7576_elements(17)); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	2 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	33 
    -- CP-element group 18:  members (9) 
      -- CP-element group 18: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2830_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2830_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2830_Update/word_access_complete/$exit
      -- CP-element group 18: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2830_Update/word_access_complete/word_0/$exit
      -- CP-element group 18: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2830_Update/word_access_complete/word_0/ca
      -- CP-element group 18: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2830_Update/ptr_deref_2830_Merge/$entry
      -- CP-element group 18: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2830_Update/ptr_deref_2830_Merge/$exit
      -- CP-element group 18: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2830_Update/ptr_deref_2830_Merge/merge_req
      -- CP-element group 18: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2830_Update/ptr_deref_2830_Merge/merge_ack
      -- 
    ca_7930_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2830_load_0_ack_1, ack => convTransposeD_CP_7576_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	2 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (5) 
      -- CP-element group 19: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/LOAD_padding_2833_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/LOAD_padding_2833_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/LOAD_padding_2833_Sample/word_access_start/$exit
      -- CP-element group 19: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/LOAD_padding_2833_Sample/word_access_start/word_0/$exit
      -- CP-element group 19: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/LOAD_padding_2833_Sample/word_access_start/word_0/ra
      -- 
    ra_7952_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_padding_2833_load_0_ack_0, ack => convTransposeD_CP_7576_elements(19)); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	2 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (12) 
      -- CP-element group 20: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/LOAD_padding_2833_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/LOAD_padding_2833_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/LOAD_padding_2833_Update/word_access_complete/$exit
      -- CP-element group 20: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/LOAD_padding_2833_Update/word_access_complete/word_0/$exit
      -- CP-element group 20: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/LOAD_padding_2833_Update/word_access_complete/word_0/ca
      -- CP-element group 20: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/LOAD_padding_2833_Update/LOAD_padding_2833_Merge/$entry
      -- CP-element group 20: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/LOAD_padding_2833_Update/LOAD_padding_2833_Merge/$exit
      -- CP-element group 20: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/LOAD_padding_2833_Update/LOAD_padding_2833_Merge/merge_req
      -- CP-element group 20: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/LOAD_padding_2833_Update/LOAD_padding_2833_Merge/merge_ack
      -- CP-element group 20: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/type_cast_2837_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/type_cast_2837_Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/type_cast_2837_Sample/rr
      -- 
    ca_7963_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_padding_2833_load_0_ack_1, ack => convTransposeD_CP_7576_elements(20)); -- 
    rr_7976_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7976_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(20), ack => type_cast_2837_inst_req_0); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/type_cast_2837_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/type_cast_2837_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/type_cast_2837_Sample/ra
      -- 
    ra_7977_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2837_inst_ack_0, ack => convTransposeD_CP_7576_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	2 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	33 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/type_cast_2837_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/type_cast_2837_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/type_cast_2837_Update/ca
      -- 
    ca_7982_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2837_inst_ack_1, ack => convTransposeD_CP_7576_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	2 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (5) 
      -- CP-element group 23: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2847_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2847_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2847_Sample/word_access_start/$exit
      -- CP-element group 23: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2847_Sample/word_access_start/word_0/$exit
      -- CP-element group 23: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2847_Sample/word_access_start/word_0/ra
      -- 
    ra_8016_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2847_load_0_ack_0, ack => convTransposeD_CP_7576_elements(23)); -- 
    -- CP-element group 24:  transition  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	2 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (12) 
      -- CP-element group 24: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2847_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2847_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2847_Update/word_access_complete/$exit
      -- CP-element group 24: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2847_Update/word_access_complete/word_0/$exit
      -- CP-element group 24: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2847_Update/word_access_complete/word_0/ca
      -- CP-element group 24: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2847_Update/ptr_deref_2847_Merge/$entry
      -- CP-element group 24: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2847_Update/ptr_deref_2847_Merge/$exit
      -- CP-element group 24: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2847_Update/ptr_deref_2847_Merge/merge_req
      -- CP-element group 24: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2847_Update/ptr_deref_2847_Merge/merge_ack
      -- CP-element group 24: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/type_cast_2851_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/type_cast_2851_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/type_cast_2851_Sample/rr
      -- 
    ca_8027_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2847_load_0_ack_1, ack => convTransposeD_CP_7576_elements(24)); -- 
    rr_8040_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8040_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(24), ack => type_cast_2851_inst_req_0); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/type_cast_2851_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/type_cast_2851_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/type_cast_2851_Sample/ra
      -- 
    ra_8041_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2851_inst_ack_0, ack => convTransposeD_CP_7576_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	2 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	33 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/type_cast_2851_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/type_cast_2851_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/type_cast_2851_Update/ca
      -- 
    ca_8046_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2851_inst_ack_1, ack => convTransposeD_CP_7576_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	2 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (5) 
      -- CP-element group 27: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2863_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2863_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2863_Sample/word_access_start/$exit
      -- CP-element group 27: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2863_Sample/word_access_start/word_0/$exit
      -- CP-element group 27: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2863_Sample/word_access_start/word_0/ra
      -- 
    ra_8080_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2863_load_0_ack_0, ack => convTransposeD_CP_7576_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	2 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	33 
    -- CP-element group 28:  members (9) 
      -- CP-element group 28: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2863_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2863_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2863_Update/word_access_complete/$exit
      -- CP-element group 28: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2863_Update/word_access_complete/word_0/$exit
      -- CP-element group 28: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2863_Update/word_access_complete/word_0/ca
      -- CP-element group 28: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2863_Update/ptr_deref_2863_Merge/$entry
      -- CP-element group 28: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2863_Update/ptr_deref_2863_Merge/$exit
      -- CP-element group 28: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2863_Update/ptr_deref_2863_Merge/merge_req
      -- CP-element group 28: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2863_Update/ptr_deref_2863_Merge/merge_ack
      -- 
    ca_8091_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2863_load_0_ack_1, ack => convTransposeD_CP_7576_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	2 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (5) 
      -- CP-element group 29: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2875_Sample/word_access_start/word_0/$exit
      -- CP-element group 29: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2875_Sample/word_access_start/$exit
      -- CP-element group 29: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2875_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2875_Sample/word_access_start/word_0/ra
      -- CP-element group 29: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2875_sample_completed_
      -- 
    ra_8130_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2875_load_0_ack_0, ack => convTransposeD_CP_7576_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	2 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	33 
    -- CP-element group 30:  members (9) 
      -- CP-element group 30: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2875_Update/word_access_complete/$exit
      -- CP-element group 30: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2875_Update/ptr_deref_2875_Merge/$entry
      -- CP-element group 30: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2875_Update/word_access_complete/word_0/ca
      -- CP-element group 30: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2875_Update/word_access_complete/word_0/$exit
      -- CP-element group 30: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2875_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2875_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2875_Update/ptr_deref_2875_Merge/merge_ack
      -- CP-element group 30: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2875_Update/ptr_deref_2875_Merge/merge_req
      -- CP-element group 30: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2875_Update/ptr_deref_2875_Merge/$exit
      -- 
    ca_8141_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2875_load_0_ack_1, ack => convTransposeD_CP_7576_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	2 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (5) 
      -- CP-element group 31: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2887_Sample/$exit
      -- CP-element group 31: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2887_Sample/word_access_start/word_0/ra
      -- CP-element group 31: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2887_sample_completed_
      -- CP-element group 31: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2887_Sample/word_access_start/$exit
      -- CP-element group 31: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2887_Sample/word_access_start/word_0/$exit
      -- 
    ra_8180_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2887_load_0_ack_0, ack => convTransposeD_CP_7576_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	2 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (9) 
      -- CP-element group 32: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2887_Update/word_access_complete/$exit
      -- CP-element group 32: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2887_Update/$exit
      -- CP-element group 32: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2887_Update/ptr_deref_2887_Merge/merge_ack
      -- CP-element group 32: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2887_update_completed_
      -- CP-element group 32: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2887_Update/ptr_deref_2887_Merge/$exit
      -- CP-element group 32: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2887_Update/ptr_deref_2887_Merge/merge_req
      -- CP-element group 32: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2887_Update/word_access_complete/word_0/ca
      -- CP-element group 32: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2887_Update/ptr_deref_2887_Merge/$entry
      -- CP-element group 32: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/ptr_deref_2887_Update/word_access_complete/word_0/$exit
      -- 
    ca_8191_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2887_load_0_ack_1, ack => convTransposeD_CP_7576_elements(32)); -- 
    -- CP-element group 33:  join  fork  transition  place  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	30 
    -- CP-element group 33: 	22 
    -- CP-element group 33: 	28 
    -- CP-element group 33: 	16 
    -- CP-element group 33: 	26 
    -- CP-element group 33: 	32 
    -- CP-element group 33: 	18 
    -- CP-element group 33: 	6 
    -- CP-element group 33: 	10 
    -- CP-element group 33: 	12 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	75 
    -- CP-element group 33: 	76 
    -- CP-element group 33: 	78 
    -- CP-element group 33: 	79 
    -- CP-element group 33:  members (20) 
      -- CP-element group 33: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888__exit__
      -- CP-element group 33: 	 branch_block_stmt_2745/entry_whilex_xbodyx_xouter
      -- CP-element group 33: 	 branch_block_stmt_2745/assign_stmt_2757_to_assign_stmt_2888/$exit
      -- CP-element group 33: 	 branch_block_stmt_2745/entry_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 33: 	 branch_block_stmt_2745/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2891/$entry
      -- CP-element group 33: 	 branch_block_stmt_2745/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2891/phi_stmt_2891_sources/$entry
      -- CP-element group 33: 	 branch_block_stmt_2745/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2891/phi_stmt_2891_sources/type_cast_2894/$entry
      -- CP-element group 33: 	 branch_block_stmt_2745/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2891/phi_stmt_2891_sources/type_cast_2894/SplitProtocol/$entry
      -- CP-element group 33: 	 branch_block_stmt_2745/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2891/phi_stmt_2891_sources/type_cast_2894/SplitProtocol/Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_2745/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2891/phi_stmt_2891_sources/type_cast_2894/SplitProtocol/Sample/rr
      -- CP-element group 33: 	 branch_block_stmt_2745/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2891/phi_stmt_2891_sources/type_cast_2894/SplitProtocol/Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_2745/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2891/phi_stmt_2891_sources/type_cast_2894/SplitProtocol/Update/cr
      -- CP-element group 33: 	 branch_block_stmt_2745/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2897/$entry
      -- CP-element group 33: 	 branch_block_stmt_2745/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2897/phi_stmt_2897_sources/$entry
      -- CP-element group 33: 	 branch_block_stmt_2745/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2897/phi_stmt_2897_sources/type_cast_2900/$entry
      -- CP-element group 33: 	 branch_block_stmt_2745/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2897/phi_stmt_2897_sources/type_cast_2900/SplitProtocol/$entry
      -- CP-element group 33: 	 branch_block_stmt_2745/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2897/phi_stmt_2897_sources/type_cast_2900/SplitProtocol/Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_2745/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2897/phi_stmt_2897_sources/type_cast_2900/SplitProtocol/Sample/rr
      -- CP-element group 33: 	 branch_block_stmt_2745/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2897/phi_stmt_2897_sources/type_cast_2900/SplitProtocol/Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_2745/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2897/phi_stmt_2897_sources/type_cast_2900/SplitProtocol/Update/cr
      -- 
    rr_8625_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8625_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(33), ack => type_cast_2894_inst_req_0); -- 
    cr_8630_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8630_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(33), ack => type_cast_2894_inst_req_1); -- 
    rr_8648_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8648_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(33), ack => type_cast_2900_inst_req_0); -- 
    cr_8653_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8653_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(33), ack => type_cast_2900_inst_req_1); -- 
    convTransposeD_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= convTransposeD_CP_7576_elements(30) & convTransposeD_CP_7576_elements(22) & convTransposeD_CP_7576_elements(28) & convTransposeD_CP_7576_elements(16) & convTransposeD_CP_7576_elements(26) & convTransposeD_CP_7576_elements(32) & convTransposeD_CP_7576_elements(18) & convTransposeD_CP_7576_elements(6) & convTransposeD_CP_7576_elements(10) & convTransposeD_CP_7576_elements(12);
      gj_convTransposeD_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7576_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	92 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_2745/assign_stmt_2908_to_assign_stmt_3015/type_cast_2907_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_2745/assign_stmt_2908_to_assign_stmt_3015/type_cast_2907_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_2745/assign_stmt_2908_to_assign_stmt_3015/type_cast_2907_Sample/ra
      -- 
    ra_8208_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2907_inst_ack_0, ack => convTransposeD_CP_7576_elements(34)); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	92 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	38 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_2745/assign_stmt_2908_to_assign_stmt_3015/type_cast_2907_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_2745/assign_stmt_2908_to_assign_stmt_3015/type_cast_2907_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_2745/assign_stmt_2908_to_assign_stmt_3015/type_cast_2907_Update/ca
      -- 
    ca_8213_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2907_inst_ack_1, ack => convTransposeD_CP_7576_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	92 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_2745/assign_stmt_2908_to_assign_stmt_3015/type_cast_2912_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_2745/assign_stmt_2908_to_assign_stmt_3015/type_cast_2912_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_2745/assign_stmt_2908_to_assign_stmt_3015/type_cast_2912_Sample/ra
      -- 
    ra_8222_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2912_inst_ack_0, ack => convTransposeD_CP_7576_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	92 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_2745/assign_stmt_2908_to_assign_stmt_3015/type_cast_2912_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_2745/assign_stmt_2908_to_assign_stmt_3015/type_cast_2912_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_2745/assign_stmt_2908_to_assign_stmt_3015/type_cast_2912_Update/ca
      -- 
    ca_8227_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2912_inst_ack_1, ack => convTransposeD_CP_7576_elements(37)); -- 
    -- CP-element group 38:  join  transition  place  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: 	35 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	96 
    -- CP-element group 38:  members (6) 
      -- CP-element group 38: 	 branch_block_stmt_2745/assign_stmt_2908_to_assign_stmt_3015__exit__
      -- CP-element group 38: 	 branch_block_stmt_2745/whilex_xbodyx_xouter_whilex_xbody
      -- CP-element group 38: 	 branch_block_stmt_2745/assign_stmt_2908_to_assign_stmt_3015/$exit
      -- CP-element group 38: 	 branch_block_stmt_2745/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$entry
      -- CP-element group 38: 	 branch_block_stmt_2745/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_3018/$entry
      -- CP-element group 38: 	 branch_block_stmt_2745/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_3018/phi_stmt_3018_sources/$entry
      -- 
    convTransposeD_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7576_elements(37) & convTransposeD_CP_7576_elements(35);
      gj_convTransposeD_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7576_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	98 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/type_cast_3034_Sample/ra
      -- CP-element group 39: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/type_cast_3034_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/type_cast_3034_sample_completed_
      -- 
    ra_8239_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3034_inst_ack_0, ack => convTransposeD_CP_7576_elements(39)); -- 
    -- CP-element group 40:  fork  transition  input  output  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	98 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	49 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (9) 
      -- CP-element group 40: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/type_cast_3064_sample_start_
      -- CP-element group 40: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/type_cast_3064_Sample/rr
      -- CP-element group 40: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/type_cast_3064_Sample/$entry
      -- CP-element group 40: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/type_cast_3034_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/type_cast_3034_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/type_cast_3034_Update/ca
      -- CP-element group 40: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/type_cast_3095_sample_start_
      -- CP-element group 40: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/type_cast_3095_Sample/$entry
      -- CP-element group 40: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/type_cast_3095_Sample/rr
      -- 
    ca_8244_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3034_inst_ack_1, ack => convTransposeD_CP_7576_elements(40)); -- 
    rr_8362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(40), ack => type_cast_3095_inst_req_0); -- 
    rr_8252_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8252_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(40), ack => type_cast_3064_inst_req_0); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/type_cast_3064_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/type_cast_3064_Sample/ra
      -- CP-element group 41: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/type_cast_3064_Sample/$exit
      -- 
    ra_8253_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3064_inst_ack_0, ack => convTransposeD_CP_7576_elements(41)); -- 
    -- CP-element group 42:  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	98 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (16) 
      -- CP-element group 42: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/type_cast_3064_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/array_obj_ref_3070_index_resize_1/$entry
      -- CP-element group 42: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/array_obj_ref_3070_index_scale_1/$entry
      -- CP-element group 42: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/array_obj_ref_3070_index_resized_1
      -- CP-element group 42: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/array_obj_ref_3070_index_scaled_1
      -- CP-element group 42: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/array_obj_ref_3070_final_index_sum_regn_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/array_obj_ref_3070_index_resize_1/$exit
      -- CP-element group 42: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/array_obj_ref_3070_index_scale_1/$exit
      -- CP-element group 42: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/array_obj_ref_3070_final_index_sum_regn_Sample/req
      -- CP-element group 42: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/array_obj_ref_3070_index_scale_1/scale_rename_ack
      -- CP-element group 42: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/type_cast_3064_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/array_obj_ref_3070_index_resize_1/index_resize_req
      -- CP-element group 42: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/array_obj_ref_3070_index_resize_1/index_resize_ack
      -- CP-element group 42: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/type_cast_3064_Update/ca
      -- CP-element group 42: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/array_obj_ref_3070_index_scale_1/scale_rename_req
      -- CP-element group 42: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/array_obj_ref_3070_index_computed_1
      -- 
    ca_8258_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3064_inst_ack_1, ack => convTransposeD_CP_7576_elements(42)); -- 
    req_8283_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8283_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(42), ack => array_obj_ref_3070_index_offset_req_0); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	60 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/array_obj_ref_3070_final_index_sum_regn_Sample/ack
      -- CP-element group 43: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/array_obj_ref_3070_final_index_sum_regn_sample_complete
      -- CP-element group 43: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/array_obj_ref_3070_final_index_sum_regn_Sample/$exit
      -- 
    ack_8284_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3070_index_offset_ack_0, ack => convTransposeD_CP_7576_elements(43)); -- 
    -- CP-element group 44:  transition  input  output  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	98 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (11) 
      -- CP-element group 44: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/array_obj_ref_3070_final_index_sum_regn_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/array_obj_ref_3070_root_address_calculated
      -- CP-element group 44: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/array_obj_ref_3070_offset_calculated
      -- CP-element group 44: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/addr_of_3071_sample_start_
      -- CP-element group 44: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/array_obj_ref_3070_base_plus_offset/$entry
      -- CP-element group 44: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/array_obj_ref_3070_base_plus_offset/$exit
      -- CP-element group 44: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/array_obj_ref_3070_base_plus_offset/sum_rename_req
      -- CP-element group 44: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/array_obj_ref_3070_base_plus_offset/sum_rename_ack
      -- CP-element group 44: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/addr_of_3071_request/$entry
      -- CP-element group 44: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/addr_of_3071_request/req
      -- CP-element group 44: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/array_obj_ref_3070_final_index_sum_regn_Update/ack
      -- 
    ack_8289_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3070_index_offset_ack_1, ack => convTransposeD_CP_7576_elements(44)); -- 
    req_8298_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8298_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(44), ack => addr_of_3071_final_reg_req_0); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	44 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/addr_of_3071_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/addr_of_3071_request/$exit
      -- CP-element group 45: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/addr_of_3071_request/ack
      -- 
    ack_8299_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3071_final_reg_ack_0, ack => convTransposeD_CP_7576_elements(45)); -- 
    -- CP-element group 46:  join  fork  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	98 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (24) 
      -- CP-element group 46: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3075_base_addr_resize/base_resize_ack
      -- CP-element group 46: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3075_word_address_calculated
      -- CP-element group 46: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3075_base_plus_offset/$entry
      -- CP-element group 46: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3075_base_plus_offset/$exit
      -- CP-element group 46: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3075_base_addr_resize/base_resize_req
      -- CP-element group 46: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/addr_of_3071_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/addr_of_3071_complete/ack
      -- CP-element group 46: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3075_base_plus_offset/sum_rename_req
      -- CP-element group 46: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3075_base_address_resized
      -- CP-element group 46: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3075_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3075_Sample/word_access_start/$entry
      -- CP-element group 46: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3075_base_address_calculated
      -- CP-element group 46: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3075_base_plus_offset/sum_rename_ack
      -- CP-element group 46: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3075_word_addrgen/$entry
      -- CP-element group 46: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3075_word_addrgen/$exit
      -- CP-element group 46: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3075_word_addrgen/root_register_req
      -- CP-element group 46: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3075_word_addrgen/root_register_ack
      -- CP-element group 46: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/addr_of_3071_complete/$exit
      -- CP-element group 46: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3075_base_addr_resize/$entry
      -- CP-element group 46: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3075_base_addr_resize/$exit
      -- CP-element group 46: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3075_root_address_calculated
      -- CP-element group 46: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3075_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3075_Sample/word_access_start/word_0/$entry
      -- CP-element group 46: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3075_Sample/word_access_start/word_0/rr
      -- 
    ack_8304_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3071_final_reg_ack_1, ack => convTransposeD_CP_7576_elements(46)); -- 
    rr_8337_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8337_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(46), ack => ptr_deref_3075_load_0_req_0); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (5) 
      -- CP-element group 47: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3075_Sample/word_access_start/$exit
      -- CP-element group 47: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3075_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3075_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3075_Sample/word_access_start/word_0/$exit
      -- CP-element group 47: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3075_Sample/word_access_start/word_0/ra
      -- 
    ra_8338_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3075_load_0_ack_0, ack => convTransposeD_CP_7576_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	98 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	55 
    -- CP-element group 48:  members (9) 
      -- CP-element group 48: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3075_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3075_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3075_Update/word_access_complete/$exit
      -- CP-element group 48: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3075_Update/word_access_complete/word_0/$exit
      -- CP-element group 48: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3075_Update/word_access_complete/word_0/ca
      -- CP-element group 48: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3075_Update/ptr_deref_3075_Merge/$entry
      -- CP-element group 48: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3075_Update/ptr_deref_3075_Merge/$exit
      -- CP-element group 48: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3075_Update/ptr_deref_3075_Merge/merge_req
      -- CP-element group 48: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3075_Update/ptr_deref_3075_Merge/merge_ack
      -- 
    ca_8349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3075_load_0_ack_1, ack => convTransposeD_CP_7576_elements(48)); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	40 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/type_cast_3095_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/type_cast_3095_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/type_cast_3095_Sample/ra
      -- 
    ra_8363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3095_inst_ack_0, ack => convTransposeD_CP_7576_elements(49)); -- 
    -- CP-element group 50:  transition  input  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	98 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (16) 
      -- CP-element group 50: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/type_cast_3095_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/type_cast_3095_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/type_cast_3095_Update/ca
      -- CP-element group 50: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/array_obj_ref_3101_index_resized_1
      -- CP-element group 50: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/array_obj_ref_3101_index_scaled_1
      -- CP-element group 50: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/array_obj_ref_3101_index_computed_1
      -- CP-element group 50: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/array_obj_ref_3101_index_resize_1/$entry
      -- CP-element group 50: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/array_obj_ref_3101_index_resize_1/$exit
      -- CP-element group 50: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/array_obj_ref_3101_index_resize_1/index_resize_req
      -- CP-element group 50: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/array_obj_ref_3101_index_resize_1/index_resize_ack
      -- CP-element group 50: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/array_obj_ref_3101_index_scale_1/$entry
      -- CP-element group 50: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/array_obj_ref_3101_index_scale_1/$exit
      -- CP-element group 50: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/array_obj_ref_3101_index_scale_1/scale_rename_req
      -- CP-element group 50: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/array_obj_ref_3101_index_scale_1/scale_rename_ack
      -- CP-element group 50: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/array_obj_ref_3101_final_index_sum_regn_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/array_obj_ref_3101_final_index_sum_regn_Sample/req
      -- 
    ca_8368_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3095_inst_ack_1, ack => convTransposeD_CP_7576_elements(50)); -- 
    req_8393_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8393_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(50), ack => array_obj_ref_3101_index_offset_req_0); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	60 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/array_obj_ref_3101_final_index_sum_regn_sample_complete
      -- CP-element group 51: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/array_obj_ref_3101_final_index_sum_regn_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/array_obj_ref_3101_final_index_sum_regn_Sample/ack
      -- 
    ack_8394_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3101_index_offset_ack_0, ack => convTransposeD_CP_7576_elements(51)); -- 
    -- CP-element group 52:  transition  input  output  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	98 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	53 
    -- CP-element group 52:  members (11) 
      -- CP-element group 52: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/addr_of_3102_request/$entry
      -- CP-element group 52: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/addr_of_3102_sample_start_
      -- CP-element group 52: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/array_obj_ref_3101_root_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/array_obj_ref_3101_offset_calculated
      -- CP-element group 52: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/array_obj_ref_3101_final_index_sum_regn_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/array_obj_ref_3101_final_index_sum_regn_Update/ack
      -- CP-element group 52: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/array_obj_ref_3101_base_plus_offset/$entry
      -- CP-element group 52: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/array_obj_ref_3101_base_plus_offset/$exit
      -- CP-element group 52: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/array_obj_ref_3101_base_plus_offset/sum_rename_req
      -- CP-element group 52: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/array_obj_ref_3101_base_plus_offset/sum_rename_ack
      -- CP-element group 52: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/addr_of_3102_request/req
      -- 
    ack_8399_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3101_index_offset_ack_1, ack => convTransposeD_CP_7576_elements(52)); -- 
    req_8408_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8408_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(52), ack => addr_of_3102_final_reg_req_0); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	52 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/addr_of_3102_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/addr_of_3102_request/$exit
      -- CP-element group 53: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/addr_of_3102_request/ack
      -- 
    ack_8409_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3102_final_reg_ack_0, ack => convTransposeD_CP_7576_elements(53)); -- 
    -- CP-element group 54:  fork  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	98 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54:  members (19) 
      -- CP-element group 54: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/addr_of_3102_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/addr_of_3102_complete/$exit
      -- CP-element group 54: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/addr_of_3102_complete/ack
      -- CP-element group 54: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3105_base_address_calculated
      -- CP-element group 54: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3105_word_address_calculated
      -- CP-element group 54: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3105_root_address_calculated
      -- CP-element group 54: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3105_base_address_resized
      -- CP-element group 54: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3105_base_addr_resize/$entry
      -- CP-element group 54: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3105_base_addr_resize/$exit
      -- CP-element group 54: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3105_base_addr_resize/base_resize_req
      -- CP-element group 54: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3105_base_addr_resize/base_resize_ack
      -- CP-element group 54: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3105_base_plus_offset/$entry
      -- CP-element group 54: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3105_base_plus_offset/$exit
      -- CP-element group 54: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3105_base_plus_offset/sum_rename_req
      -- CP-element group 54: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3105_base_plus_offset/sum_rename_ack
      -- CP-element group 54: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3105_word_addrgen/$entry
      -- CP-element group 54: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3105_word_addrgen/$exit
      -- CP-element group 54: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3105_word_addrgen/root_register_req
      -- CP-element group 54: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3105_word_addrgen/root_register_ack
      -- 
    ack_8414_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3102_final_reg_ack_1, ack => convTransposeD_CP_7576_elements(54)); -- 
    -- CP-element group 55:  join  transition  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	48 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (9) 
      -- CP-element group 55: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3105_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3105_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3105_Sample/ptr_deref_3105_Split/$entry
      -- CP-element group 55: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3105_Sample/ptr_deref_3105_Split/$exit
      -- CP-element group 55: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3105_Sample/ptr_deref_3105_Split/split_req
      -- CP-element group 55: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3105_Sample/ptr_deref_3105_Split/split_ack
      -- CP-element group 55: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3105_Sample/word_access_start/$entry
      -- CP-element group 55: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3105_Sample/word_access_start/word_0/$entry
      -- CP-element group 55: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3105_Sample/word_access_start/word_0/rr
      -- 
    rr_8452_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8452_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(55), ack => ptr_deref_3105_store_0_req_0); -- 
    convTransposeD_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7576_elements(48) & convTransposeD_CP_7576_elements(54);
      gj_convTransposeD_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7576_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (5) 
      -- CP-element group 56: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3105_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3105_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3105_Sample/word_access_start/$exit
      -- CP-element group 56: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3105_Sample/word_access_start/word_0/$exit
      -- CP-element group 56: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3105_Sample/word_access_start/word_0/ra
      -- 
    ra_8453_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3105_store_0_ack_0, ack => convTransposeD_CP_7576_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	98 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	60 
    -- CP-element group 57:  members (5) 
      -- CP-element group 57: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3105_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3105_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3105_Update/word_access_complete/$exit
      -- CP-element group 57: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3105_Update/word_access_complete/word_0/$exit
      -- CP-element group 57: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3105_Update/word_access_complete/word_0/ca
      -- 
    ca_8464_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3105_store_0_ack_1, ack => convTransposeD_CP_7576_elements(57)); -- 
    -- CP-element group 58:  transition  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	98 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/type_cast_3111_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/type_cast_3111_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/type_cast_3111_Sample/ra
      -- 
    ra_8473_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3111_inst_ack_0, ack => convTransposeD_CP_7576_elements(58)); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	98 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/type_cast_3111_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/type_cast_3111_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/type_cast_3111_Update/ca
      -- 
    ca_8478_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3111_inst_ack_1, ack => convTransposeD_CP_7576_elements(59)); -- 
    -- CP-element group 60:  branch  join  transition  place  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	57 
    -- CP-element group 60: 	51 
    -- CP-element group 60: 	43 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60: 	62 
    -- CP-element group 60:  members (10) 
      -- CP-element group 60: 	 branch_block_stmt_2745/R_cmp_3125_place
      -- CP-element group 60: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123__exit__
      -- CP-element group 60: 	 branch_block_stmt_2745/if_stmt_3124__entry__
      -- CP-element group 60: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/$exit
      -- CP-element group 60: 	 branch_block_stmt_2745/if_stmt_3124_dead_link/$entry
      -- CP-element group 60: 	 branch_block_stmt_2745/if_stmt_3124_eval_test/$entry
      -- CP-element group 60: 	 branch_block_stmt_2745/if_stmt_3124_eval_test/$exit
      -- CP-element group 60: 	 branch_block_stmt_2745/if_stmt_3124_eval_test/branch_req
      -- CP-element group 60: 	 branch_block_stmt_2745/if_stmt_3124_if_link/$entry
      -- CP-element group 60: 	 branch_block_stmt_2745/if_stmt_3124_else_link/$entry
      -- 
    branch_req_8486_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_8486_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(60), ack => if_stmt_3124_branch_req_0); -- 
    convTransposeD_cp_element_group_60: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_60"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeD_CP_7576_elements(57) & convTransposeD_CP_7576_elements(51) & convTransposeD_CP_7576_elements(43) & convTransposeD_CP_7576_elements(59);
      gj_convTransposeD_cp_element_group_60 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7576_elements(60), clk => clk, reset => reset); --
    end block;
    -- CP-element group 61:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	93 
    -- CP-element group 61: 	94 
    -- CP-element group 61:  members (24) 
      -- CP-element group 61: 	 branch_block_stmt_2745/whilex_xbody_ifx_xthen
      -- CP-element group 61: 	 branch_block_stmt_2745/merge_stmt_3130__exit__
      -- CP-element group 61: 	 branch_block_stmt_2745/assign_stmt_3136__entry__
      -- CP-element group 61: 	 branch_block_stmt_2745/assign_stmt_3136__exit__
      -- CP-element group 61: 	 branch_block_stmt_2745/ifx_xthen_whilex_xbody
      -- CP-element group 61: 	 branch_block_stmt_2745/if_stmt_3124_if_link/$exit
      -- CP-element group 61: 	 branch_block_stmt_2745/if_stmt_3124_if_link/if_choice_transition
      -- CP-element group 61: 	 branch_block_stmt_2745/assign_stmt_3136/$entry
      -- CP-element group 61: 	 branch_block_stmt_2745/assign_stmt_3136/$exit
      -- CP-element group 61: 	 branch_block_stmt_2745/ifx_xthen_whilex_xbody_PhiReq/$entry
      -- CP-element group 61: 	 branch_block_stmt_2745/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3018/$entry
      -- CP-element group 61: 	 branch_block_stmt_2745/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3018/phi_stmt_3018_sources/$entry
      -- CP-element group 61: 	 branch_block_stmt_2745/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3018/phi_stmt_3018_sources/type_cast_3024/$entry
      -- CP-element group 61: 	 branch_block_stmt_2745/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3018/phi_stmt_3018_sources/type_cast_3024/SplitProtocol/$entry
      -- CP-element group 61: 	 branch_block_stmt_2745/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3018/phi_stmt_3018_sources/type_cast_3024/SplitProtocol/Sample/$entry
      -- CP-element group 61: 	 branch_block_stmt_2745/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3018/phi_stmt_3018_sources/type_cast_3024/SplitProtocol/Sample/rr
      -- CP-element group 61: 	 branch_block_stmt_2745/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3018/phi_stmt_3018_sources/type_cast_3024/SplitProtocol/Update/$entry
      -- CP-element group 61: 	 branch_block_stmt_2745/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3018/phi_stmt_3018_sources/type_cast_3024/SplitProtocol/Update/cr
      -- CP-element group 61: 	 branch_block_stmt_2745/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 61: 	 branch_block_stmt_2745/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 61: 	 branch_block_stmt_2745/merge_stmt_3130_PhiReqMerge
      -- CP-element group 61: 	 branch_block_stmt_2745/merge_stmt_3130_PhiAck/$entry
      -- CP-element group 61: 	 branch_block_stmt_2745/merge_stmt_3130_PhiAck/$exit
      -- CP-element group 61: 	 branch_block_stmt_2745/merge_stmt_3130_PhiAck/dummy
      -- 
    if_choice_transition_8491_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3124_branch_ack_1, ack => convTransposeD_CP_7576_elements(61)); -- 
    rr_8729_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8729_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(61), ack => type_cast_3024_inst_req_0); -- 
    cr_8734_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8734_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(61), ack => type_cast_3024_inst_req_1); -- 
    -- CP-element group 62:  fork  transition  place  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	60 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62: 	64 
    -- CP-element group 62:  members (18) 
      -- CP-element group 62: 	 branch_block_stmt_2745/whilex_xbody_ifx_xelse
      -- CP-element group 62: 	 branch_block_stmt_2745/merge_stmt_3138__exit__
      -- CP-element group 62: 	 branch_block_stmt_2745/assign_stmt_3144_to_assign_stmt_3154__entry__
      -- CP-element group 62: 	 branch_block_stmt_2745/if_stmt_3124_else_link/$exit
      -- CP-element group 62: 	 branch_block_stmt_2745/if_stmt_3124_else_link/else_choice_transition
      -- CP-element group 62: 	 branch_block_stmt_2745/assign_stmt_3144_to_assign_stmt_3154/$entry
      -- CP-element group 62: 	 branch_block_stmt_2745/assign_stmt_3144_to_assign_stmt_3154/type_cast_3148_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_2745/assign_stmt_3144_to_assign_stmt_3154/type_cast_3148_update_start_
      -- CP-element group 62: 	 branch_block_stmt_2745/assign_stmt_3144_to_assign_stmt_3154/type_cast_3148_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_2745/assign_stmt_3144_to_assign_stmt_3154/type_cast_3148_Sample/rr
      -- CP-element group 62: 	 branch_block_stmt_2745/assign_stmt_3144_to_assign_stmt_3154/type_cast_3148_Update/$entry
      -- CP-element group 62: 	 branch_block_stmt_2745/assign_stmt_3144_to_assign_stmt_3154/type_cast_3148_Update/cr
      -- CP-element group 62: 	 branch_block_stmt_2745/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 62: 	 branch_block_stmt_2745/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 62: 	 branch_block_stmt_2745/merge_stmt_3138_PhiReqMerge
      -- CP-element group 62: 	 branch_block_stmt_2745/merge_stmt_3138_PhiAck/$entry
      -- CP-element group 62: 	 branch_block_stmt_2745/merge_stmt_3138_PhiAck/$exit
      -- CP-element group 62: 	 branch_block_stmt_2745/merge_stmt_3138_PhiAck/dummy
      -- 
    else_choice_transition_8495_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3124_branch_ack_0, ack => convTransposeD_CP_7576_elements(62)); -- 
    rr_8511_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8511_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(62), ack => type_cast_3148_inst_req_0); -- 
    cr_8516_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8516_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(62), ack => type_cast_3148_inst_req_1); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_2745/assign_stmt_3144_to_assign_stmt_3154/type_cast_3148_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_2745/assign_stmt_3144_to_assign_stmt_3154/type_cast_3148_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_2745/assign_stmt_3144_to_assign_stmt_3154/type_cast_3148_Sample/ra
      -- 
    ra_8512_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3148_inst_ack_0, ack => convTransposeD_CP_7576_elements(63)); -- 
    -- CP-element group 64:  branch  transition  place  input  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	62 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64: 	66 
    -- CP-element group 64:  members (13) 
      -- CP-element group 64: 	 branch_block_stmt_2745/R_cmp81_3156_place
      -- CP-element group 64: 	 branch_block_stmt_2745/assign_stmt_3144_to_assign_stmt_3154__exit__
      -- CP-element group 64: 	 branch_block_stmt_2745/if_stmt_3155__entry__
      -- CP-element group 64: 	 branch_block_stmt_2745/assign_stmt_3144_to_assign_stmt_3154/$exit
      -- CP-element group 64: 	 branch_block_stmt_2745/assign_stmt_3144_to_assign_stmt_3154/type_cast_3148_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_2745/assign_stmt_3144_to_assign_stmt_3154/type_cast_3148_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_2745/assign_stmt_3144_to_assign_stmt_3154/type_cast_3148_Update/ca
      -- CP-element group 64: 	 branch_block_stmt_2745/if_stmt_3155_dead_link/$entry
      -- CP-element group 64: 	 branch_block_stmt_2745/if_stmt_3155_eval_test/$entry
      -- CP-element group 64: 	 branch_block_stmt_2745/if_stmt_3155_eval_test/$exit
      -- CP-element group 64: 	 branch_block_stmt_2745/if_stmt_3155_eval_test/branch_req
      -- CP-element group 64: 	 branch_block_stmt_2745/if_stmt_3155_if_link/$entry
      -- CP-element group 64: 	 branch_block_stmt_2745/if_stmt_3155_else_link/$entry
      -- 
    ca_8517_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3148_inst_ack_1, ack => convTransposeD_CP_7576_elements(64)); -- 
    branch_req_8525_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_8525_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(64), ack => if_stmt_3155_branch_req_0); -- 
    -- CP-element group 65:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	67 
    -- CP-element group 65: 	68 
    -- CP-element group 65:  members (18) 
      -- CP-element group 65: 	 branch_block_stmt_2745/ifx_xelse_ifx_xthen83
      -- CP-element group 65: 	 branch_block_stmt_2745/merge_stmt_3161__exit__
      -- CP-element group 65: 	 branch_block_stmt_2745/assign_stmt_3167_to_assign_stmt_3177__entry__
      -- CP-element group 65: 	 branch_block_stmt_2745/if_stmt_3155_if_link/$exit
      -- CP-element group 65: 	 branch_block_stmt_2745/if_stmt_3155_if_link/if_choice_transition
      -- CP-element group 65: 	 branch_block_stmt_2745/assign_stmt_3167_to_assign_stmt_3177/$entry
      -- CP-element group 65: 	 branch_block_stmt_2745/assign_stmt_3167_to_assign_stmt_3177/type_cast_3176_sample_start_
      -- CP-element group 65: 	 branch_block_stmt_2745/assign_stmt_3167_to_assign_stmt_3177/type_cast_3176_update_start_
      -- CP-element group 65: 	 branch_block_stmt_2745/assign_stmt_3167_to_assign_stmt_3177/type_cast_3176_Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_2745/assign_stmt_3167_to_assign_stmt_3177/type_cast_3176_Sample/rr
      -- CP-element group 65: 	 branch_block_stmt_2745/assign_stmt_3167_to_assign_stmt_3177/type_cast_3176_Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_2745/assign_stmt_3167_to_assign_stmt_3177/type_cast_3176_Update/cr
      -- CP-element group 65: 	 branch_block_stmt_2745/ifx_xelse_ifx_xthen83_PhiReq/$entry
      -- CP-element group 65: 	 branch_block_stmt_2745/ifx_xelse_ifx_xthen83_PhiReq/$exit
      -- CP-element group 65: 	 branch_block_stmt_2745/merge_stmt_3161_PhiReqMerge
      -- CP-element group 65: 	 branch_block_stmt_2745/merge_stmt_3161_PhiAck/$entry
      -- CP-element group 65: 	 branch_block_stmt_2745/merge_stmt_3161_PhiAck/$exit
      -- CP-element group 65: 	 branch_block_stmt_2745/merge_stmt_3161_PhiAck/dummy
      -- 
    if_choice_transition_8530_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3155_branch_ack_1, ack => convTransposeD_CP_7576_elements(65)); -- 
    rr_8547_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8547_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(65), ack => type_cast_3176_inst_req_0); -- 
    cr_8552_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8552_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(65), ack => type_cast_3176_inst_req_1); -- 
    -- CP-element group 66:  fork  transition  place  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	64 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	103 
    -- CP-element group 66: 	99 
    -- CP-element group 66: 	100 
    -- CP-element group 66: 	102 
    -- CP-element group 66:  members (20) 
      -- CP-element group 66: 	 branch_block_stmt_2745/ifx_xelse_ifx_xend
      -- CP-element group 66: 	 branch_block_stmt_2745/if_stmt_3155_else_link/$exit
      -- CP-element group 66: 	 branch_block_stmt_2745/if_stmt_3155_else_link/else_choice_transition
      -- CP-element group 66: 	 branch_block_stmt_2745/ifx_xelse_ifx_xend_PhiReq/$entry
      -- CP-element group 66: 	 branch_block_stmt_2745/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3180/$entry
      -- CP-element group 66: 	 branch_block_stmt_2745/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3180/phi_stmt_3180_sources/$entry
      -- CP-element group 66: 	 branch_block_stmt_2745/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3180/phi_stmt_3180_sources/type_cast_3185/$entry
      -- CP-element group 66: 	 branch_block_stmt_2745/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3180/phi_stmt_3180_sources/type_cast_3185/SplitProtocol/$entry
      -- CP-element group 66: 	 branch_block_stmt_2745/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3180/phi_stmt_3180_sources/type_cast_3185/SplitProtocol/Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_2745/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3180/phi_stmt_3180_sources/type_cast_3185/SplitProtocol/Sample/rr
      -- CP-element group 66: 	 branch_block_stmt_2745/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3180/phi_stmt_3180_sources/type_cast_3185/SplitProtocol/Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_2745/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3180/phi_stmt_3180_sources/type_cast_3185/SplitProtocol/Update/cr
      -- CP-element group 66: 	 branch_block_stmt_2745/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3186/$entry
      -- CP-element group 66: 	 branch_block_stmt_2745/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3186/phi_stmt_3186_sources/$entry
      -- CP-element group 66: 	 branch_block_stmt_2745/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3186/phi_stmt_3186_sources/type_cast_3191/$entry
      -- CP-element group 66: 	 branch_block_stmt_2745/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3186/phi_stmt_3186_sources/type_cast_3191/SplitProtocol/$entry
      -- CP-element group 66: 	 branch_block_stmt_2745/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3186/phi_stmt_3186_sources/type_cast_3191/SplitProtocol/Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_2745/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3186/phi_stmt_3186_sources/type_cast_3191/SplitProtocol/Sample/rr
      -- CP-element group 66: 	 branch_block_stmt_2745/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3186/phi_stmt_3186_sources/type_cast_3191/SplitProtocol/Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_2745/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3186/phi_stmt_3186_sources/type_cast_3191/SplitProtocol/Update/cr
      -- 
    else_choice_transition_8534_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3155_branch_ack_0, ack => convTransposeD_CP_7576_elements(66)); -- 
    rr_8803_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8803_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(66), ack => type_cast_3185_inst_req_0); -- 
    cr_8808_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8808_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(66), ack => type_cast_3185_inst_req_1); -- 
    rr_8826_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8826_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(66), ack => type_cast_3191_inst_req_0); -- 
    cr_8831_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8831_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(66), ack => type_cast_3191_inst_req_1); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	65 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_2745/assign_stmt_3167_to_assign_stmt_3177/type_cast_3176_sample_completed_
      -- CP-element group 67: 	 branch_block_stmt_2745/assign_stmt_3167_to_assign_stmt_3177/type_cast_3176_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_2745/assign_stmt_3167_to_assign_stmt_3177/type_cast_3176_Sample/ra
      -- 
    ra_8548_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3176_inst_ack_0, ack => convTransposeD_CP_7576_elements(67)); -- 
    -- CP-element group 68:  fork  transition  place  input  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	65 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	109 
    -- CP-element group 68: 	110 
    -- CP-element group 68: 	106 
    -- CP-element group 68: 	107 
    -- CP-element group 68:  members (23) 
      -- CP-element group 68: 	 branch_block_stmt_2745/assign_stmt_3167_to_assign_stmt_3177__exit__
      -- CP-element group 68: 	 branch_block_stmt_2745/ifx_xthen83_ifx_xend
      -- CP-element group 68: 	 branch_block_stmt_2745/assign_stmt_3167_to_assign_stmt_3177/$exit
      -- CP-element group 68: 	 branch_block_stmt_2745/assign_stmt_3167_to_assign_stmt_3177/type_cast_3176_update_completed_
      -- CP-element group 68: 	 branch_block_stmt_2745/assign_stmt_3167_to_assign_stmt_3177/type_cast_3176_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_2745/assign_stmt_3167_to_assign_stmt_3177/type_cast_3176_Update/ca
      -- CP-element group 68: 	 branch_block_stmt_2745/ifx_xthen83_ifx_xend_PhiReq/$entry
      -- CP-element group 68: 	 branch_block_stmt_2745/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3180/$entry
      -- CP-element group 68: 	 branch_block_stmt_2745/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3180/phi_stmt_3180_sources/$entry
      -- CP-element group 68: 	 branch_block_stmt_2745/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3180/phi_stmt_3180_sources/type_cast_3183/$entry
      -- CP-element group 68: 	 branch_block_stmt_2745/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3180/phi_stmt_3180_sources/type_cast_3183/SplitProtocol/$entry
      -- CP-element group 68: 	 branch_block_stmt_2745/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3180/phi_stmt_3180_sources/type_cast_3183/SplitProtocol/Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_2745/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3180/phi_stmt_3180_sources/type_cast_3183/SplitProtocol/Sample/rr
      -- CP-element group 68: 	 branch_block_stmt_2745/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3180/phi_stmt_3180_sources/type_cast_3183/SplitProtocol/Update/$entry
      -- CP-element group 68: 	 branch_block_stmt_2745/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3180/phi_stmt_3180_sources/type_cast_3183/SplitProtocol/Update/cr
      -- CP-element group 68: 	 branch_block_stmt_2745/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3186/$entry
      -- CP-element group 68: 	 branch_block_stmt_2745/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3186/phi_stmt_3186_sources/$entry
      -- CP-element group 68: 	 branch_block_stmt_2745/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3186/phi_stmt_3186_sources/type_cast_3189/$entry
      -- CP-element group 68: 	 branch_block_stmt_2745/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3186/phi_stmt_3186_sources/type_cast_3189/SplitProtocol/$entry
      -- CP-element group 68: 	 branch_block_stmt_2745/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3186/phi_stmt_3186_sources/type_cast_3189/SplitProtocol/Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_2745/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3186/phi_stmt_3186_sources/type_cast_3189/SplitProtocol/Sample/rr
      -- CP-element group 68: 	 branch_block_stmt_2745/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3186/phi_stmt_3186_sources/type_cast_3189/SplitProtocol/Update/$entry
      -- CP-element group 68: 	 branch_block_stmt_2745/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3186/phi_stmt_3186_sources/type_cast_3189/SplitProtocol/Update/cr
      -- 
    ca_8553_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3176_inst_ack_1, ack => convTransposeD_CP_7576_elements(68)); -- 
    rr_8852_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8852_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(68), ack => type_cast_3183_inst_req_0); -- 
    cr_8857_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8857_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(68), ack => type_cast_3183_inst_req_1); -- 
    rr_8875_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8875_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(68), ack => type_cast_3189_inst_req_0); -- 
    cr_8880_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8880_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(68), ack => type_cast_3189_inst_req_1); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	116 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_2745/assign_stmt_3197_to_assign_stmt_3202/type_cast_3196_sample_completed_
      -- CP-element group 69: 	 branch_block_stmt_2745/assign_stmt_3197_to_assign_stmt_3202/type_cast_3196_Sample/$exit
      -- CP-element group 69: 	 branch_block_stmt_2745/assign_stmt_3197_to_assign_stmt_3202/type_cast_3196_Sample/ra
      -- 
    ra_8565_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3196_inst_ack_0, ack => convTransposeD_CP_7576_elements(69)); -- 
    -- CP-element group 70:  branch  transition  place  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	116 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (13) 
      -- CP-element group 70: 	 branch_block_stmt_2745/R_cmp92_3204_place
      -- CP-element group 70: 	 branch_block_stmt_2745/if_stmt_3203_eval_test/$entry
      -- CP-element group 70: 	 branch_block_stmt_2745/assign_stmt_3197_to_assign_stmt_3202__exit__
      -- CP-element group 70: 	 branch_block_stmt_2745/if_stmt_3203__entry__
      -- CP-element group 70: 	 branch_block_stmt_2745/assign_stmt_3197_to_assign_stmt_3202/$exit
      -- CP-element group 70: 	 branch_block_stmt_2745/assign_stmt_3197_to_assign_stmt_3202/type_cast_3196_update_completed_
      -- CP-element group 70: 	 branch_block_stmt_2745/assign_stmt_3197_to_assign_stmt_3202/type_cast_3196_Update/$exit
      -- CP-element group 70: 	 branch_block_stmt_2745/assign_stmt_3197_to_assign_stmt_3202/type_cast_3196_Update/ca
      -- CP-element group 70: 	 branch_block_stmt_2745/if_stmt_3203_dead_link/$entry
      -- CP-element group 70: 	 branch_block_stmt_2745/if_stmt_3203_eval_test/$exit
      -- CP-element group 70: 	 branch_block_stmt_2745/if_stmt_3203_eval_test/branch_req
      -- CP-element group 70: 	 branch_block_stmt_2745/if_stmt_3203_if_link/$entry
      -- CP-element group 70: 	 branch_block_stmt_2745/if_stmt_3203_else_link/$entry
      -- 
    ca_8570_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3196_inst_ack_1, ack => convTransposeD_CP_7576_elements(70)); -- 
    branch_req_8578_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_8578_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(70), ack => if_stmt_3203_branch_req_0); -- 
    -- CP-element group 71:  merge  transition  place  input  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (15) 
      -- CP-element group 71: 	 branch_block_stmt_2745/ifx_xend_whilex_xend
      -- CP-element group 71: 	 branch_block_stmt_2745/merge_stmt_3209__exit__
      -- CP-element group 71: 	 branch_block_stmt_2745/assign_stmt_3213__entry__
      -- CP-element group 71: 	 branch_block_stmt_2745/if_stmt_3203_if_link/$exit
      -- CP-element group 71: 	 branch_block_stmt_2745/if_stmt_3203_if_link/if_choice_transition
      -- CP-element group 71: 	 branch_block_stmt_2745/assign_stmt_3213/$entry
      -- CP-element group 71: 	 branch_block_stmt_2745/assign_stmt_3213/WPIPE_Block3_done_3211_sample_start_
      -- CP-element group 71: 	 branch_block_stmt_2745/assign_stmt_3213/WPIPE_Block3_done_3211_Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_2745/assign_stmt_3213/WPIPE_Block3_done_3211_Sample/req
      -- CP-element group 71: 	 branch_block_stmt_2745/ifx_xend_whilex_xend_PhiReq/$entry
      -- CP-element group 71: 	 branch_block_stmt_2745/ifx_xend_whilex_xend_PhiReq/$exit
      -- CP-element group 71: 	 branch_block_stmt_2745/merge_stmt_3209_PhiReqMerge
      -- CP-element group 71: 	 branch_block_stmt_2745/merge_stmt_3209_PhiAck/$entry
      -- CP-element group 71: 	 branch_block_stmt_2745/merge_stmt_3209_PhiAck/$exit
      -- CP-element group 71: 	 branch_block_stmt_2745/merge_stmt_3209_PhiAck/dummy
      -- 
    if_choice_transition_8583_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3203_branch_ack_1, ack => convTransposeD_CP_7576_elements(71)); -- 
    req_8600_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8600_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(71), ack => WPIPE_Block3_done_3211_inst_req_0); -- 
    -- CP-element group 72:  fork  transition  place  input  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	82 
    -- CP-element group 72: 	83 
    -- CP-element group 72: 	85 
    -- CP-element group 72: 	86 
    -- CP-element group 72:  members (20) 
      -- CP-element group 72: 	 branch_block_stmt_2745/ifx_xend_whilex_xbodyx_xouter
      -- CP-element group 72: 	 branch_block_stmt_2745/if_stmt_3203_else_link/$exit
      -- CP-element group 72: 	 branch_block_stmt_2745/if_stmt_3203_else_link/else_choice_transition
      -- CP-element group 72: 	 branch_block_stmt_2745/ifx_xend_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 72: 	 branch_block_stmt_2745/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2891/$entry
      -- CP-element group 72: 	 branch_block_stmt_2745/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2891/phi_stmt_2891_sources/$entry
      -- CP-element group 72: 	 branch_block_stmt_2745/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2891/phi_stmt_2891_sources/type_cast_2896/$entry
      -- CP-element group 72: 	 branch_block_stmt_2745/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2891/phi_stmt_2891_sources/type_cast_2896/SplitProtocol/$entry
      -- CP-element group 72: 	 branch_block_stmt_2745/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2891/phi_stmt_2891_sources/type_cast_2896/SplitProtocol/Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_2745/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2891/phi_stmt_2891_sources/type_cast_2896/SplitProtocol/Sample/rr
      -- CP-element group 72: 	 branch_block_stmt_2745/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2891/phi_stmt_2891_sources/type_cast_2896/SplitProtocol/Update/$entry
      -- CP-element group 72: 	 branch_block_stmt_2745/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2891/phi_stmt_2891_sources/type_cast_2896/SplitProtocol/Update/cr
      -- CP-element group 72: 	 branch_block_stmt_2745/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2897/$entry
      -- CP-element group 72: 	 branch_block_stmt_2745/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2897/phi_stmt_2897_sources/$entry
      -- CP-element group 72: 	 branch_block_stmt_2745/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2897/phi_stmt_2897_sources/type_cast_2902/$entry
      -- CP-element group 72: 	 branch_block_stmt_2745/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2897/phi_stmt_2897_sources/type_cast_2902/SplitProtocol/$entry
      -- CP-element group 72: 	 branch_block_stmt_2745/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2897/phi_stmt_2897_sources/type_cast_2902/SplitProtocol/Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_2745/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2897/phi_stmt_2897_sources/type_cast_2902/SplitProtocol/Sample/rr
      -- CP-element group 72: 	 branch_block_stmt_2745/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2897/phi_stmt_2897_sources/type_cast_2902/SplitProtocol/Update/$entry
      -- CP-element group 72: 	 branch_block_stmt_2745/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2897/phi_stmt_2897_sources/type_cast_2902/SplitProtocol/Update/cr
      -- 
    else_choice_transition_8587_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3203_branch_ack_0, ack => convTransposeD_CP_7576_elements(72)); -- 
    rr_8674_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8674_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(72), ack => type_cast_2896_inst_req_0); -- 
    cr_8679_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8679_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(72), ack => type_cast_2896_inst_req_1); -- 
    rr_8697_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8697_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(72), ack => type_cast_2902_inst_req_0); -- 
    cr_8702_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8702_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(72), ack => type_cast_2902_inst_req_1); -- 
    -- CP-element group 73:  transition  input  output  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (6) 
      -- CP-element group 73: 	 branch_block_stmt_2745/assign_stmt_3213/WPIPE_Block3_done_3211_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_2745/assign_stmt_3213/WPIPE_Block3_done_3211_update_start_
      -- CP-element group 73: 	 branch_block_stmt_2745/assign_stmt_3213/WPIPE_Block3_done_3211_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_2745/assign_stmt_3213/WPIPE_Block3_done_3211_Sample/ack
      -- CP-element group 73: 	 branch_block_stmt_2745/assign_stmt_3213/WPIPE_Block3_done_3211_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_2745/assign_stmt_3213/WPIPE_Block3_done_3211_Update/req
      -- 
    ack_8601_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_done_3211_inst_ack_0, ack => convTransposeD_CP_7576_elements(73)); -- 
    req_8605_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8605_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(73), ack => WPIPE_Block3_done_3211_inst_req_1); -- 
    -- CP-element group 74:  transition  place  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (16) 
      -- CP-element group 74: 	 branch_block_stmt_2745/branch_block_stmt_2745__exit__
      -- CP-element group 74: 	 branch_block_stmt_2745/$exit
      -- CP-element group 74: 	 $exit
      -- CP-element group 74: 	 branch_block_stmt_2745/assign_stmt_3213__exit__
      -- CP-element group 74: 	 branch_block_stmt_2745/return__
      -- CP-element group 74: 	 branch_block_stmt_2745/merge_stmt_3215__exit__
      -- CP-element group 74: 	 branch_block_stmt_2745/assign_stmt_3213/$exit
      -- CP-element group 74: 	 branch_block_stmt_2745/assign_stmt_3213/WPIPE_Block3_done_3211_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_2745/assign_stmt_3213/WPIPE_Block3_done_3211_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_2745/assign_stmt_3213/WPIPE_Block3_done_3211_Update/ack
      -- CP-element group 74: 	 branch_block_stmt_2745/return___PhiReq/$entry
      -- CP-element group 74: 	 branch_block_stmt_2745/return___PhiReq/$exit
      -- CP-element group 74: 	 branch_block_stmt_2745/merge_stmt_3215_PhiReqMerge
      -- CP-element group 74: 	 branch_block_stmt_2745/merge_stmt_3215_PhiAck/$entry
      -- CP-element group 74: 	 branch_block_stmt_2745/merge_stmt_3215_PhiAck/$exit
      -- CP-element group 74: 	 branch_block_stmt_2745/merge_stmt_3215_PhiAck/dummy
      -- 
    ack_8606_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_done_3211_inst_ack_1, ack => convTransposeD_CP_7576_elements(74)); -- 
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	33 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (2) 
      -- CP-element group 75: 	 branch_block_stmt_2745/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2891/phi_stmt_2891_sources/type_cast_2894/SplitProtocol/Sample/$exit
      -- CP-element group 75: 	 branch_block_stmt_2745/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2891/phi_stmt_2891_sources/type_cast_2894/SplitProtocol/Sample/ra
      -- 
    ra_8626_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2894_inst_ack_0, ack => convTransposeD_CP_7576_elements(75)); -- 
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	33 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76:  members (2) 
      -- CP-element group 76: 	 branch_block_stmt_2745/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2891/phi_stmt_2891_sources/type_cast_2894/SplitProtocol/Update/$exit
      -- CP-element group 76: 	 branch_block_stmt_2745/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2891/phi_stmt_2891_sources/type_cast_2894/SplitProtocol/Update/ca
      -- 
    ca_8631_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2894_inst_ack_1, ack => convTransposeD_CP_7576_elements(76)); -- 
    -- CP-element group 77:  join  transition  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: 	76 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	81 
    -- CP-element group 77:  members (5) 
      -- CP-element group 77: 	 branch_block_stmt_2745/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2891/$exit
      -- CP-element group 77: 	 branch_block_stmt_2745/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2891/phi_stmt_2891_sources/$exit
      -- CP-element group 77: 	 branch_block_stmt_2745/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2891/phi_stmt_2891_sources/type_cast_2894/$exit
      -- CP-element group 77: 	 branch_block_stmt_2745/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2891/phi_stmt_2891_sources/type_cast_2894/SplitProtocol/$exit
      -- CP-element group 77: 	 branch_block_stmt_2745/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2891/phi_stmt_2891_req
      -- 
    phi_stmt_2891_req_8632_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2891_req_8632_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(77), ack => phi_stmt_2891_req_0); -- 
    convTransposeD_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7576_elements(75) & convTransposeD_CP_7576_elements(76);
      gj_convTransposeD_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7576_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	33 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	80 
    -- CP-element group 78:  members (2) 
      -- CP-element group 78: 	 branch_block_stmt_2745/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2897/phi_stmt_2897_sources/type_cast_2900/SplitProtocol/Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_2745/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2897/phi_stmt_2897_sources/type_cast_2900/SplitProtocol/Sample/ra
      -- 
    ra_8649_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2900_inst_ack_0, ack => convTransposeD_CP_7576_elements(78)); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	33 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_2745/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2897/phi_stmt_2897_sources/type_cast_2900/SplitProtocol/Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_2745/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2897/phi_stmt_2897_sources/type_cast_2900/SplitProtocol/Update/ca
      -- 
    ca_8654_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2900_inst_ack_1, ack => convTransposeD_CP_7576_elements(79)); -- 
    -- CP-element group 80:  join  transition  output  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (5) 
      -- CP-element group 80: 	 branch_block_stmt_2745/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2897/$exit
      -- CP-element group 80: 	 branch_block_stmt_2745/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2897/phi_stmt_2897_sources/$exit
      -- CP-element group 80: 	 branch_block_stmt_2745/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2897/phi_stmt_2897_sources/type_cast_2900/$exit
      -- CP-element group 80: 	 branch_block_stmt_2745/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2897/phi_stmt_2897_sources/type_cast_2900/SplitProtocol/$exit
      -- CP-element group 80: 	 branch_block_stmt_2745/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2897/phi_stmt_2897_req
      -- 
    phi_stmt_2897_req_8655_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2897_req_8655_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(80), ack => phi_stmt_2897_req_0); -- 
    convTransposeD_cp_element_group_80: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_80"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7576_elements(78) & convTransposeD_CP_7576_elements(79);
      gj_convTransposeD_cp_element_group_80 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7576_elements(80), clk => clk, reset => reset); --
    end block;
    -- CP-element group 81:  join  transition  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	77 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	89 
    -- CP-element group 81:  members (1) 
      -- CP-element group 81: 	 branch_block_stmt_2745/entry_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7576_elements(77) & convTransposeD_CP_7576_elements(80);
      gj_convTransposeD_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7576_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	72 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	84 
    -- CP-element group 82:  members (2) 
      -- CP-element group 82: 	 branch_block_stmt_2745/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2891/phi_stmt_2891_sources/type_cast_2896/SplitProtocol/Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_2745/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2891/phi_stmt_2891_sources/type_cast_2896/SplitProtocol/Sample/ra
      -- 
    ra_8675_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2896_inst_ack_0, ack => convTransposeD_CP_7576_elements(82)); -- 
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	72 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_2745/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2891/phi_stmt_2891_sources/type_cast_2896/SplitProtocol/Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_2745/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2891/phi_stmt_2891_sources/type_cast_2896/SplitProtocol/Update/ca
      -- 
    ca_8680_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2896_inst_ack_1, ack => convTransposeD_CP_7576_elements(83)); -- 
    -- CP-element group 84:  join  transition  output  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	88 
    -- CP-element group 84:  members (5) 
      -- CP-element group 84: 	 branch_block_stmt_2745/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2891/$exit
      -- CP-element group 84: 	 branch_block_stmt_2745/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2891/phi_stmt_2891_sources/$exit
      -- CP-element group 84: 	 branch_block_stmt_2745/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2891/phi_stmt_2891_sources/type_cast_2896/$exit
      -- CP-element group 84: 	 branch_block_stmt_2745/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2891/phi_stmt_2891_sources/type_cast_2896/SplitProtocol/$exit
      -- CP-element group 84: 	 branch_block_stmt_2745/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2891/phi_stmt_2891_req
      -- 
    phi_stmt_2891_req_8681_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2891_req_8681_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(84), ack => phi_stmt_2891_req_1); -- 
    convTransposeD_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7576_elements(82) & convTransposeD_CP_7576_elements(83);
      gj_convTransposeD_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7576_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	72 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (2) 
      -- CP-element group 85: 	 branch_block_stmt_2745/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2897/phi_stmt_2897_sources/type_cast_2902/SplitProtocol/Sample/$exit
      -- CP-element group 85: 	 branch_block_stmt_2745/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2897/phi_stmt_2897_sources/type_cast_2902/SplitProtocol/Sample/ra
      -- 
    ra_8698_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2902_inst_ack_0, ack => convTransposeD_CP_7576_elements(85)); -- 
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	72 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_2745/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2897/phi_stmt_2897_sources/type_cast_2902/SplitProtocol/Update/$exit
      -- CP-element group 86: 	 branch_block_stmt_2745/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2897/phi_stmt_2897_sources/type_cast_2902/SplitProtocol/Update/ca
      -- 
    ca_8703_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2902_inst_ack_1, ack => convTransposeD_CP_7576_elements(86)); -- 
    -- CP-element group 87:  join  transition  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (5) 
      -- CP-element group 87: 	 branch_block_stmt_2745/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2897/$exit
      -- CP-element group 87: 	 branch_block_stmt_2745/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2897/phi_stmt_2897_sources/$exit
      -- CP-element group 87: 	 branch_block_stmt_2745/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2897/phi_stmt_2897_sources/type_cast_2902/$exit
      -- CP-element group 87: 	 branch_block_stmt_2745/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2897/phi_stmt_2897_sources/type_cast_2902/SplitProtocol/$exit
      -- CP-element group 87: 	 branch_block_stmt_2745/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2897/phi_stmt_2897_req
      -- 
    phi_stmt_2897_req_8704_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2897_req_8704_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(87), ack => phi_stmt_2897_req_1); -- 
    convTransposeD_cp_element_group_87: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_87"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7576_elements(85) & convTransposeD_CP_7576_elements(86);
      gj_convTransposeD_cp_element_group_87 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7576_elements(87), clk => clk, reset => reset); --
    end block;
    -- CP-element group 88:  join  transition  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	84 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	89 
    -- CP-element group 88:  members (1) 
      -- CP-element group 88: 	 branch_block_stmt_2745/ifx_xend_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_88: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_88"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7576_elements(84) & convTransposeD_CP_7576_elements(87);
      gj_convTransposeD_cp_element_group_88 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7576_elements(88), clk => clk, reset => reset); --
    end block;
    -- CP-element group 89:  merge  fork  transition  place  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	81 
    -- CP-element group 89: 	88 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	90 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (2) 
      -- CP-element group 89: 	 branch_block_stmt_2745/merge_stmt_2890_PhiReqMerge
      -- CP-element group 89: 	 branch_block_stmt_2745/merge_stmt_2890_PhiAck/$entry
      -- 
    convTransposeD_CP_7576_elements(89) <= OrReduce(convTransposeD_CP_7576_elements(81) & convTransposeD_CP_7576_elements(88));
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	89 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	92 
    -- CP-element group 90:  members (1) 
      -- CP-element group 90: 	 branch_block_stmt_2745/merge_stmt_2890_PhiAck/phi_stmt_2891_ack
      -- 
    phi_stmt_2891_ack_8709_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2891_ack_0, ack => convTransposeD_CP_7576_elements(90)); -- 
    -- CP-element group 91:  transition  input  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (1) 
      -- CP-element group 91: 	 branch_block_stmt_2745/merge_stmt_2890_PhiAck/phi_stmt_2897_ack
      -- 
    phi_stmt_2897_ack_8710_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2897_ack_0, ack => convTransposeD_CP_7576_elements(91)); -- 
    -- CP-element group 92:  join  fork  transition  place  output  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	90 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	36 
    -- CP-element group 92: 	37 
    -- CP-element group 92: 	34 
    -- CP-element group 92: 	35 
    -- CP-element group 92:  members (16) 
      -- CP-element group 92: 	 branch_block_stmt_2745/assign_stmt_2908_to_assign_stmt_3015/type_cast_2912_Sample/rr
      -- CP-element group 92: 	 branch_block_stmt_2745/assign_stmt_2908_to_assign_stmt_3015/type_cast_2907_Update/cr
      -- CP-element group 92: 	 branch_block_stmt_2745/assign_stmt_2908_to_assign_stmt_3015/$entry
      -- CP-element group 92: 	 branch_block_stmt_2745/assign_stmt_2908_to_assign_stmt_3015/type_cast_2912_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2745/assign_stmt_2908_to_assign_stmt_3015/type_cast_2907_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2745/assign_stmt_2908_to_assign_stmt_3015/type_cast_2912_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_2745/assign_stmt_2908_to_assign_stmt_3015/type_cast_2907_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_2745/assign_stmt_2908_to_assign_stmt_3015/type_cast_2912_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2745/assign_stmt_2908_to_assign_stmt_3015/type_cast_2907_Sample/rr
      -- CP-element group 92: 	 branch_block_stmt_2745/assign_stmt_2908_to_assign_stmt_3015/type_cast_2907_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2745/assign_stmt_2908_to_assign_stmt_3015/type_cast_2912_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_2745/assign_stmt_2908_to_assign_stmt_3015/type_cast_2907_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_2745/assign_stmt_2908_to_assign_stmt_3015/type_cast_2912_Update/cr
      -- CP-element group 92: 	 branch_block_stmt_2745/merge_stmt_2890__exit__
      -- CP-element group 92: 	 branch_block_stmt_2745/assign_stmt_2908_to_assign_stmt_3015__entry__
      -- CP-element group 92: 	 branch_block_stmt_2745/merge_stmt_2890_PhiAck/$exit
      -- 
    rr_8221_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8221_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(92), ack => type_cast_2912_inst_req_0); -- 
    cr_8212_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8212_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(92), ack => type_cast_2907_inst_req_1); -- 
    rr_8207_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8207_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(92), ack => type_cast_2907_inst_req_0); -- 
    cr_8226_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8226_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(92), ack => type_cast_2912_inst_req_1); -- 
    convTransposeD_cp_element_group_92: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_92"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7576_elements(90) & convTransposeD_CP_7576_elements(91);
      gj_convTransposeD_cp_element_group_92 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7576_elements(92), clk => clk, reset => reset); --
    end block;
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	61 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (2) 
      -- CP-element group 93: 	 branch_block_stmt_2745/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3018/phi_stmt_3018_sources/type_cast_3024/SplitProtocol/Sample/$exit
      -- CP-element group 93: 	 branch_block_stmt_2745/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3018/phi_stmt_3018_sources/type_cast_3024/SplitProtocol/Sample/ra
      -- 
    ra_8730_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3024_inst_ack_0, ack => convTransposeD_CP_7576_elements(93)); -- 
    -- CP-element group 94:  transition  input  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	61 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94:  members (2) 
      -- CP-element group 94: 	 branch_block_stmt_2745/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3018/phi_stmt_3018_sources/type_cast_3024/SplitProtocol/Update/$exit
      -- CP-element group 94: 	 branch_block_stmt_2745/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3018/phi_stmt_3018_sources/type_cast_3024/SplitProtocol/Update/ca
      -- 
    ca_8735_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3024_inst_ack_1, ack => convTransposeD_CP_7576_elements(94)); -- 
    -- CP-element group 95:  join  transition  output  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	97 
    -- CP-element group 95:  members (6) 
      -- CP-element group 95: 	 branch_block_stmt_2745/ifx_xthen_whilex_xbody_PhiReq/$exit
      -- CP-element group 95: 	 branch_block_stmt_2745/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3018/$exit
      -- CP-element group 95: 	 branch_block_stmt_2745/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3018/phi_stmt_3018_sources/$exit
      -- CP-element group 95: 	 branch_block_stmt_2745/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3018/phi_stmt_3018_sources/type_cast_3024/$exit
      -- CP-element group 95: 	 branch_block_stmt_2745/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3018/phi_stmt_3018_sources/type_cast_3024/SplitProtocol/$exit
      -- CP-element group 95: 	 branch_block_stmt_2745/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3018/phi_stmt_3018_req
      -- 
    phi_stmt_3018_req_8736_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3018_req_8736_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(95), ack => phi_stmt_3018_req_1); -- 
    convTransposeD_cp_element_group_95: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_95"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7576_elements(93) & convTransposeD_CP_7576_elements(94);
      gj_convTransposeD_cp_element_group_95 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7576_elements(95), clk => clk, reset => reset); --
    end block;
    -- CP-element group 96:  transition  output  delay-element  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	38 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (5) 
      -- CP-element group 96: 	 branch_block_stmt_2745/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$exit
      -- CP-element group 96: 	 branch_block_stmt_2745/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_3018/$exit
      -- CP-element group 96: 	 branch_block_stmt_2745/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_3018/phi_stmt_3018_sources/$exit
      -- CP-element group 96: 	 branch_block_stmt_2745/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_3018/phi_stmt_3018_sources/type_cast_3022_konst_delay_trans
      -- CP-element group 96: 	 branch_block_stmt_2745/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_3018/phi_stmt_3018_req
      -- 
    phi_stmt_3018_req_8747_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3018_req_8747_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(96), ack => phi_stmt_3018_req_0); -- 
    -- Element group convTransposeD_CP_7576_elements(96) is a control-delay.
    cp_element_96_delay: control_delay_element  generic map(name => " 96_delay", delay_value => 1)  port map(req => convTransposeD_CP_7576_elements(38), ack => convTransposeD_CP_7576_elements(96), clk => clk, reset =>reset);
    -- CP-element group 97:  merge  transition  place  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97:  members (2) 
      -- CP-element group 97: 	 branch_block_stmt_2745/merge_stmt_3017_PhiReqMerge
      -- CP-element group 97: 	 branch_block_stmt_2745/merge_stmt_3017_PhiAck/$entry
      -- 
    convTransposeD_CP_7576_elements(97) <= OrReduce(convTransposeD_CP_7576_elements(95) & convTransposeD_CP_7576_elements(96));
    -- CP-element group 98:  fork  transition  place  input  output  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	46 
    -- CP-element group 98: 	52 
    -- CP-element group 98: 	57 
    -- CP-element group 98: 	48 
    -- CP-element group 98: 	42 
    -- CP-element group 98: 	44 
    -- CP-element group 98: 	39 
    -- CP-element group 98: 	40 
    -- CP-element group 98: 	58 
    -- CP-element group 98: 	59 
    -- CP-element group 98: 	54 
    -- CP-element group 98: 	50 
    -- CP-element group 98:  members (45) 
      -- CP-element group 98: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/type_cast_3034_Sample/rr
      -- CP-element group 98: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/type_cast_3064_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3075_update_start_
      -- CP-element group 98: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/array_obj_ref_3070_final_index_sum_regn_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/array_obj_ref_3070_final_index_sum_regn_Update/req
      -- CP-element group 98: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/addr_of_3071_update_start_
      -- CP-element group 98: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/array_obj_ref_3070_final_index_sum_regn_update_start
      -- CP-element group 98: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/type_cast_3034_Sample/$entry
      -- CP-element group 98: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/type_cast_3034_update_start_
      -- CP-element group 98: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/addr_of_3071_complete/req
      -- CP-element group 98: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/type_cast_3034_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/type_cast_3064_update_start_
      -- CP-element group 98: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/type_cast_3034_Update/cr
      -- CP-element group 98: 	 branch_block_stmt_2745/merge_stmt_3017__exit__
      -- CP-element group 98: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123__entry__
      -- CP-element group 98: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/type_cast_3034_sample_start_
      -- CP-element group 98: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/addr_of_3071_complete/$entry
      -- CP-element group 98: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/type_cast_3064_Update/cr
      -- CP-element group 98: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/$entry
      -- CP-element group 98: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3075_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3075_Update/word_access_complete/$entry
      -- CP-element group 98: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3075_Update/word_access_complete/word_0/$entry
      -- CP-element group 98: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3075_Update/word_access_complete/word_0/cr
      -- CP-element group 98: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/type_cast_3095_update_start_
      -- CP-element group 98: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/type_cast_3095_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/type_cast_3095_Update/cr
      -- CP-element group 98: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/addr_of_3102_update_start_
      -- CP-element group 98: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/array_obj_ref_3101_final_index_sum_regn_update_start
      -- CP-element group 98: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/array_obj_ref_3101_final_index_sum_regn_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/array_obj_ref_3101_final_index_sum_regn_Update/req
      -- CP-element group 98: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/addr_of_3102_complete/$entry
      -- CP-element group 98: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/addr_of_3102_complete/req
      -- CP-element group 98: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3105_update_start_
      -- CP-element group 98: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3105_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3105_Update/word_access_complete/$entry
      -- CP-element group 98: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3105_Update/word_access_complete/word_0/$entry
      -- CP-element group 98: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/ptr_deref_3105_Update/word_access_complete/word_0/cr
      -- CP-element group 98: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/type_cast_3111_sample_start_
      -- CP-element group 98: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/type_cast_3111_update_start_
      -- CP-element group 98: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/type_cast_3111_Sample/$entry
      -- CP-element group 98: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/type_cast_3111_Sample/rr
      -- CP-element group 98: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/type_cast_3111_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_2745/assign_stmt_3031_to_assign_stmt_3123/type_cast_3111_Update/cr
      -- CP-element group 98: 	 branch_block_stmt_2745/merge_stmt_3017_PhiAck/$exit
      -- CP-element group 98: 	 branch_block_stmt_2745/merge_stmt_3017_PhiAck/phi_stmt_3018_ack
      -- 
    phi_stmt_3018_ack_8752_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3018_ack_0, ack => convTransposeD_CP_7576_elements(98)); -- 
    rr_8238_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8238_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(98), ack => type_cast_3034_inst_req_0); -- 
    req_8288_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8288_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(98), ack => array_obj_ref_3070_index_offset_req_1); -- 
    req_8303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(98), ack => addr_of_3071_final_reg_req_1); -- 
    cr_8243_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8243_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(98), ack => type_cast_3034_inst_req_1); -- 
    cr_8257_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8257_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(98), ack => type_cast_3064_inst_req_1); -- 
    cr_8348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(98), ack => ptr_deref_3075_load_0_req_1); -- 
    cr_8367_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8367_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(98), ack => type_cast_3095_inst_req_1); -- 
    req_8398_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8398_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(98), ack => array_obj_ref_3101_index_offset_req_1); -- 
    req_8413_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8413_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(98), ack => addr_of_3102_final_reg_req_1); -- 
    cr_8463_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8463_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(98), ack => ptr_deref_3105_store_0_req_1); -- 
    rr_8472_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8472_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(98), ack => type_cast_3111_inst_req_0); -- 
    cr_8477_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8477_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(98), ack => type_cast_3111_inst_req_1); -- 
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	66 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	101 
    -- CP-element group 99:  members (2) 
      -- CP-element group 99: 	 branch_block_stmt_2745/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3180/phi_stmt_3180_sources/type_cast_3185/SplitProtocol/Sample/$exit
      -- CP-element group 99: 	 branch_block_stmt_2745/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3180/phi_stmt_3180_sources/type_cast_3185/SplitProtocol/Sample/ra
      -- 
    ra_8804_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3185_inst_ack_0, ack => convTransposeD_CP_7576_elements(99)); -- 
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	66 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	101 
    -- CP-element group 100:  members (2) 
      -- CP-element group 100: 	 branch_block_stmt_2745/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3180/phi_stmt_3180_sources/type_cast_3185/SplitProtocol/Update/$exit
      -- CP-element group 100: 	 branch_block_stmt_2745/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3180/phi_stmt_3180_sources/type_cast_3185/SplitProtocol/Update/ca
      -- 
    ca_8809_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3185_inst_ack_1, ack => convTransposeD_CP_7576_elements(100)); -- 
    -- CP-element group 101:  join  transition  output  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	99 
    -- CP-element group 101: 	100 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	105 
    -- CP-element group 101:  members (5) 
      -- CP-element group 101: 	 branch_block_stmt_2745/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3180/$exit
      -- CP-element group 101: 	 branch_block_stmt_2745/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3180/phi_stmt_3180_sources/$exit
      -- CP-element group 101: 	 branch_block_stmt_2745/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3180/phi_stmt_3180_sources/type_cast_3185/$exit
      -- CP-element group 101: 	 branch_block_stmt_2745/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3180/phi_stmt_3180_sources/type_cast_3185/SplitProtocol/$exit
      -- CP-element group 101: 	 branch_block_stmt_2745/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3180/phi_stmt_3180_req
      -- 
    phi_stmt_3180_req_8810_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3180_req_8810_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(101), ack => phi_stmt_3180_req_1); -- 
    convTransposeD_cp_element_group_101: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_101"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7576_elements(99) & convTransposeD_CP_7576_elements(100);
      gj_convTransposeD_cp_element_group_101 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7576_elements(101), clk => clk, reset => reset); --
    end block;
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	66 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	104 
    -- CP-element group 102:  members (2) 
      -- CP-element group 102: 	 branch_block_stmt_2745/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3186/phi_stmt_3186_sources/type_cast_3191/SplitProtocol/Sample/$exit
      -- CP-element group 102: 	 branch_block_stmt_2745/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3186/phi_stmt_3186_sources/type_cast_3191/SplitProtocol/Sample/ra
      -- 
    ra_8827_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3191_inst_ack_0, ack => convTransposeD_CP_7576_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	66 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (2) 
      -- CP-element group 103: 	 branch_block_stmt_2745/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3186/phi_stmt_3186_sources/type_cast_3191/SplitProtocol/Update/$exit
      -- CP-element group 103: 	 branch_block_stmt_2745/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3186/phi_stmt_3186_sources/type_cast_3191/SplitProtocol/Update/ca
      -- 
    ca_8832_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3191_inst_ack_1, ack => convTransposeD_CP_7576_elements(103)); -- 
    -- CP-element group 104:  join  transition  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	103 
    -- CP-element group 104: 	102 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	105 
    -- CP-element group 104:  members (5) 
      -- CP-element group 104: 	 branch_block_stmt_2745/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3186/$exit
      -- CP-element group 104: 	 branch_block_stmt_2745/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3186/phi_stmt_3186_sources/$exit
      -- CP-element group 104: 	 branch_block_stmt_2745/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3186/phi_stmt_3186_sources/type_cast_3191/$exit
      -- CP-element group 104: 	 branch_block_stmt_2745/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3186/phi_stmt_3186_sources/type_cast_3191/SplitProtocol/$exit
      -- CP-element group 104: 	 branch_block_stmt_2745/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3186/phi_stmt_3186_req
      -- 
    phi_stmt_3186_req_8833_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3186_req_8833_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(104), ack => phi_stmt_3186_req_1); -- 
    convTransposeD_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7576_elements(103) & convTransposeD_CP_7576_elements(102);
      gj_convTransposeD_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7576_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  join  transition  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	104 
    -- CP-element group 105: 	101 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	113 
    -- CP-element group 105:  members (1) 
      -- CP-element group 105: 	 branch_block_stmt_2745/ifx_xelse_ifx_xend_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_105: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_105"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7576_elements(104) & convTransposeD_CP_7576_elements(101);
      gj_convTransposeD_cp_element_group_105 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7576_elements(105), clk => clk, reset => reset); --
    end block;
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	68 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	108 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_2745/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3180/phi_stmt_3180_sources/type_cast_3183/SplitProtocol/Sample/$exit
      -- CP-element group 106: 	 branch_block_stmt_2745/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3180/phi_stmt_3180_sources/type_cast_3183/SplitProtocol/Sample/ra
      -- 
    ra_8853_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3183_inst_ack_0, ack => convTransposeD_CP_7576_elements(106)); -- 
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	68 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107:  members (2) 
      -- CP-element group 107: 	 branch_block_stmt_2745/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3180/phi_stmt_3180_sources/type_cast_3183/SplitProtocol/Update/$exit
      -- CP-element group 107: 	 branch_block_stmt_2745/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3180/phi_stmt_3180_sources/type_cast_3183/SplitProtocol/Update/ca
      -- 
    ca_8858_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3183_inst_ack_1, ack => convTransposeD_CP_7576_elements(107)); -- 
    -- CP-element group 108:  join  transition  output  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	106 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	112 
    -- CP-element group 108:  members (5) 
      -- CP-element group 108: 	 branch_block_stmt_2745/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3180/$exit
      -- CP-element group 108: 	 branch_block_stmt_2745/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3180/phi_stmt_3180_sources/$exit
      -- CP-element group 108: 	 branch_block_stmt_2745/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3180/phi_stmt_3180_sources/type_cast_3183/$exit
      -- CP-element group 108: 	 branch_block_stmt_2745/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3180/phi_stmt_3180_sources/type_cast_3183/SplitProtocol/$exit
      -- CP-element group 108: 	 branch_block_stmt_2745/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3180/phi_stmt_3180_req
      -- 
    phi_stmt_3180_req_8859_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3180_req_8859_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(108), ack => phi_stmt_3180_req_0); -- 
    convTransposeD_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7576_elements(106) & convTransposeD_CP_7576_elements(107);
      gj_convTransposeD_cp_element_group_108 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7576_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	68 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (2) 
      -- CP-element group 109: 	 branch_block_stmt_2745/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3186/phi_stmt_3186_sources/type_cast_3189/SplitProtocol/Sample/$exit
      -- CP-element group 109: 	 branch_block_stmt_2745/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3186/phi_stmt_3186_sources/type_cast_3189/SplitProtocol/Sample/ra
      -- 
    ra_8876_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3189_inst_ack_0, ack => convTransposeD_CP_7576_elements(109)); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	68 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (2) 
      -- CP-element group 110: 	 branch_block_stmt_2745/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3186/phi_stmt_3186_sources/type_cast_3189/SplitProtocol/Update/$exit
      -- CP-element group 110: 	 branch_block_stmt_2745/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3186/phi_stmt_3186_sources/type_cast_3189/SplitProtocol/Update/ca
      -- 
    ca_8881_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3189_inst_ack_1, ack => convTransposeD_CP_7576_elements(110)); -- 
    -- CP-element group 111:  join  transition  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111:  members (5) 
      -- CP-element group 111: 	 branch_block_stmt_2745/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3186/$exit
      -- CP-element group 111: 	 branch_block_stmt_2745/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3186/phi_stmt_3186_sources/$exit
      -- CP-element group 111: 	 branch_block_stmt_2745/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3186/phi_stmt_3186_sources/type_cast_3189/$exit
      -- CP-element group 111: 	 branch_block_stmt_2745/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3186/phi_stmt_3186_sources/type_cast_3189/SplitProtocol/$exit
      -- CP-element group 111: 	 branch_block_stmt_2745/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3186/phi_stmt_3186_req
      -- 
    phi_stmt_3186_req_8882_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3186_req_8882_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(111), ack => phi_stmt_3186_req_0); -- 
    convTransposeD_cp_element_group_111: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_111"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7576_elements(109) & convTransposeD_CP_7576_elements(110);
      gj_convTransposeD_cp_element_group_111 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7576_elements(111), clk => clk, reset => reset); --
    end block;
    -- CP-element group 112:  join  transition  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	111 
    -- CP-element group 112: 	108 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	113 
    -- CP-element group 112:  members (1) 
      -- CP-element group 112: 	 branch_block_stmt_2745/ifx_xthen83_ifx_xend_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_112: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_112"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7576_elements(111) & convTransposeD_CP_7576_elements(108);
      gj_convTransposeD_cp_element_group_112 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7576_elements(112), clk => clk, reset => reset); --
    end block;
    -- CP-element group 113:  merge  fork  transition  place  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	105 
    -- CP-element group 113: 	112 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	114 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (2) 
      -- CP-element group 113: 	 branch_block_stmt_2745/merge_stmt_3179_PhiReqMerge
      -- CP-element group 113: 	 branch_block_stmt_2745/merge_stmt_3179_PhiAck/$entry
      -- 
    convTransposeD_CP_7576_elements(113) <= OrReduce(convTransposeD_CP_7576_elements(105) & convTransposeD_CP_7576_elements(112));
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	113 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	116 
    -- CP-element group 114:  members (1) 
      -- CP-element group 114: 	 branch_block_stmt_2745/merge_stmt_3179_PhiAck/phi_stmt_3180_ack
      -- 
    phi_stmt_3180_ack_8887_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3180_ack_0, ack => convTransposeD_CP_7576_elements(114)); -- 
    -- CP-element group 115:  transition  input  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	116 
    -- CP-element group 115:  members (1) 
      -- CP-element group 115: 	 branch_block_stmt_2745/merge_stmt_3179_PhiAck/phi_stmt_3186_ack
      -- 
    phi_stmt_3186_ack_8888_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3186_ack_0, ack => convTransposeD_CP_7576_elements(115)); -- 
    -- CP-element group 116:  join  fork  transition  place  output  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	114 
    -- CP-element group 116: 	115 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	69 
    -- CP-element group 116: 	70 
    -- CP-element group 116:  members (10) 
      -- CP-element group 116: 	 branch_block_stmt_2745/merge_stmt_3179__exit__
      -- CP-element group 116: 	 branch_block_stmt_2745/assign_stmt_3197_to_assign_stmt_3202__entry__
      -- CP-element group 116: 	 branch_block_stmt_2745/assign_stmt_3197_to_assign_stmt_3202/$entry
      -- CP-element group 116: 	 branch_block_stmt_2745/assign_stmt_3197_to_assign_stmt_3202/type_cast_3196_sample_start_
      -- CP-element group 116: 	 branch_block_stmt_2745/assign_stmt_3197_to_assign_stmt_3202/type_cast_3196_update_start_
      -- CP-element group 116: 	 branch_block_stmt_2745/assign_stmt_3197_to_assign_stmt_3202/type_cast_3196_Sample/$entry
      -- CP-element group 116: 	 branch_block_stmt_2745/assign_stmt_3197_to_assign_stmt_3202/type_cast_3196_Sample/rr
      -- CP-element group 116: 	 branch_block_stmt_2745/assign_stmt_3197_to_assign_stmt_3202/type_cast_3196_Update/$entry
      -- CP-element group 116: 	 branch_block_stmt_2745/assign_stmt_3197_to_assign_stmt_3202/type_cast_3196_Update/cr
      -- CP-element group 116: 	 branch_block_stmt_2745/merge_stmt_3179_PhiAck/$exit
      -- 
    rr_8564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(116), ack => type_cast_3196_inst_req_0); -- 
    cr_8569_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8569_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7576_elements(116), ack => type_cast_3196_inst_req_1); -- 
    convTransposeD_cp_element_group_116: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_116"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7576_elements(114) & convTransposeD_CP_7576_elements(115);
      gj_convTransposeD_cp_element_group_116 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7576_elements(116), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i32_i32_2977_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2998_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_3058_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_3089_wire : std_logic_vector(31 downto 0);
    signal LOAD_padding_2833_data_0 : std_logic_vector(7 downto 0);
    signal LOAD_padding_2833_word_address_0 : std_logic_vector(0 downto 0);
    signal R_idxprom65_3100_resized : std_logic_vector(13 downto 0);
    signal R_idxprom65_3100_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_3069_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_3069_scaled : std_logic_vector(13 downto 0);
    signal add21_3040 : std_logic_vector(31 downto 0);
    signal add29_2938 : std_logic_vector(31 downto 0);
    signal add40_2953 : std_logic_vector(31 downto 0);
    signal add55_3010 : std_logic_vector(31 downto 0);
    signal add57_3045 : std_logic_vector(31 downto 0);
    signal add70_3118 : std_logic_vector(31 downto 0);
    signal add_2923 : std_logic_vector(31 downto 0);
    signal array_obj_ref_3070_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3070_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3070_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3070_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3070_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3070_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3101_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3101_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3101_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3101_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3101_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3101_root_address : std_logic_vector(13 downto 0);
    signal arrayidx66_3103 : std_logic_vector(31 downto 0);
    signal arrayidx_3072 : std_logic_vector(31 downto 0);
    signal call_2748 : std_logic_vector(15 downto 0);
    signal cmp81_3154 : std_logic_vector(0 downto 0);
    signal cmp92_3202 : std_logic_vector(0 downto 0);
    signal cmp_3123 : std_logic_vector(0 downto 0);
    signal conv13105_3035 : std_logic_vector(31 downto 0);
    signal conv16_2908 : std_logic_vector(31 downto 0);
    signal conv19_2913 : std_logic_vector(31 downto 0);
    signal conv26_2819 : std_logic_vector(31 downto 0);
    signal conv31_2838 : std_logic_vector(31 downto 0);
    signal conv37_2852 : std_logic_vector(31 downto 0);
    signal conv4_2793 : std_logic_vector(15 downto 0);
    signal conv50_2979 : std_logic_vector(31 downto 0);
    signal conv53_3000 : std_logic_vector(31 downto 0);
    signal conv69_3112 : std_logic_vector(31 downto 0);
    signal conv79_3149 : std_logic_vector(31 downto 0);
    signal conv88_3177 : std_logic_vector(15 downto 0);
    signal conv90_3197 : std_logic_vector(31 downto 0);
    signal conv_2771 : std_logic_vector(15 downto 0);
    signal div3_2789 : std_logic_vector(31 downto 0);
    signal div87_3173 : std_logic_vector(31 downto 0);
    signal div_2767 : std_logic_vector(31 downto 0);
    signal iNsTr_10_2884 : std_logic_vector(31 downto 0);
    signal iNsTr_2_2757 : std_logic_vector(31 downto 0);
    signal iNsTr_3_2779 : std_logic_vector(31 downto 0);
    signal iNsTr_4_2801 : std_logic_vector(31 downto 0);
    signal iNsTr_5_2811 : std_logic_vector(31 downto 0);
    signal iNsTr_6_2827 : std_logic_vector(31 downto 0);
    signal iNsTr_7_2844 : std_logic_vector(31 downto 0);
    signal iNsTr_8_2860 : std_logic_vector(31 downto 0);
    signal iNsTr_9_2872 : std_logic_vector(31 downto 0);
    signal idxprom65_3096 : std_logic_vector(63 downto 0);
    signal idxprom_3065 : std_logic_vector(63 downto 0);
    signal inc85_3167 : std_logic_vector(15 downto 0);
    signal inc_3144 : std_logic_vector(15 downto 0);
    signal indvar_3018 : std_logic_vector(15 downto 0);
    signal indvarx_xnext_3136 : std_logic_vector(15 downto 0);
    signal input_dim0x_x0_3186 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2x_xph_2897 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1x_xph_2891 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_3180 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_3031 : std_logic_vector(15 downto 0);
    signal mul20_2928 : std_logic_vector(31 downto 0);
    signal mul27_2933 : std_logic_vector(31 downto 0);
    signal mul38_2948 : std_logic_vector(31 downto 0);
    signal mul54_3005 : std_logic_vector(31 downto 0);
    signal mul56_3015 : std_logic_vector(31 downto 0);
    signal mul_2918 : std_logic_vector(31 downto 0);
    signal ptr_deref_2760_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2760_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2760_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2760_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2760_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2782_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2782_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2782_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2782_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2782_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2804_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2804_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2804_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2804_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2804_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2814_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2814_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2814_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2814_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2814_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2830_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2830_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2830_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2830_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2830_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2847_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2847_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2847_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2847_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2847_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2863_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2863_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2863_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2863_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2863_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2875_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2875_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2875_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2875_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2875_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2887_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2887_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2887_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2887_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2887_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_3075_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_3075_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3075_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3075_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3075_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3105_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_3105_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3105_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3105_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_3105_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3105_word_offset_0 : std_logic_vector(13 downto 0);
    signal sext106_2991 : std_logic_vector(31 downto 0);
    signal sext108_3051 : std_logic_vector(31 downto 0);
    signal sext109_3082 : std_logic_vector(31 downto 0);
    signal sext_2970 : std_logic_vector(31 downto 0);
    signal shr64_3091 : std_logic_vector(31 downto 0);
    signal shr_3060 : std_logic_vector(31 downto 0);
    signal sub32_2985 : std_logic_vector(31 downto 0);
    signal sub43_2958 : std_logic_vector(31 downto 0);
    signal sub44_2964 : std_logic_vector(31 downto 0);
    signal sub_2943 : std_logic_vector(31 downto 0);
    signal tmp14_2805 : std_logic_vector(31 downto 0);
    signal tmp25_2815 : std_logic_vector(7 downto 0);
    signal tmp28_2831 : std_logic_vector(31 downto 0);
    signal tmp2_2783 : std_logic_vector(31 downto 0);
    signal tmp30_2834 : std_logic_vector(7 downto 0);
    signal tmp36_2848 : std_logic_vector(7 downto 0);
    signal tmp39_2864 : std_logic_vector(31 downto 0);
    signal tmp48_2876 : std_logic_vector(31 downto 0);
    signal tmp51_2888 : std_logic_vector(31 downto 0);
    signal tmp61_3076 : std_logic_vector(63 downto 0);
    signal tmp_2761 : std_logic_vector(31 downto 0);
    signal type_cast_2765_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2787_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2894_wire : std_logic_vector(15 downto 0);
    signal type_cast_2896_wire : std_logic_vector(15 downto 0);
    signal type_cast_2900_wire : std_logic_vector(15 downto 0);
    signal type_cast_2902_wire : std_logic_vector(15 downto 0);
    signal type_cast_2906_wire : std_logic_vector(31 downto 0);
    signal type_cast_2911_wire : std_logic_vector(31 downto 0);
    signal type_cast_2962_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2968_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2973_wire : std_logic_vector(31 downto 0);
    signal type_cast_2976_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2983_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2989_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2994_wire : std_logic_vector(31 downto 0);
    signal type_cast_2997_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3022_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3024_wire : std_logic_vector(15 downto 0);
    signal type_cast_3029_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3049_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3054_wire : std_logic_vector(31 downto 0);
    signal type_cast_3057_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3063_wire : std_logic_vector(63 downto 0);
    signal type_cast_3080_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3085_wire : std_logic_vector(31 downto 0);
    signal type_cast_3088_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3094_wire : std_logic_vector(63 downto 0);
    signal type_cast_3110_wire : std_logic_vector(31 downto 0);
    signal type_cast_3116_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3134_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3142_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3147_wire : std_logic_vector(31 downto 0);
    signal type_cast_3165_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3171_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3183_wire : std_logic_vector(15 downto 0);
    signal type_cast_3185_wire : std_logic_vector(15 downto 0);
    signal type_cast_3189_wire : std_logic_vector(15 downto 0);
    signal type_cast_3191_wire : std_logic_vector(15 downto 0);
    signal type_cast_3195_wire : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    LOAD_padding_2833_word_address_0 <= "0";
    array_obj_ref_3070_constant_part_of_offset <= "00000000000000";
    array_obj_ref_3070_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_3070_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_3070_resized_base_address <= "00000000000000";
    array_obj_ref_3101_constant_part_of_offset <= "00000000000000";
    array_obj_ref_3101_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_3101_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_3101_resized_base_address <= "00000000000000";
    iNsTr_10_2884 <= "00000000000000000000000000000100";
    iNsTr_2_2757 <= "00000000000000000000000000000011";
    iNsTr_3_2779 <= "00000000000000000000000000000100";
    iNsTr_4_2801 <= "00000000000000000000000000000101";
    iNsTr_5_2811 <= "00000000000000000000000000000000";
    iNsTr_6_2827 <= "00000000000000000000000000000100";
    iNsTr_7_2844 <= "00000000000000000000000000000001";
    iNsTr_8_2860 <= "00000000000000000000000000000101";
    iNsTr_9_2872 <= "00000000000000000000000000000101";
    ptr_deref_2760_word_offset_0 <= "0000000";
    ptr_deref_2782_word_offset_0 <= "0000000";
    ptr_deref_2804_word_offset_0 <= "0000000";
    ptr_deref_2814_word_offset_0 <= "0";
    ptr_deref_2830_word_offset_0 <= "0000000";
    ptr_deref_2847_word_offset_0 <= "0";
    ptr_deref_2863_word_offset_0 <= "0000000";
    ptr_deref_2875_word_offset_0 <= "0000000";
    ptr_deref_2887_word_offset_0 <= "0000000";
    ptr_deref_3075_word_offset_0 <= "00000000000000";
    ptr_deref_3105_word_offset_0 <= "00000000000000";
    type_cast_2765_wire_constant <= "00000000000000000000000000000001";
    type_cast_2787_wire_constant <= "00000000000000000000000000000001";
    type_cast_2962_wire_constant <= "00000000000000000000000000010000";
    type_cast_2968_wire_constant <= "11111111111111110000000000000000";
    type_cast_2976_wire_constant <= "00000000000000000000000000010000";
    type_cast_2983_wire_constant <= "00000000000000000000000000010000";
    type_cast_2989_wire_constant <= "11111111111111110000000000000000";
    type_cast_2997_wire_constant <= "00000000000000000000000000010000";
    type_cast_3022_wire_constant <= "0000000000000000";
    type_cast_3029_wire_constant <= "0000000000000100";
    type_cast_3049_wire_constant <= "00000000000000000000000000010000";
    type_cast_3057_wire_constant <= "00000000000000000000000000010010";
    type_cast_3080_wire_constant <= "00000000000000000000000000010000";
    type_cast_3088_wire_constant <= "00000000000000000000000000010010";
    type_cast_3116_wire_constant <= "00000000000000000000000000000100";
    type_cast_3134_wire_constant <= "0000000000000001";
    type_cast_3142_wire_constant <= "0000000000000001";
    type_cast_3165_wire_constant <= "0000000000000001";
    type_cast_3171_wire_constant <= "00000000000000000000000000000001";
    phi_stmt_2891: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2894_wire & type_cast_2896_wire;
      req <= phi_stmt_2891_req_0 & phi_stmt_2891_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2891",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2891_ack_0,
          idata => idata,
          odata => input_dim1x_x1x_xph_2891,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2891
    phi_stmt_2897: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2900_wire & type_cast_2902_wire;
      req <= phi_stmt_2897_req_0 & phi_stmt_2897_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2897",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2897_ack_0,
          idata => idata,
          odata => input_dim0x_x2x_xph_2897,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2897
    phi_stmt_3018: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3022_wire_constant & type_cast_3024_wire;
      req <= phi_stmt_3018_req_0 & phi_stmt_3018_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3018",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3018_ack_0,
          idata => idata,
          odata => indvar_3018,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3018
    phi_stmt_3180: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3183_wire & type_cast_3185_wire;
      req <= phi_stmt_3180_req_0 & phi_stmt_3180_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3180",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3180_ack_0,
          idata => idata,
          odata => input_dim1x_x2_3180,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3180
    phi_stmt_3186: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3189_wire & type_cast_3191_wire;
      req <= phi_stmt_3186_req_0 & phi_stmt_3186_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3186",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3186_ack_0,
          idata => idata,
          odata => input_dim0x_x0_3186,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3186
    addr_of_3071_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_3071_final_reg_req_0;
      addr_of_3071_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_3071_final_reg_req_1;
      addr_of_3071_final_reg_ack_1<= rack(0);
      addr_of_3071_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_3071_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_3070_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_3072,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_3102_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_3102_final_reg_req_0;
      addr_of_3102_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_3102_final_reg_req_1;
      addr_of_3102_final_reg_ack_1<= rack(0);
      addr_of_3102_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_3102_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_3101_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx66_3103,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2770_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2770_inst_req_0;
      type_cast_2770_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2770_inst_req_1;
      type_cast_2770_inst_ack_1<= rack(0);
      type_cast_2770_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2770_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div_2767,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_2771,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2792_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2792_inst_req_0;
      type_cast_2792_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2792_inst_req_1;
      type_cast_2792_inst_ack_1<= rack(0);
      type_cast_2792_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2792_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div3_2789,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv4_2793,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2818_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2818_inst_req_0;
      type_cast_2818_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2818_inst_req_1;
      type_cast_2818_inst_ack_1<= rack(0);
      type_cast_2818_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2818_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp25_2815,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv26_2819,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2837_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2837_inst_req_0;
      type_cast_2837_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2837_inst_req_1;
      type_cast_2837_inst_ack_1<= rack(0);
      type_cast_2837_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2837_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp30_2834,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv31_2838,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2851_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2851_inst_req_0;
      type_cast_2851_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2851_inst_req_1;
      type_cast_2851_inst_ack_1<= rack(0);
      type_cast_2851_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2851_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp36_2848,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv37_2852,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2894_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2894_inst_req_0;
      type_cast_2894_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2894_inst_req_1;
      type_cast_2894_inst_ack_1<= rack(0);
      type_cast_2894_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2894_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv4_2793,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2894_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2896_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2896_inst_req_0;
      type_cast_2896_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2896_inst_req_1;
      type_cast_2896_inst_ack_1<= rack(0);
      type_cast_2896_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2896_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_3180,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2896_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2900_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2900_inst_req_0;
      type_cast_2900_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2900_inst_req_1;
      type_cast_2900_inst_ack_1<= rack(0);
      type_cast_2900_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2900_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv_2771,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2900_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2902_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2902_inst_req_0;
      type_cast_2902_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2902_inst_req_1;
      type_cast_2902_inst_ack_1<= rack(0);
      type_cast_2902_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2902_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x0_3186,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2902_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2907_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2907_inst_req_0;
      type_cast_2907_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2907_inst_req_1;
      type_cast_2907_inst_ack_1<= rack(0);
      type_cast_2907_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2907_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2906_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv16_2908,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2912_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2912_inst_req_0;
      type_cast_2912_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2912_inst_req_1;
      type_cast_2912_inst_ack_1<= rack(0);
      type_cast_2912_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2912_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2911_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv19_2913,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2973_inst
    process(sext_2970) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext_2970(31 downto 0);
      type_cast_2973_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2978_inst
    process(ASHR_i32_i32_2977_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2977_wire(31 downto 0);
      conv50_2979 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2994_inst
    process(sext106_2991) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext106_2991(31 downto 0);
      type_cast_2994_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2999_inst
    process(ASHR_i32_i32_2998_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2998_wire(31 downto 0);
      conv53_3000 <= tmp_var; -- 
    end process;
    type_cast_3024_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3024_inst_req_0;
      type_cast_3024_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3024_inst_req_1;
      type_cast_3024_inst_ack_1<= rack(0);
      type_cast_3024_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3024_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_3136,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3024_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3034_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3034_inst_req_0;
      type_cast_3034_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3034_inst_req_1;
      type_cast_3034_inst_ack_1<= rack(0);
      type_cast_3034_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3034_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_3031,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv13105_3035,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3054_inst
    process(sext108_3051) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext108_3051(31 downto 0);
      type_cast_3054_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3059_inst
    process(ASHR_i32_i32_3058_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3058_wire(31 downto 0);
      shr_3060 <= tmp_var; -- 
    end process;
    type_cast_3064_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3064_inst_req_0;
      type_cast_3064_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3064_inst_req_1;
      type_cast_3064_inst_ack_1<= rack(0);
      type_cast_3064_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3064_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3063_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_3065,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3085_inst
    process(sext109_3082) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext109_3082(31 downto 0);
      type_cast_3085_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3090_inst
    process(ASHR_i32_i32_3089_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3089_wire(31 downto 0);
      shr64_3091 <= tmp_var; -- 
    end process;
    type_cast_3095_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3095_inst_req_0;
      type_cast_3095_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3095_inst_req_1;
      type_cast_3095_inst_ack_1<= rack(0);
      type_cast_3095_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3095_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3094_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom65_3096,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3111_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3111_inst_req_0;
      type_cast_3111_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3111_inst_req_1;
      type_cast_3111_inst_ack_1<= rack(0);
      type_cast_3111_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3111_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3110_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv69_3112,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3148_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3148_inst_req_0;
      type_cast_3148_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3148_inst_req_1;
      type_cast_3148_inst_ack_1<= rack(0);
      type_cast_3148_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3148_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3147_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv79_3149,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3176_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3176_inst_req_0;
      type_cast_3176_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3176_inst_req_1;
      type_cast_3176_inst_ack_1<= rack(0);
      type_cast_3176_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3176_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div87_3173,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv88_3177,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3183_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3183_inst_req_0;
      type_cast_3183_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3183_inst_req_1;
      type_cast_3183_inst_ack_1<= rack(0);
      type_cast_3183_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3183_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv88_3177,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3183_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3185_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3185_inst_req_0;
      type_cast_3185_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3185_inst_req_1;
      type_cast_3185_inst_ack_1<= rack(0);
      type_cast_3185_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3185_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc_3144,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3185_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3189_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3189_inst_req_0;
      type_cast_3189_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3189_inst_req_1;
      type_cast_3189_inst_ack_1<= rack(0);
      type_cast_3189_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3189_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc85_3167,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3189_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3191_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3191_inst_req_0;
      type_cast_3191_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3191_inst_req_1;
      type_cast_3191_inst_ack_1<= rack(0);
      type_cast_3191_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3191_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x2x_xph_2897,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3191_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3196_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3196_inst_req_0;
      type_cast_3196_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3196_inst_req_1;
      type_cast_3196_inst_ack_1<= rack(0);
      type_cast_3196_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3196_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3195_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv90_3197,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence LOAD_padding_2833_gather_scatter
    process(LOAD_padding_2833_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_padding_2833_data_0;
      ov(7 downto 0) := iv;
      tmp30_2834 <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3070_index_1_rename
    process(R_idxprom_3069_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_3069_resized;
      ov(13 downto 0) := iv;
      R_idxprom_3069_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3070_index_1_resize
    process(idxprom_3065) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_3065;
      ov := iv(13 downto 0);
      R_idxprom_3069_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3070_root_address_inst
    process(array_obj_ref_3070_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_3070_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_3070_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3101_index_1_rename
    process(R_idxprom65_3100_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom65_3100_resized;
      ov(13 downto 0) := iv;
      R_idxprom65_3100_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3101_index_1_resize
    process(idxprom65_3096) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom65_3096;
      ov := iv(13 downto 0);
      R_idxprom65_3100_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3101_root_address_inst
    process(array_obj_ref_3101_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_3101_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_3101_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2760_addr_0
    process(ptr_deref_2760_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2760_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2760_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2760_base_resize
    process(iNsTr_2_2757) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_2_2757;
      ov := iv(6 downto 0);
      ptr_deref_2760_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2760_gather_scatter
    process(ptr_deref_2760_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2760_data_0;
      ov(31 downto 0) := iv;
      tmp_2761 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2760_root_address_inst
    process(ptr_deref_2760_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2760_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2760_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2782_addr_0
    process(ptr_deref_2782_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2782_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2782_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2782_base_resize
    process(iNsTr_3_2779) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_3_2779;
      ov := iv(6 downto 0);
      ptr_deref_2782_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2782_gather_scatter
    process(ptr_deref_2782_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2782_data_0;
      ov(31 downto 0) := iv;
      tmp2_2783 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2782_root_address_inst
    process(ptr_deref_2782_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2782_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2782_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2804_addr_0
    process(ptr_deref_2804_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2804_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2804_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2804_base_resize
    process(iNsTr_4_2801) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_4_2801;
      ov := iv(6 downto 0);
      ptr_deref_2804_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2804_gather_scatter
    process(ptr_deref_2804_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2804_data_0;
      ov(31 downto 0) := iv;
      tmp14_2805 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2804_root_address_inst
    process(ptr_deref_2804_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2804_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2804_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2814_addr_0
    process(ptr_deref_2814_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2814_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_2814_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2814_base_resize
    process(iNsTr_5_2811) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_5_2811;
      ov := iv(0 downto 0);
      ptr_deref_2814_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2814_gather_scatter
    process(ptr_deref_2814_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2814_data_0;
      ov(7 downto 0) := iv;
      tmp25_2815 <= ov(7 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2814_root_address_inst
    process(ptr_deref_2814_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2814_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_2814_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2830_addr_0
    process(ptr_deref_2830_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2830_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2830_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2830_base_resize
    process(iNsTr_6_2827) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_6_2827;
      ov := iv(6 downto 0);
      ptr_deref_2830_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2830_gather_scatter
    process(ptr_deref_2830_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2830_data_0;
      ov(31 downto 0) := iv;
      tmp28_2831 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2830_root_address_inst
    process(ptr_deref_2830_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2830_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2830_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2847_addr_0
    process(ptr_deref_2847_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2847_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_2847_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2847_base_resize
    process(iNsTr_7_2844) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_7_2844;
      ov := iv(0 downto 0);
      ptr_deref_2847_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2847_gather_scatter
    process(ptr_deref_2847_data_0) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2847_data_0;
      ov(7 downto 0) := iv;
      tmp36_2848 <= ov(7 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2847_root_address_inst
    process(ptr_deref_2847_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2847_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_2847_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2863_addr_0
    process(ptr_deref_2863_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2863_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2863_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2863_base_resize
    process(iNsTr_8_2860) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_8_2860;
      ov := iv(6 downto 0);
      ptr_deref_2863_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2863_gather_scatter
    process(ptr_deref_2863_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2863_data_0;
      ov(31 downto 0) := iv;
      tmp39_2864 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2863_root_address_inst
    process(ptr_deref_2863_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2863_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2863_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2875_addr_0
    process(ptr_deref_2875_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2875_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2875_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2875_base_resize
    process(iNsTr_9_2872) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_9_2872;
      ov := iv(6 downto 0);
      ptr_deref_2875_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2875_gather_scatter
    process(ptr_deref_2875_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2875_data_0;
      ov(31 downto 0) := iv;
      tmp48_2876 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2875_root_address_inst
    process(ptr_deref_2875_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2875_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2875_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2887_addr_0
    process(ptr_deref_2887_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2887_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2887_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2887_base_resize
    process(iNsTr_10_2884) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_10_2884;
      ov := iv(6 downto 0);
      ptr_deref_2887_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2887_gather_scatter
    process(ptr_deref_2887_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2887_data_0;
      ov(31 downto 0) := iv;
      tmp51_2888 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2887_root_address_inst
    process(ptr_deref_2887_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2887_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2887_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3075_addr_0
    process(ptr_deref_3075_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3075_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_3075_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3075_base_resize
    process(arrayidx_3072) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_3072;
      ov := iv(13 downto 0);
      ptr_deref_3075_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3075_gather_scatter
    process(ptr_deref_3075_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3075_data_0;
      ov(63 downto 0) := iv;
      tmp61_3076 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3075_root_address_inst
    process(ptr_deref_3075_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3075_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_3075_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3105_addr_0
    process(ptr_deref_3105_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3105_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_3105_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3105_base_resize
    process(arrayidx66_3103) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx66_3103;
      ov := iv(13 downto 0);
      ptr_deref_3105_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3105_gather_scatter
    process(tmp61_3076) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp61_3076;
      ov(63 downto 0) := iv;
      ptr_deref_3105_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3105_root_address_inst
    process(ptr_deref_3105_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3105_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_3105_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_3124_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_3123;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3124_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3124_branch_req_0,
          ack0 => if_stmt_3124_branch_ack_0,
          ack1 => if_stmt_3124_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3155_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp81_3154;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3155_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3155_branch_req_0,
          ack0 => if_stmt_3155_branch_ack_0,
          ack1 => if_stmt_3155_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3203_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp92_3202;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3203_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3203_branch_req_0,
          ack0 => if_stmt_3203_branch_ack_0,
          ack1 => if_stmt_3203_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_3135_inst
    process(indvar_3018) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_3018, type_cast_3134_wire_constant, tmp_var);
      indvarx_xnext_3136 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3143_inst
    process(input_dim1x_x1x_xph_2891) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_2891, type_cast_3142_wire_constant, tmp_var);
      inc_3144 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3166_inst
    process(input_dim0x_x2x_xph_2897) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim0x_x2x_xph_2897, type_cast_3165_wire_constant, tmp_var);
      inc85_3167 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2922_inst
    process(mul_2918, conv16_2908) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul_2918, conv16_2908, tmp_var);
      add_2923 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2937_inst
    process(mul27_2933, tmp28_2831) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul27_2933, tmp28_2831, tmp_var);
      add29_2938 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2952_inst
    process(mul38_2948, tmp39_2864) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul38_2948, tmp39_2864, tmp_var);
      add40_2953 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2969_inst
    process(sub44_2964) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub44_2964, type_cast_2968_wire_constant, tmp_var);
      sext_2970 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2990_inst
    process(sub32_2985) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub32_2985, type_cast_2989_wire_constant, tmp_var);
      sext106_2991 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3009_inst
    process(conv50_2979, mul54_3005) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv50_2979, mul54_3005, tmp_var);
      add55_3010 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3039_inst
    process(mul20_2928, conv13105_3035) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul20_2928, conv13105_3035, tmp_var);
      add21_3040 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3044_inst
    process(mul56_3015, conv13105_3035) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul56_3015, conv13105_3035, tmp_var);
      add57_3045 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3117_inst
    process(conv69_3112) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv69_3112, type_cast_3116_wire_constant, tmp_var);
      add70_3118 <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2977_inst
    process(type_cast_2973_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2973_wire, type_cast_2976_wire_constant, tmp_var);
      ASHR_i32_i32_2977_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2998_inst
    process(type_cast_2994_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2994_wire, type_cast_2997_wire_constant, tmp_var);
      ASHR_i32_i32_2998_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3058_inst
    process(type_cast_3054_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3054_wire, type_cast_3057_wire_constant, tmp_var);
      ASHR_i32_i32_3058_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3089_inst
    process(type_cast_3085_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3085_wire, type_cast_3088_wire_constant, tmp_var);
      ASHR_i32_i32_3089_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_3153_inst
    process(conv79_3149, tmp2_2783) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv79_3149, tmp2_2783, tmp_var);
      cmp81_3154 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_3201_inst
    process(conv90_3197, tmp_2761) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv90_3197, tmp_2761, tmp_var);
      cmp92_3202 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2766_inst
    process(tmp_2761) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp_2761, type_cast_2765_wire_constant, tmp_var);
      div_2767 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2788_inst
    process(tmp2_2783) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp2_2783, type_cast_2787_wire_constant, tmp_var);
      div3_2789 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_3172_inst
    process(tmp2_2783) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp2_2783, type_cast_3171_wire_constant, tmp_var);
      div87_3173 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_3030_inst
    process(indvar_3018) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_3018, type_cast_3029_wire_constant, tmp_var);
      input_dim2x_x1_3031 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2917_inst
    process(tmp2_2783, conv19_2913) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp2_2783, conv19_2913, tmp_var);
      mul_2918 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2927_inst
    process(add_2923, tmp14_2805) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add_2923, tmp14_2805, tmp_var);
      mul20_2928 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2932_inst
    process(conv26_2819, conv19_2913) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv26_2819, conv19_2913, tmp_var);
      mul27_2933 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2947_inst
    process(conv37_2852, conv16_2908) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv37_2852, conv16_2908, tmp_var);
      mul38_2948 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3004_inst
    process(tmp51_2888, conv53_3000) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp51_2888, conv53_3000, tmp_var);
      mul54_3005 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3014_inst
    process(add55_3010, tmp48_2876) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add55_3010, tmp48_2876, tmp_var);
      mul56_3015 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2963_inst
    process(sub43_2958) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(sub43_2958, type_cast_2962_wire_constant, tmp_var);
      sub44_2964 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2984_inst
    process(sub_2943) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(sub_2943, type_cast_2983_wire_constant, tmp_var);
      sub32_2985 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_3050_inst
    process(add21_3040) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add21_3040, type_cast_3049_wire_constant, tmp_var);
      sext108_3051 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_3081_inst
    process(add57_3045) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add57_3045, type_cast_3080_wire_constant, tmp_var);
      sext109_3082 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_2942_inst
    process(add29_2938, conv31_2838) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(add29_2938, conv31_2838, tmp_var);
      sub_2943 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_2957_inst
    process(add40_2953, conv31_2838) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(add40_2953, conv31_2838, tmp_var);
      sub43_2958 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_3122_inst
    process(add70_3118, tmp14_2805) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add70_3118, tmp14_2805, tmp_var);
      cmp_3123 <= tmp_var; --
    end process;
    -- shared split operator group (35) : array_obj_ref_3070_index_offset 
    ApIntAdd_group_35: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_3069_scaled;
      array_obj_ref_3070_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_3070_index_offset_req_0;
      array_obj_ref_3070_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_3070_index_offset_req_1;
      array_obj_ref_3070_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_35_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_35_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_35",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 35
    -- shared split operator group (36) : array_obj_ref_3101_index_offset 
    ApIntAdd_group_36: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom65_3100_scaled;
      array_obj_ref_3101_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_3101_index_offset_req_0;
      array_obj_ref_3101_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_3101_index_offset_req_1;
      array_obj_ref_3101_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_36_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_36_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_36",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 36
    -- unary operator type_cast_2906_inst
    process(input_dim1x_x1x_xph_2891) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim1x_x1x_xph_2891, tmp_var);
      type_cast_2906_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2911_inst
    process(input_dim0x_x2x_xph_2897) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim0x_x2x_xph_2897, tmp_var);
      type_cast_2911_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3063_inst
    process(shr_3060) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr_3060, tmp_var);
      type_cast_3063_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3094_inst
    process(shr64_3091) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr64_3091, tmp_var);
      type_cast_3094_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3110_inst
    process(input_dim2x_x1_3031) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim2x_x1_3031, tmp_var);
      type_cast_3110_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3147_inst
    process(inc_3144) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc_3144, tmp_var);
      type_cast_3147_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3195_inst
    process(input_dim0x_x0_3186) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim0x_x0_3186, tmp_var);
      type_cast_3195_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : LOAD_padding_2833_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_padding_2833_load_0_req_0;
      LOAD_padding_2833_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_padding_2833_load_0_req_1;
      LOAD_padding_2833_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_padding_2833_word_address_0;
      LOAD_padding_2833_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_7_lr_req(0),
          mack => memory_space_7_lr_ack(0),
          maddr => memory_space_7_lr_addr(0 downto 0),
          mtag => memory_space_7_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 8,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_7_lc_req(0),
          mack => memory_space_7_lc_ack(0),
          mdata => memory_space_7_lc_data(7 downto 0),
          mtag => memory_space_7_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_2760_load_0 ptr_deref_2782_load_0 ptr_deref_2804_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(20 downto 0);
      signal data_out: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_2760_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_2782_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2804_load_0_req_0;
      ptr_deref_2760_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_2782_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2804_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_2760_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_2782_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2804_load_0_req_1;
      ptr_deref_2760_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_2782_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2804_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      LoadGroup1_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2760_word_address_0 & ptr_deref_2782_word_address_0 & ptr_deref_2804_word_address_0;
      ptr_deref_2760_data_0 <= data_out(95 downto 64);
      ptr_deref_2782_data_0 <= data_out(63 downto 32);
      ptr_deref_2804_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 7,
        num_reqs => 3,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(6 downto 0),
          mtag => memory_space_1_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 32,
        num_reqs => 3,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(31 downto 0),
          mtag => memory_space_1_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : ptr_deref_2814_load_0 ptr_deref_2847_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_2814_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2847_load_0_req_0;
      ptr_deref_2814_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2847_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_2814_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2847_load_0_req_1;
      ptr_deref_2814_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2847_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup2_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup2_gI: SplitGuardInterface generic map(name => "LoadGroup2_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2814_word_address_0 & ptr_deref_2847_word_address_0;
      ptr_deref_2814_data_0 <= data_out(15 downto 8);
      ptr_deref_2847_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup2", addr_width => 1,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_8_lr_req(0),
          mack => memory_space_8_lr_ack(0),
          maddr => memory_space_8_lr_addr(0 downto 0),
          mtag => memory_space_8_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup2 load-complete ",
        data_width => 8,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_8_lc_req(0),
          mack => memory_space_8_lc_ack(0),
          mdata => memory_space_8_lc_data(7 downto 0),
          mtag => memory_space_8_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared load operator group (3) : ptr_deref_2830_load_0 ptr_deref_2863_load_0 
    LoadGroup3: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_2830_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2863_load_0_req_0;
      ptr_deref_2830_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2863_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_2830_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2863_load_0_req_1;
      ptr_deref_2830_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2863_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup3_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup3_gI: SplitGuardInterface generic map(name => "LoadGroup3_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2830_word_address_0 & ptr_deref_2863_word_address_0;
      ptr_deref_2830_data_0 <= data_out(63 downto 32);
      ptr_deref_2863_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup3", addr_width => 7,
        num_reqs => 2,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(6 downto 0),
          mtag => memory_space_2_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup3 load-complete ",
        data_width => 32,
        num_reqs => 2,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(31 downto 0),
          mtag => memory_space_2_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 3
    -- shared load operator group (4) : ptr_deref_2875_load_0 ptr_deref_2887_load_0 
    LoadGroup4: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_2875_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2887_load_0_req_0;
      ptr_deref_2875_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2887_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_2875_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2887_load_0_req_1;
      ptr_deref_2875_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2887_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup4_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup4_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup4_gI: SplitGuardInterface generic map(name => "LoadGroup4_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2875_word_address_0 & ptr_deref_2887_word_address_0;
      ptr_deref_2875_data_0 <= data_out(63 downto 32);
      ptr_deref_2887_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup4", addr_width => 7,
        num_reqs => 2,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(6 downto 0),
          mtag => memory_space_3_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup4 load-complete ",
        data_width => 32,
        num_reqs => 2,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(31 downto 0),
          mtag => memory_space_3_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 4
    -- shared load operator group (5) : ptr_deref_3075_load_0 
    LoadGroup5: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_3075_load_0_req_0;
      ptr_deref_3075_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_3075_load_0_req_1;
      ptr_deref_3075_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup5_gI: SplitGuardInterface generic map(name => "LoadGroup5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_3075_word_address_0;
      ptr_deref_3075_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup5", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_4_lr_req(0),
          mack => memory_space_4_lr_ack(0),
          maddr => memory_space_4_lr_addr(13 downto 0),
          mtag => memory_space_4_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup5 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_4_lc_req(0),
          mack => memory_space_4_lc_ack(0),
          mdata => memory_space_4_lc_data(63 downto 0),
          mtag => memory_space_4_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 5
    -- shared store operator group (0) : ptr_deref_3105_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_3105_store_0_req_0;
      ptr_deref_3105_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_3105_store_0_req_1;
      ptr_deref_3105_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_3105_word_address_0;
      data_in <= ptr_deref_3105_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_6_sr_req(0),
          mack => memory_space_6_sr_ack(0),
          maddr => memory_space_6_sr_addr(13 downto 0),
          mdata => memory_space_6_sr_data(63 downto 0),
          mtag => memory_space_6_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_6_sc_req(0),
          mack => memory_space_6_sc_ack(0),
          mtag => memory_space_6_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block3_start_2747_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block3_start_2747_inst_req_0;
      RPIPE_Block3_start_2747_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block3_start_2747_inst_req_1;
      RPIPE_Block3_start_2747_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call_2748 <= data_out(15 downto 0);
      Block3_start_read_0_gI: SplitGuardInterface generic map(name => "Block3_start_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block3_start_read_0: InputPortRevised -- 
        generic map ( name => "Block3_start_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block3_start_pipe_read_req(0),
          oack => Block3_start_pipe_read_ack(0),
          odata => Block3_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block3_done_3211_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block3_done_3211_inst_req_0;
      WPIPE_Block3_done_3211_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block3_done_3211_inst_req_1;
      WPIPE_Block3_done_3211_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= call_2748;
      Block3_done_write_0_gI: SplitGuardInterface generic map(name => "Block3_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block3_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block3_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block3_done_pipe_write_req(0),
          oack => Block3_done_pipe_write_ack(0),
          odata => Block3_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeD_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity sendOutput is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_6_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_6_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(2 downto 0);
    ConvTranspose_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity sendOutput;
architecture sendOutput_arch of sendOutput is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal sendOutput_CP_3122_start: Boolean;
  signal sendOutput_CP_3122_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal type_cast_1163_inst_req_0 : boolean;
  signal array_obj_ref_1192_index_offset_ack_1 : boolean;
  signal ptr_deref_1197_load_0_req_0 : boolean;
  signal ptr_deref_1106_load_0_ack_0 : boolean;
  signal if_stmt_1136_branch_req_0 : boolean;
  signal array_obj_ref_1192_index_offset_req_1 : boolean;
  signal ptr_deref_1197_load_0_ack_0 : boolean;
  signal ptr_deref_1094_load_0_ack_1 : boolean;
  signal type_cast_1163_inst_ack_0 : boolean;
  signal ptr_deref_1106_load_0_req_0 : boolean;
  signal ptr_deref_1094_load_0_ack_0 : boolean;
  signal ptr_deref_1106_load_0_ack_1 : boolean;
  signal type_cast_1201_inst_req_1 : boolean;
  signal ptr_deref_1094_load_0_req_0 : boolean;
  signal type_cast_1201_inst_req_0 : boolean;
  signal ptr_deref_1094_load_0_req_1 : boolean;
  signal type_cast_1163_inst_ack_1 : boolean;
  signal ptr_deref_1106_load_0_req_1 : boolean;
  signal type_cast_1231_inst_req_0 : boolean;
  signal type_cast_1231_inst_ack_0 : boolean;
  signal type_cast_1231_inst_req_1 : boolean;
  signal type_cast_1231_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1279_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1279_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1276_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1276_inst_ack_1 : boolean;
  signal type_cast_1271_inst_req_1 : boolean;
  signal type_cast_1271_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1279_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1279_inst_ack_0 : boolean;
  signal ptr_deref_1197_load_0_ack_1 : boolean;
  signal addr_of_1193_final_reg_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1273_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1273_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1282_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1282_inst_ack_0 : boolean;
  signal ptr_deref_1118_load_0_req_0 : boolean;
  signal type_cast_1221_inst_req_1 : boolean;
  signal type_cast_1221_inst_ack_1 : boolean;
  signal type_cast_1271_inst_ack_0 : boolean;
  signal ptr_deref_1118_load_0_ack_0 : boolean;
  signal type_cast_1211_inst_ack_0 : boolean;
  signal type_cast_1251_inst_ack_1 : boolean;
  signal type_cast_1251_inst_req_0 : boolean;
  signal type_cast_1251_inst_ack_0 : boolean;
  signal type_cast_1261_inst_req_1 : boolean;
  signal type_cast_1261_inst_ack_1 : boolean;
  signal addr_of_1193_final_reg_ack_1 : boolean;
  signal type_cast_1211_inst_ack_1 : boolean;
  signal type_cast_1271_inst_req_0 : boolean;
  signal type_cast_1261_inst_req_0 : boolean;
  signal type_cast_1241_inst_req_1 : boolean;
  signal type_cast_1241_inst_ack_1 : boolean;
  signal array_obj_ref_1192_index_offset_req_0 : boolean;
  signal ptr_deref_1118_load_0_req_1 : boolean;
  signal array_obj_ref_1192_index_offset_ack_0 : boolean;
  signal type_cast_1241_inst_req_0 : boolean;
  signal type_cast_1241_inst_ack_0 : boolean;
  signal type_cast_1251_inst_req_1 : boolean;
  signal type_cast_1163_inst_req_1 : boolean;
  signal addr_of_1193_final_reg_req_1 : boolean;
  signal type_cast_1261_inst_ack_0 : boolean;
  signal ptr_deref_1118_load_0_ack_1 : boolean;
  signal type_cast_1211_inst_req_1 : boolean;
  signal ptr_deref_1197_load_0_req_1 : boolean;
  signal if_stmt_1136_branch_ack_1 : boolean;
  signal type_cast_1201_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1282_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1282_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1273_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1273_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1276_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1276_inst_ack_0 : boolean;
  signal type_cast_1211_inst_req_0 : boolean;
  signal addr_of_1193_final_reg_req_0 : boolean;
  signal if_stmt_1136_branch_ack_0 : boolean;
  signal type_cast_1221_inst_req_0 : boolean;
  signal type_cast_1221_inst_ack_0 : boolean;
  signal type_cast_1201_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1285_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1285_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1285_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1285_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1288_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1288_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1288_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1288_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1291_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1291_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1291_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1291_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1294_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1294_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1294_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1294_inst_ack_1 : boolean;
  signal if_stmt_1308_branch_req_0 : boolean;
  signal if_stmt_1308_branch_ack_1 : boolean;
  signal if_stmt_1308_branch_ack_0 : boolean;
  signal phi_stmt_1180_req_0 : boolean;
  signal type_cast_1186_inst_req_0 : boolean;
  signal type_cast_1186_inst_ack_0 : boolean;
  signal type_cast_1186_inst_req_1 : boolean;
  signal type_cast_1186_inst_ack_1 : boolean;
  signal phi_stmt_1180_req_1 : boolean;
  signal phi_stmt_1180_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "sendOutput_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  sendOutput_CP_3122_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "sendOutput_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendOutput_CP_3122_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= sendOutput_CP_3122_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendOutput_CP_3122_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  sendOutput_CP_3122: Block -- control-path 
    signal sendOutput_CP_3122_elements: BooleanArray(66 downto 0);
    -- 
  begin -- 
    sendOutput_CP_3122_elements(0) <= sendOutput_CP_3122_start;
    sendOutput_CP_3122_symbol <= sendOutput_CP_3122_elements(66);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	3 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	5 
    -- CP-element group 0: 	6 
    -- CP-element group 0:  members (83) 
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1106_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1094_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1106_Sample/word_access_start/$entry
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1106_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1094_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1094_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1094_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1094_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1106_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/$entry
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1094_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1106_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1106_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1094_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135__entry__
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1118_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1106_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1094_Sample/word_access_start/$entry
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1106_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1094_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_1083/branch_block_stmt_1083__entry__
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1106_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1106_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1106_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1094_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1118_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1094_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1106_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1106_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1094_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1094_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1106_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1118_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1094_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1118_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1106_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1094_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1094_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1094_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1094_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1094_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1094_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1094_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1106_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1094_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1106_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1118_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_1083/$entry
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1118_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1094_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1118_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1118_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1118_Sample/word_access_start/$entry
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1118_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1118_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1118_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1118_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1118_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1106_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1094_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1106_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1118_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1118_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1118_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1106_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1118_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1106_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1118_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1106_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1118_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1106_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1118_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1118_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1106_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1118_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1118_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1106_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1118_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1106_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1094_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1094_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1118_sample_start_
      -- CP-element group 0: 	 $entry
      -- 
    rr_3235_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3235_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3122_elements(0), ack => ptr_deref_1106_load_0_req_0); -- 
    rr_3185_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3185_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3122_elements(0), ack => ptr_deref_1094_load_0_req_0); -- 
    cr_3196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3122_elements(0), ack => ptr_deref_1094_load_0_req_1); -- 
    cr_3246_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3246_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3122_elements(0), ack => ptr_deref_1106_load_0_req_1); -- 
    rr_3285_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3285_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3122_elements(0), ack => ptr_deref_1118_load_0_req_0); -- 
    cr_3296_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3296_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3122_elements(0), ack => ptr_deref_1118_load_0_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (5) 
      -- CP-element group 1: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1094_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1094_Sample/word_access_start/word_0/$exit
      -- CP-element group 1: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1094_Sample/word_access_start/$exit
      -- CP-element group 1: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1094_Sample/word_access_start/word_0/ra
      -- CP-element group 1: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1094_sample_completed_
      -- 
    ra_3186_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1094_load_0_ack_0, ack => sendOutput_CP_3122_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	7 
    -- CP-element group 2:  members (9) 
      -- CP-element group 2: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1094_Update/ptr_deref_1094_Merge/$exit
      -- CP-element group 2: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1094_Update/ptr_deref_1094_Merge/$entry
      -- CP-element group 2: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1094_Update/ptr_deref_1094_Merge/merge_req
      -- CP-element group 2: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1094_Update/ptr_deref_1094_Merge/merge_ack
      -- CP-element group 2: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1094_Update/word_access_complete/word_0/ca
      -- CP-element group 2: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1094_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1094_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1094_Update/word_access_complete/word_0/$exit
      -- CP-element group 2: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1094_Update/word_access_complete/$exit
      -- 
    ca_3197_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1094_load_0_ack_1, ack => sendOutput_CP_3122_elements(2)); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	0 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (5) 
      -- CP-element group 3: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1106_Sample/word_access_start/$exit
      -- CP-element group 3: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1106_Sample/word_access_start/word_0/ra
      -- CP-element group 3: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1106_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1106_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1106_Sample/word_access_start/word_0/$exit
      -- 
    ra_3236_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1106_load_0_ack_0, ack => sendOutput_CP_3122_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (9) 
      -- CP-element group 4: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1106_Update/word_access_complete/$exit
      -- CP-element group 4: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1106_Update/word_access_complete/word_0/ca
      -- CP-element group 4: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1106_Update/word_access_complete/word_0/$exit
      -- CP-element group 4: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1106_Update/ptr_deref_1106_Merge/$entry
      -- CP-element group 4: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1106_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1106_Update/ptr_deref_1106_Merge/merge_ack
      -- CP-element group 4: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1106_Update/ptr_deref_1106_Merge/$exit
      -- CP-element group 4: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1106_Update/ptr_deref_1106_Merge/merge_req
      -- CP-element group 4: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1106_update_completed_
      -- 
    ca_3247_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1106_load_0_ack_1, ack => sendOutput_CP_3122_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (5) 
      -- CP-element group 5: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1118_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1118_Sample/word_access_start/$exit
      -- CP-element group 5: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1118_Sample/word_access_start/word_0/$exit
      -- CP-element group 5: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1118_Sample/word_access_start/word_0/ra
      -- CP-element group 5: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1118_sample_completed_
      -- 
    ra_3286_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1118_load_0_ack_0, ack => sendOutput_CP_3122_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	0 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1118_Update/ptr_deref_1118_Merge/merge_ack
      -- CP-element group 6: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1118_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1118_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1118_Update/word_access_complete/$exit
      -- CP-element group 6: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1118_Update/word_access_complete/word_0/$exit
      -- CP-element group 6: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1118_Update/ptr_deref_1118_Merge/merge_req
      -- CP-element group 6: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1118_Update/word_access_complete/word_0/ca
      -- CP-element group 6: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1118_Update/ptr_deref_1118_Merge/$entry
      -- CP-element group 6: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/ptr_deref_1118_Update/ptr_deref_1118_Merge/$exit
      -- 
    ca_3297_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1118_load_0_ack_1, ack => sendOutput_CP_3122_elements(6)); -- 
    -- CP-element group 7:  branch  join  transition  place  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	2 
    -- CP-element group 7: 	4 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7: 	9 
    -- CP-element group 7:  members (10) 
      -- CP-element group 7: 	 branch_block_stmt_1083/if_stmt_1136_dead_link/$entry
      -- CP-element group 7: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135/$exit
      -- CP-element group 7: 	 branch_block_stmt_1083/if_stmt_1136_else_link/$entry
      -- CP-element group 7: 	 branch_block_stmt_1083/if_stmt_1136_eval_test/branch_req
      -- CP-element group 7: 	 branch_block_stmt_1083/if_stmt_1136__entry__
      -- CP-element group 7: 	 branch_block_stmt_1083/R_cmp73_1137_place
      -- CP-element group 7: 	 branch_block_stmt_1083/assign_stmt_1091_to_assign_stmt_1135__exit__
      -- CP-element group 7: 	 branch_block_stmt_1083/if_stmt_1136_if_link/$entry
      -- CP-element group 7: 	 branch_block_stmt_1083/if_stmt_1136_eval_test/$entry
      -- CP-element group 7: 	 branch_block_stmt_1083/if_stmt_1136_eval_test/$exit
      -- 
    branch_req_3310_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3310_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3122_elements(7), ack => if_stmt_1136_branch_req_0); -- 
    sendOutput_cp_element_group_7: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "sendOutput_cp_element_group_7"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= sendOutput_CP_3122_elements(2) & sendOutput_CP_3122_elements(4) & sendOutput_CP_3122_elements(6);
      gj_sendOutput_cp_element_group_7 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_3122_elements(7), clk => clk, reset => reset); --
    end block;
    -- CP-element group 8:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	10 
    -- CP-element group 8: 	11 
    -- CP-element group 8:  members (18) 
      -- CP-element group 8: 	 branch_block_stmt_1083/assign_stmt_1148_to_assign_stmt_1177/type_cast_1163_Sample/rr
      -- CP-element group 8: 	 branch_block_stmt_1083/merge_stmt_1142__exit__
      -- CP-element group 8: 	 branch_block_stmt_1083/assign_stmt_1148_to_assign_stmt_1177__entry__
      -- CP-element group 8: 	 branch_block_stmt_1083/assign_stmt_1148_to_assign_stmt_1177/type_cast_1163_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_1083/if_stmt_1136_if_link/$exit
      -- CP-element group 8: 	 branch_block_stmt_1083/assign_stmt_1148_to_assign_stmt_1177/type_cast_1163_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_1083/entry_bbx_xnph
      -- CP-element group 8: 	 branch_block_stmt_1083/assign_stmt_1148_to_assign_stmt_1177/type_cast_1163_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_1083/assign_stmt_1148_to_assign_stmt_1177/type_cast_1163_update_start_
      -- CP-element group 8: 	 branch_block_stmt_1083/assign_stmt_1148_to_assign_stmt_1177/type_cast_1163_Update/cr
      -- CP-element group 8: 	 branch_block_stmt_1083/assign_stmt_1148_to_assign_stmt_1177/$entry
      -- CP-element group 8: 	 branch_block_stmt_1083/if_stmt_1136_if_link/if_choice_transition
      -- CP-element group 8: 	 branch_block_stmt_1083/entry_bbx_xnph_PhiReq/$entry
      -- CP-element group 8: 	 branch_block_stmt_1083/entry_bbx_xnph_PhiReq/$exit
      -- CP-element group 8: 	 branch_block_stmt_1083/merge_stmt_1142_PhiReqMerge
      -- CP-element group 8: 	 branch_block_stmt_1083/merge_stmt_1142_PhiAck/$entry
      -- CP-element group 8: 	 branch_block_stmt_1083/merge_stmt_1142_PhiAck/$exit
      -- CP-element group 8: 	 branch_block_stmt_1083/merge_stmt_1142_PhiAck/dummy
      -- 
    if_choice_transition_3315_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1136_branch_ack_1, ack => sendOutput_CP_3122_elements(8)); -- 
    rr_3332_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3332_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3122_elements(8), ack => type_cast_1163_inst_req_0); -- 
    cr_3337_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3337_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3122_elements(8), ack => type_cast_1163_inst_req_1); -- 
    -- CP-element group 9:  transition  place  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	7 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	66 
    -- CP-element group 9:  members (5) 
      -- CP-element group 9: 	 branch_block_stmt_1083/if_stmt_1136_else_link/$exit
      -- CP-element group 9: 	 branch_block_stmt_1083/entry_forx_xend
      -- CP-element group 9: 	 branch_block_stmt_1083/if_stmt_1136_else_link/else_choice_transition
      -- CP-element group 9: 	 branch_block_stmt_1083/entry_forx_xend_PhiReq/$entry
      -- CP-element group 9: 	 branch_block_stmt_1083/entry_forx_xend_PhiReq/$exit
      -- 
    else_choice_transition_3319_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1136_branch_ack_0, ack => sendOutput_CP_3122_elements(9)); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	8 
    -- CP-element group 10: successors 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_1083/assign_stmt_1148_to_assign_stmt_1177/type_cast_1163_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_1083/assign_stmt_1148_to_assign_stmt_1177/type_cast_1163_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_1083/assign_stmt_1148_to_assign_stmt_1177/type_cast_1163_sample_completed_
      -- 
    ra_3333_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1163_inst_ack_0, ack => sendOutput_CP_3122_elements(10)); -- 
    -- CP-element group 11:  transition  place  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	8 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	60 
    -- CP-element group 11:  members (9) 
      -- CP-element group 11: 	 branch_block_stmt_1083/assign_stmt_1148_to_assign_stmt_1177__exit__
      -- CP-element group 11: 	 branch_block_stmt_1083/bbx_xnph_forx_xbody
      -- CP-element group 11: 	 branch_block_stmt_1083/assign_stmt_1148_to_assign_stmt_1177/type_cast_1163_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_1083/assign_stmt_1148_to_assign_stmt_1177/type_cast_1163_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_1083/assign_stmt_1148_to_assign_stmt_1177/type_cast_1163_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_1083/assign_stmt_1148_to_assign_stmt_1177/$exit
      -- CP-element group 11: 	 branch_block_stmt_1083/bbx_xnph_forx_xbody_PhiReq/$entry
      -- CP-element group 11: 	 branch_block_stmt_1083/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1180/$entry
      -- CP-element group 11: 	 branch_block_stmt_1083/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1180/phi_stmt_1180_sources/$entry
      -- 
    ca_3338_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1163_inst_ack_1, ack => sendOutput_CP_3122_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	65 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	57 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/array_obj_ref_1192_final_index_sum_regn_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/array_obj_ref_1192_final_index_sum_regn_sample_complete
      -- CP-element group 12: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/array_obj_ref_1192_final_index_sum_regn_Sample/ack
      -- 
    ack_3367_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1192_index_offset_ack_0, ack => sendOutput_CP_3122_elements(12)); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	65 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (11) 
      -- CP-element group 13: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/array_obj_ref_1192_final_index_sum_regn_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/array_obj_ref_1192_final_index_sum_regn_Update/ack
      -- CP-element group 13: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/array_obj_ref_1192_base_plus_offset/$exit
      -- CP-element group 13: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/array_obj_ref_1192_base_plus_offset/$entry
      -- CP-element group 13: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/addr_of_1193_request/$entry
      -- CP-element group 13: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/array_obj_ref_1192_base_plus_offset/sum_rename_req
      -- CP-element group 13: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/addr_of_1193_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/array_obj_ref_1192_base_plus_offset/sum_rename_ack
      -- CP-element group 13: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/array_obj_ref_1192_offset_calculated
      -- CP-element group 13: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/array_obj_ref_1192_root_address_calculated
      -- CP-element group 13: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/addr_of_1193_request/req
      -- 
    ack_3372_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1192_index_offset_ack_1, ack => sendOutput_CP_3122_elements(13)); -- 
    req_3381_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3381_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3122_elements(13), ack => addr_of_1193_final_reg_req_0); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/addr_of_1193_request/$exit
      -- CP-element group 14: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/addr_of_1193_request/ack
      -- CP-element group 14: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/addr_of_1193_sample_completed_
      -- 
    ack_3382_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1193_final_reg_ack_0, ack => sendOutput_CP_3122_elements(14)); -- 
    -- CP-element group 15:  join  fork  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	65 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (24) 
      -- CP-element group 15: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/ptr_deref_1197_base_addr_resize/base_resize_ack
      -- CP-element group 15: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/ptr_deref_1197_base_addr_resize/$exit
      -- CP-element group 15: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/ptr_deref_1197_word_addrgen/$exit
      -- CP-element group 15: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/ptr_deref_1197_base_plus_offset/$exit
      -- CP-element group 15: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/ptr_deref_1197_Sample/word_access_start/word_0/rr
      -- CP-element group 15: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/ptr_deref_1197_word_addrgen/$entry
      -- CP-element group 15: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/ptr_deref_1197_base_addr_resize/base_resize_req
      -- CP-element group 15: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/ptr_deref_1197_word_addrgen/root_register_req
      -- CP-element group 15: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/ptr_deref_1197_base_plus_offset/sum_rename_req
      -- CP-element group 15: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/ptr_deref_1197_base_plus_offset/sum_rename_ack
      -- CP-element group 15: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/ptr_deref_1197_base_addr_resize/$entry
      -- CP-element group 15: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/ptr_deref_1197_word_addrgen/root_register_ack
      -- CP-element group 15: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/ptr_deref_1197_base_address_resized
      -- CP-element group 15: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/ptr_deref_1197_base_plus_offset/$entry
      -- CP-element group 15: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/ptr_deref_1197_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/ptr_deref_1197_word_address_calculated
      -- CP-element group 15: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/ptr_deref_1197_root_address_calculated
      -- CP-element group 15: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/ptr_deref_1197_base_address_calculated
      -- CP-element group 15: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/addr_of_1193_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/ptr_deref_1197_Sample/word_access_start/word_0/$entry
      -- CP-element group 15: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/ptr_deref_1197_Sample/word_access_start/$entry
      -- CP-element group 15: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/addr_of_1193_complete/ack
      -- CP-element group 15: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/ptr_deref_1197_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/addr_of_1193_complete/$exit
      -- 
    ack_3387_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1193_final_reg_ack_1, ack => sendOutput_CP_3122_elements(15)); -- 
    rr_3420_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3420_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3122_elements(15), ack => ptr_deref_1197_load_0_req_0); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (5) 
      -- CP-element group 16: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/ptr_deref_1197_Sample/word_access_start/word_0/ra
      -- CP-element group 16: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/ptr_deref_1197_Sample/word_access_start/word_0/$exit
      -- CP-element group 16: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/ptr_deref_1197_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/ptr_deref_1197_Sample/word_access_start/$exit
      -- CP-element group 16: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/ptr_deref_1197_sample_completed_
      -- 
    ra_3421_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1197_load_0_ack_0, ack => sendOutput_CP_3122_elements(16)); -- 
    -- CP-element group 17:  fork  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	65 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17: 	20 
    -- CP-element group 17: 	22 
    -- CP-element group 17: 	24 
    -- CP-element group 17: 	26 
    -- CP-element group 17: 	28 
    -- CP-element group 17: 	30 
    -- CP-element group 17: 	32 
    -- CP-element group 17:  members (33) 
      -- CP-element group 17: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/ptr_deref_1197_Update/ptr_deref_1197_Merge/merge_ack
      -- CP-element group 17: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/ptr_deref_1197_Update/ptr_deref_1197_Merge/merge_req
      -- CP-element group 17: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/ptr_deref_1197_Update/ptr_deref_1197_Merge/$entry
      -- CP-element group 17: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/ptr_deref_1197_Update/ptr_deref_1197_Merge/$exit
      -- CP-element group 17: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1231_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1201_Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/ptr_deref_1197_Update/word_access_complete/$exit
      -- CP-element group 17: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1201_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/ptr_deref_1197_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1231_Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/ptr_deref_1197_Update/word_access_complete/word_0/ca
      -- CP-element group 17: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/ptr_deref_1197_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/ptr_deref_1197_Update/word_access_complete/word_0/$exit
      -- CP-element group 17: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1251_Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1251_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1231_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1271_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1271_Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1261_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1261_Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1241_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1221_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1261_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1241_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1241_Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1221_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1211_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1271_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1251_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1211_Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1211_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1221_Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1201_sample_start_
      -- 
    ca_3432_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1197_load_0_ack_1, ack => sendOutput_CP_3122_elements(17)); -- 
    rr_3445_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3445_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3122_elements(17), ack => type_cast_1201_inst_req_0); -- 
    rr_3459_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3459_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3122_elements(17), ack => type_cast_1211_inst_req_0); -- 
    rr_3473_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3473_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3122_elements(17), ack => type_cast_1221_inst_req_0); -- 
    rr_3487_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3487_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3122_elements(17), ack => type_cast_1231_inst_req_0); -- 
    rr_3501_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3501_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3122_elements(17), ack => type_cast_1241_inst_req_0); -- 
    rr_3515_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3515_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3122_elements(17), ack => type_cast_1251_inst_req_0); -- 
    rr_3529_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3529_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3122_elements(17), ack => type_cast_1261_inst_req_0); -- 
    rr_3543_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3543_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3122_elements(17), ack => type_cast_1271_inst_req_0); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1201_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1201_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1201_Sample/ra
      -- 
    ra_3446_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1201_inst_ack_0, ack => sendOutput_CP_3122_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	65 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	54 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1201_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1201_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1201_Update/ca
      -- 
    ca_3451_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1201_inst_ack_1, ack => sendOutput_CP_3122_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	17 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1211_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1211_Sample/ra
      -- CP-element group 20: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1211_Sample/$exit
      -- 
    ra_3460_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1211_inst_ack_0, ack => sendOutput_CP_3122_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	65 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	51 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1211_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1211_Update/ca
      -- CP-element group 21: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1211_Update/$exit
      -- 
    ca_3465_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1211_inst_ack_1, ack => sendOutput_CP_3122_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	17 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1221_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1221_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1221_Sample/ra
      -- 
    ra_3474_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1221_inst_ack_0, ack => sendOutput_CP_3122_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	65 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	48 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1221_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1221_Update/ca
      -- CP-element group 23: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1221_update_completed_
      -- 
    ca_3479_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1221_inst_ack_1, ack => sendOutput_CP_3122_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	17 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1231_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1231_Sample/ra
      -- CP-element group 24: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1231_sample_completed_
      -- 
    ra_3488_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1231_inst_ack_0, ack => sendOutput_CP_3122_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	65 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	45 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1231_Update/ca
      -- CP-element group 25: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1231_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1231_Update/$exit
      -- 
    ca_3493_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1231_inst_ack_1, ack => sendOutput_CP_3122_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	17 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1241_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1241_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1241_Sample/ra
      -- 
    ra_3502_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1241_inst_ack_0, ack => sendOutput_CP_3122_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	65 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	42 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1241_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1241_Update/ca
      -- CP-element group 27: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1241_Update/$exit
      -- 
    ca_3507_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1241_inst_ack_1, ack => sendOutput_CP_3122_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	17 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1251_Sample/ra
      -- CP-element group 28: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1251_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1251_sample_completed_
      -- 
    ra_3516_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1251_inst_ack_0, ack => sendOutput_CP_3122_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	65 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	39 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1251_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1251_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1251_Update/$exit
      -- 
    ca_3521_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1251_inst_ack_1, ack => sendOutput_CP_3122_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	17 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1261_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1261_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1261_Sample/ra
      -- 
    ra_3530_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1261_inst_ack_0, ack => sendOutput_CP_3122_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	65 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	36 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1261_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1261_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1261_Update/$exit
      -- 
    ca_3535_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1261_inst_ack_1, ack => sendOutput_CP_3122_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	17 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1271_Sample/ra
      -- CP-element group 32: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1271_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1271_sample_completed_
      -- 
    ra_3544_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1271_inst_ack_0, ack => sendOutput_CP_3122_elements(32)); -- 
    -- CP-element group 33:  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	65 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (6) 
      -- CP-element group 33: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1271_Update/ca
      -- CP-element group 33: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1271_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1271_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1273_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1273_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1273_Sample/req
      -- 
    ca_3549_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1271_inst_ack_1, ack => sendOutput_CP_3122_elements(33)); -- 
    req_3557_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3557_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3122_elements(33), ack => WPIPE_ConvTranspose_output_pipe_1273_inst_req_0); -- 
    -- CP-element group 34:  transition  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34:  members (6) 
      -- CP-element group 34: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1273_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1273_Update/req
      -- CP-element group 34: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1273_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1273_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1273_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1273_Sample/ack
      -- 
    ack_3558_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1273_inst_ack_0, ack => sendOutput_CP_3122_elements(34)); -- 
    req_3562_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3562_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3122_elements(34), ack => WPIPE_ConvTranspose_output_pipe_1273_inst_req_1); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1273_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1273_Update/ack
      -- CP-element group 35: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1273_update_completed_
      -- 
    ack_3563_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1273_inst_ack_1, ack => sendOutput_CP_3122_elements(35)); -- 
    -- CP-element group 36:  join  transition  output  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	31 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	37 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1276_Sample/$entry
      -- CP-element group 36: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1276_Sample/req
      -- CP-element group 36: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1276_sample_start_
      -- 
    req_3571_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3571_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3122_elements(36), ack => WPIPE_ConvTranspose_output_pipe_1276_inst_req_0); -- 
    sendOutput_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_3122_elements(31) & sendOutput_CP_3122_elements(35);
      gj_sendOutput_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_3122_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	36 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (6) 
      -- CP-element group 37: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1276_Update/req
      -- CP-element group 37: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1276_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1276_Sample/ack
      -- CP-element group 37: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1276_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1276_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1276_update_start_
      -- 
    ack_3572_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1276_inst_ack_0, ack => sendOutput_CP_3122_elements(37)); -- 
    req_3576_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3576_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3122_elements(37), ack => WPIPE_ConvTranspose_output_pipe_1276_inst_req_1); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1276_Update/ack
      -- CP-element group 38: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1276_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1276_update_completed_
      -- 
    ack_3577_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1276_inst_ack_1, ack => sendOutput_CP_3122_elements(38)); -- 
    -- CP-element group 39:  join  transition  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	29 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1279_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1279_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1279_Sample/req
      -- 
    req_3585_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3585_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3122_elements(39), ack => WPIPE_ConvTranspose_output_pipe_1279_inst_req_0); -- 
    sendOutput_cp_element_group_39: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_39"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_3122_elements(29) & sendOutput_CP_3122_elements(38);
      gj_sendOutput_cp_element_group_39 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_3122_elements(39), clk => clk, reset => reset); --
    end block;
    -- CP-element group 40:  transition  input  output  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (6) 
      -- CP-element group 40: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1279_Update/$entry
      -- CP-element group 40: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1279_Update/req
      -- CP-element group 40: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1279_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1279_update_start_
      -- CP-element group 40: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1279_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1279_Sample/ack
      -- 
    ack_3586_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1279_inst_ack_0, ack => sendOutput_CP_3122_elements(40)); -- 
    req_3590_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3590_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3122_elements(40), ack => WPIPE_ConvTranspose_output_pipe_1279_inst_req_1); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1279_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1279_Update/ack
      -- CP-element group 41: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1279_update_completed_
      -- 
    ack_3591_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1279_inst_ack_1, ack => sendOutput_CP_3122_elements(41)); -- 
    -- CP-element group 42:  join  transition  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	27 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1282_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1282_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1282_Sample/req
      -- 
    req_3599_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3599_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3122_elements(42), ack => WPIPE_ConvTranspose_output_pipe_1282_inst_req_0); -- 
    sendOutput_cp_element_group_42: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_42"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_3122_elements(27) & sendOutput_CP_3122_elements(41);
      gj_sendOutput_cp_element_group_42 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_3122_elements(42), clk => clk, reset => reset); --
    end block;
    -- CP-element group 43:  transition  input  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (6) 
      -- CP-element group 43: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1282_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1282_update_start_
      -- CP-element group 43: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1282_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1282_Sample/ack
      -- CP-element group 43: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1282_Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1282_Update/req
      -- 
    ack_3600_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1282_inst_ack_0, ack => sendOutput_CP_3122_elements(43)); -- 
    req_3604_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3604_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3122_elements(43), ack => WPIPE_ConvTranspose_output_pipe_1282_inst_req_1); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1282_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1282_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1282_Update/ack
      -- 
    ack_3605_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1282_inst_ack_1, ack => sendOutput_CP_3122_elements(44)); -- 
    -- CP-element group 45:  join  transition  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	25 
    -- CP-element group 45: 	44 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1285_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1285_Sample/$entry
      -- CP-element group 45: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1285_Sample/req
      -- 
    req_3613_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3613_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3122_elements(45), ack => WPIPE_ConvTranspose_output_pipe_1285_inst_req_0); -- 
    sendOutput_cp_element_group_45: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_45"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_3122_elements(25) & sendOutput_CP_3122_elements(44);
      gj_sendOutput_cp_element_group_45 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_3122_elements(45), clk => clk, reset => reset); --
    end block;
    -- CP-element group 46:  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (6) 
      -- CP-element group 46: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1285_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1285_update_start_
      -- CP-element group 46: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1285_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1285_Sample/ack
      -- CP-element group 46: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1285_Update/$entry
      -- CP-element group 46: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1285_Update/req
      -- 
    ack_3614_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1285_inst_ack_0, ack => sendOutput_CP_3122_elements(46)); -- 
    req_3618_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3618_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3122_elements(46), ack => WPIPE_ConvTranspose_output_pipe_1285_inst_req_1); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1285_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1285_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1285_Update/ack
      -- 
    ack_3619_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1285_inst_ack_1, ack => sendOutput_CP_3122_elements(47)); -- 
    -- CP-element group 48:  join  transition  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	23 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1288_sample_start_
      -- CP-element group 48: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1288_Sample/$entry
      -- CP-element group 48: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1288_Sample/req
      -- 
    req_3627_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3627_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3122_elements(48), ack => WPIPE_ConvTranspose_output_pipe_1288_inst_req_0); -- 
    sendOutput_cp_element_group_48: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_48"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_3122_elements(23) & sendOutput_CP_3122_elements(47);
      gj_sendOutput_cp_element_group_48 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_3122_elements(48), clk => clk, reset => reset); --
    end block;
    -- CP-element group 49:  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (6) 
      -- CP-element group 49: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1288_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1288_update_start_
      -- CP-element group 49: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1288_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1288_Sample/ack
      -- CP-element group 49: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1288_Update/$entry
      -- CP-element group 49: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1288_Update/req
      -- 
    ack_3628_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1288_inst_ack_0, ack => sendOutput_CP_3122_elements(49)); -- 
    req_3632_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3632_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3122_elements(49), ack => WPIPE_ConvTranspose_output_pipe_1288_inst_req_1); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1288_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1288_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1288_Update/ack
      -- 
    ack_3633_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1288_inst_ack_1, ack => sendOutput_CP_3122_elements(50)); -- 
    -- CP-element group 51:  join  transition  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	21 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1291_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1291_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1291_Sample/req
      -- 
    req_3641_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3641_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3122_elements(51), ack => WPIPE_ConvTranspose_output_pipe_1291_inst_req_0); -- 
    sendOutput_cp_element_group_51: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_51"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_3122_elements(21) & sendOutput_CP_3122_elements(50);
      gj_sendOutput_cp_element_group_51 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_3122_elements(51), clk => clk, reset => reset); --
    end block;
    -- CP-element group 52:  transition  input  output  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	53 
    -- CP-element group 52:  members (6) 
      -- CP-element group 52: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1291_sample_completed_
      -- CP-element group 52: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1291_update_start_
      -- CP-element group 52: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1291_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1291_Sample/ack
      -- CP-element group 52: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1291_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1291_Update/req
      -- 
    ack_3642_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1291_inst_ack_0, ack => sendOutput_CP_3122_elements(52)); -- 
    req_3646_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3646_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3122_elements(52), ack => WPIPE_ConvTranspose_output_pipe_1291_inst_req_1); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	52 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1291_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1291_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1291_Update/ack
      -- 
    ack_3647_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1291_inst_ack_1, ack => sendOutput_CP_3122_elements(53)); -- 
    -- CP-element group 54:  join  transition  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	19 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1294_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1294_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1294_Sample/req
      -- 
    req_3655_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3655_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3122_elements(54), ack => WPIPE_ConvTranspose_output_pipe_1294_inst_req_0); -- 
    sendOutput_cp_element_group_54: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_54"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_3122_elements(19) & sendOutput_CP_3122_elements(53);
      gj_sendOutput_cp_element_group_54 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_3122_elements(54), clk => clk, reset => reset); --
    end block;
    -- CP-element group 55:  transition  input  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (6) 
      -- CP-element group 55: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1294_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1294_update_start_
      -- CP-element group 55: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1294_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1294_Sample/ack
      -- CP-element group 55: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1294_Update/$entry
      -- CP-element group 55: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1294_Update/req
      -- 
    ack_3656_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1294_inst_ack_0, ack => sendOutput_CP_3122_elements(55)); -- 
    req_3660_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3660_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3122_elements(55), ack => WPIPE_ConvTranspose_output_pipe_1294_inst_req_1); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1294_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1294_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/WPIPE_ConvTranspose_output_pipe_1294_Update/ack
      -- 
    ack_3661_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1294_inst_ack_1, ack => sendOutput_CP_3122_elements(56)); -- 
    -- CP-element group 57:  branch  join  transition  place  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	12 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57: 	59 
    -- CP-element group 57:  members (10) 
      -- CP-element group 57: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307__exit__
      -- CP-element group 57: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/$exit
      -- CP-element group 57: 	 branch_block_stmt_1083/if_stmt_1308__entry__
      -- CP-element group 57: 	 branch_block_stmt_1083/if_stmt_1308_dead_link/$entry
      -- CP-element group 57: 	 branch_block_stmt_1083/if_stmt_1308_eval_test/$entry
      -- CP-element group 57: 	 branch_block_stmt_1083/if_stmt_1308_eval_test/$exit
      -- CP-element group 57: 	 branch_block_stmt_1083/if_stmt_1308_eval_test/branch_req
      -- CP-element group 57: 	 branch_block_stmt_1083/R_exitcond1_1309_place
      -- CP-element group 57: 	 branch_block_stmt_1083/if_stmt_1308_if_link/$entry
      -- CP-element group 57: 	 branch_block_stmt_1083/if_stmt_1308_else_link/$entry
      -- 
    branch_req_3669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3122_elements(57), ack => if_stmt_1308_branch_req_0); -- 
    sendOutput_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_3122_elements(12) & sendOutput_CP_3122_elements(56);
      gj_sendOutput_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_3122_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  merge  transition  place  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	66 
    -- CP-element group 58:  members (13) 
      -- CP-element group 58: 	 branch_block_stmt_1083/merge_stmt_1314__exit__
      -- CP-element group 58: 	 branch_block_stmt_1083/forx_xendx_xloopexit_forx_xend
      -- CP-element group 58: 	 branch_block_stmt_1083/if_stmt_1308_if_link/$exit
      -- CP-element group 58: 	 branch_block_stmt_1083/if_stmt_1308_if_link/if_choice_transition
      -- CP-element group 58: 	 branch_block_stmt_1083/forx_xbody_forx_xendx_xloopexit
      -- CP-element group 58: 	 branch_block_stmt_1083/forx_xbody_forx_xendx_xloopexit_PhiReq/$entry
      -- CP-element group 58: 	 branch_block_stmt_1083/forx_xbody_forx_xendx_xloopexit_PhiReq/$exit
      -- CP-element group 58: 	 branch_block_stmt_1083/merge_stmt_1314_PhiReqMerge
      -- CP-element group 58: 	 branch_block_stmt_1083/merge_stmt_1314_PhiAck/$entry
      -- CP-element group 58: 	 branch_block_stmt_1083/merge_stmt_1314_PhiAck/$exit
      -- CP-element group 58: 	 branch_block_stmt_1083/merge_stmt_1314_PhiAck/dummy
      -- CP-element group 58: 	 branch_block_stmt_1083/forx_xendx_xloopexit_forx_xend_PhiReq/$entry
      -- CP-element group 58: 	 branch_block_stmt_1083/forx_xendx_xloopexit_forx_xend_PhiReq/$exit
      -- 
    if_choice_transition_3674_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1308_branch_ack_1, ack => sendOutput_CP_3122_elements(58)); -- 
    -- CP-element group 59:  fork  transition  place  input  output  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	57 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	61 
    -- CP-element group 59: 	62 
    -- CP-element group 59:  members (12) 
      -- CP-element group 59: 	 branch_block_stmt_1083/if_stmt_1308_else_link/$exit
      -- CP-element group 59: 	 branch_block_stmt_1083/if_stmt_1308_else_link/else_choice_transition
      -- CP-element group 59: 	 branch_block_stmt_1083/forx_xbody_forx_xbody
      -- CP-element group 59: 	 branch_block_stmt_1083/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 59: 	 branch_block_stmt_1083/forx_xbody_forx_xbody_PhiReq/phi_stmt_1180/$entry
      -- CP-element group 59: 	 branch_block_stmt_1083/forx_xbody_forx_xbody_PhiReq/phi_stmt_1180/phi_stmt_1180_sources/$entry
      -- CP-element group 59: 	 branch_block_stmt_1083/forx_xbody_forx_xbody_PhiReq/phi_stmt_1180/phi_stmt_1180_sources/type_cast_1186/$entry
      -- CP-element group 59: 	 branch_block_stmt_1083/forx_xbody_forx_xbody_PhiReq/phi_stmt_1180/phi_stmt_1180_sources/type_cast_1186/SplitProtocol/$entry
      -- CP-element group 59: 	 branch_block_stmt_1083/forx_xbody_forx_xbody_PhiReq/phi_stmt_1180/phi_stmt_1180_sources/type_cast_1186/SplitProtocol/Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_1083/forx_xbody_forx_xbody_PhiReq/phi_stmt_1180/phi_stmt_1180_sources/type_cast_1186/SplitProtocol/Sample/rr
      -- CP-element group 59: 	 branch_block_stmt_1083/forx_xbody_forx_xbody_PhiReq/phi_stmt_1180/phi_stmt_1180_sources/type_cast_1186/SplitProtocol/Update/$entry
      -- CP-element group 59: 	 branch_block_stmt_1083/forx_xbody_forx_xbody_PhiReq/phi_stmt_1180/phi_stmt_1180_sources/type_cast_1186/SplitProtocol/Update/cr
      -- 
    else_choice_transition_3678_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1308_branch_ack_0, ack => sendOutput_CP_3122_elements(59)); -- 
    rr_3722_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3722_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3122_elements(59), ack => type_cast_1186_inst_req_0); -- 
    cr_3727_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3727_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3122_elements(59), ack => type_cast_1186_inst_req_1); -- 
    -- CP-element group 60:  transition  output  delay-element  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	11 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	64 
    -- CP-element group 60:  members (5) 
      -- CP-element group 60: 	 branch_block_stmt_1083/bbx_xnph_forx_xbody_PhiReq/$exit
      -- CP-element group 60: 	 branch_block_stmt_1083/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1180/$exit
      -- CP-element group 60: 	 branch_block_stmt_1083/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1180/phi_stmt_1180_sources/$exit
      -- CP-element group 60: 	 branch_block_stmt_1083/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1180/phi_stmt_1180_sources/type_cast_1184_konst_delay_trans
      -- CP-element group 60: 	 branch_block_stmt_1083/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1180/phi_stmt_1180_req
      -- 
    phi_stmt_1180_req_3703_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1180_req_3703_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3122_elements(60), ack => phi_stmt_1180_req_0); -- 
    -- Element group sendOutput_CP_3122_elements(60) is a control-delay.
    cp_element_60_delay: control_delay_element  generic map(name => " 60_delay", delay_value => 1)  port map(req => sendOutput_CP_3122_elements(11), ack => sendOutput_CP_3122_elements(60), clk => clk, reset =>reset);
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	59 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	63 
    -- CP-element group 61:  members (2) 
      -- CP-element group 61: 	 branch_block_stmt_1083/forx_xbody_forx_xbody_PhiReq/phi_stmt_1180/phi_stmt_1180_sources/type_cast_1186/SplitProtocol/Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_1083/forx_xbody_forx_xbody_PhiReq/phi_stmt_1180/phi_stmt_1180_sources/type_cast_1186/SplitProtocol/Sample/ra
      -- 
    ra_3723_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1186_inst_ack_0, ack => sendOutput_CP_3122_elements(61)); -- 
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	59 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (2) 
      -- CP-element group 62: 	 branch_block_stmt_1083/forx_xbody_forx_xbody_PhiReq/phi_stmt_1180/phi_stmt_1180_sources/type_cast_1186/SplitProtocol/Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_1083/forx_xbody_forx_xbody_PhiReq/phi_stmt_1180/phi_stmt_1180_sources/type_cast_1186/SplitProtocol/Update/ca
      -- 
    ca_3728_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1186_inst_ack_1, ack => sendOutput_CP_3122_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	61 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (6) 
      -- CP-element group 63: 	 branch_block_stmt_1083/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 63: 	 branch_block_stmt_1083/forx_xbody_forx_xbody_PhiReq/phi_stmt_1180/$exit
      -- CP-element group 63: 	 branch_block_stmt_1083/forx_xbody_forx_xbody_PhiReq/phi_stmt_1180/phi_stmt_1180_sources/$exit
      -- CP-element group 63: 	 branch_block_stmt_1083/forx_xbody_forx_xbody_PhiReq/phi_stmt_1180/phi_stmt_1180_sources/type_cast_1186/$exit
      -- CP-element group 63: 	 branch_block_stmt_1083/forx_xbody_forx_xbody_PhiReq/phi_stmt_1180/phi_stmt_1180_sources/type_cast_1186/SplitProtocol/$exit
      -- CP-element group 63: 	 branch_block_stmt_1083/forx_xbody_forx_xbody_PhiReq/phi_stmt_1180/phi_stmt_1180_req
      -- 
    phi_stmt_1180_req_3729_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1180_req_3729_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3122_elements(63), ack => phi_stmt_1180_req_1); -- 
    sendOutput_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_3122_elements(61) & sendOutput_CP_3122_elements(62);
      gj_sendOutput_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_3122_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  merge  transition  place  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	60 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64:  members (2) 
      -- CP-element group 64: 	 branch_block_stmt_1083/merge_stmt_1179_PhiReqMerge
      -- CP-element group 64: 	 branch_block_stmt_1083/merge_stmt_1179_PhiAck/$entry
      -- 
    sendOutput_CP_3122_elements(64) <= OrReduce(sendOutput_CP_3122_elements(60) & sendOutput_CP_3122_elements(63));
    -- CP-element group 65:  fork  transition  place  input  output  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	12 
    -- CP-element group 65: 	13 
    -- CP-element group 65: 	15 
    -- CP-element group 65: 	17 
    -- CP-element group 65: 	19 
    -- CP-element group 65: 	21 
    -- CP-element group 65: 	23 
    -- CP-element group 65: 	25 
    -- CP-element group 65: 	27 
    -- CP-element group 65: 	29 
    -- CP-element group 65: 	31 
    -- CP-element group 65: 	33 
    -- CP-element group 65:  members (53) 
      -- CP-element group 65: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/array_obj_ref_1192_index_resize_1/index_resize_ack
      -- CP-element group 65: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/array_obj_ref_1192_index_scale_1/$exit
      -- CP-element group 65: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/array_obj_ref_1192_final_index_sum_regn_Update/req
      -- CP-element group 65: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/array_obj_ref_1192_index_scale_1/$entry
      -- CP-element group 65: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1201_Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/array_obj_ref_1192_index_resize_1/$exit
      -- CP-element group 65: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/ptr_deref_1197_Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307__entry__
      -- CP-element group 65: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/array_obj_ref_1192_index_scale_1/scale_rename_req
      -- CP-element group 65: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/ptr_deref_1197_Update/word_access_complete/$entry
      -- CP-element group 65: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/array_obj_ref_1192_index_resize_1/$entry
      -- CP-element group 65: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1201_Update/cr
      -- CP-element group 65: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/array_obj_ref_1192_final_index_sum_regn_Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1211_update_start_
      -- CP-element group 65: 	 branch_block_stmt_1083/merge_stmt_1179__exit__
      -- CP-element group 65: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/array_obj_ref_1192_index_resized_1
      -- CP-element group 65: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/array_obj_ref_1192_index_scaled_1
      -- CP-element group 65: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/array_obj_ref_1192_index_resize_1/index_resize_req
      -- CP-element group 65: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1231_Update/cr
      -- CP-element group 65: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1271_Update/cr
      -- CP-element group 65: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1221_Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/array_obj_ref_1192_index_computed_1
      -- CP-element group 65: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/array_obj_ref_1192_index_scale_1/scale_rename_ack
      -- CP-element group 65: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1211_Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1221_Update/cr
      -- CP-element group 65: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1271_Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1221_update_start_
      -- CP-element group 65: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/ptr_deref_1197_Update/word_access_complete/word_0/$entry
      -- CP-element group 65: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/ptr_deref_1197_update_start_
      -- CP-element group 65: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1261_update_start_
      -- CP-element group 65: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1241_update_start_
      -- CP-element group 65: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/$entry
      -- CP-element group 65: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1261_Update/cr
      -- CP-element group 65: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1251_update_start_
      -- CP-element group 65: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/array_obj_ref_1192_final_index_sum_regn_update_start
      -- CP-element group 65: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/addr_of_1193_complete/$entry
      -- CP-element group 65: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/array_obj_ref_1192_final_index_sum_regn_Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1241_Update/cr
      -- CP-element group 65: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1231_update_start_
      -- CP-element group 65: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/array_obj_ref_1192_final_index_sum_regn_Sample/req
      -- CP-element group 65: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1241_Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1251_Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1251_Update/cr
      -- CP-element group 65: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/addr_of_1193_update_start_
      -- CP-element group 65: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1271_update_start_
      -- CP-element group 65: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1231_Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/addr_of_1193_complete/req
      -- CP-element group 65: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1261_Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1211_Update/cr
      -- CP-element group 65: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/ptr_deref_1197_Update/word_access_complete/word_0/cr
      -- CP-element group 65: 	 branch_block_stmt_1083/assign_stmt_1194_to_assign_stmt_1307/type_cast_1201_update_start_
      -- CP-element group 65: 	 branch_block_stmt_1083/merge_stmt_1179_PhiAck/$exit
      -- CP-element group 65: 	 branch_block_stmt_1083/merge_stmt_1179_PhiAck/phi_stmt_1180_ack
      -- 
    phi_stmt_1180_ack_3734_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1180_ack_0, ack => sendOutput_CP_3122_elements(65)); -- 
    req_3371_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3371_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3122_elements(65), ack => array_obj_ref_1192_index_offset_req_1); -- 
    cr_3450_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3450_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3122_elements(65), ack => type_cast_1201_inst_req_1); -- 
    cr_3492_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3492_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3122_elements(65), ack => type_cast_1231_inst_req_1); -- 
    cr_3548_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3548_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3122_elements(65), ack => type_cast_1271_inst_req_1); -- 
    cr_3478_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3478_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3122_elements(65), ack => type_cast_1221_inst_req_1); -- 
    cr_3534_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3534_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3122_elements(65), ack => type_cast_1261_inst_req_1); -- 
    cr_3506_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3506_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3122_elements(65), ack => type_cast_1241_inst_req_1); -- 
    req_3366_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3366_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3122_elements(65), ack => array_obj_ref_1192_index_offset_req_0); -- 
    cr_3520_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3520_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3122_elements(65), ack => type_cast_1251_inst_req_1); -- 
    req_3386_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3386_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3122_elements(65), ack => addr_of_1193_final_reg_req_1); -- 
    cr_3464_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3464_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3122_elements(65), ack => type_cast_1211_inst_req_1); -- 
    cr_3431_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3431_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3122_elements(65), ack => ptr_deref_1197_load_0_req_1); -- 
    -- CP-element group 66:  merge  transition  place  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	9 
    -- CP-element group 66: 	58 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (16) 
      -- CP-element group 66: 	 branch_block_stmt_1083/return__
      -- CP-element group 66: 	 branch_block_stmt_1083/merge_stmt_1316__exit__
      -- CP-element group 66: 	 branch_block_stmt_1083/merge_stmt_1318__exit__
      -- CP-element group 66: 	 branch_block_stmt_1083/branch_block_stmt_1083__exit__
      -- CP-element group 66: 	 branch_block_stmt_1083/$exit
      -- CP-element group 66: 	 $exit
      -- CP-element group 66: 	 branch_block_stmt_1083/merge_stmt_1316_PhiReqMerge
      -- CP-element group 66: 	 branch_block_stmt_1083/merge_stmt_1316_PhiAck/$entry
      -- CP-element group 66: 	 branch_block_stmt_1083/merge_stmt_1316_PhiAck/$exit
      -- CP-element group 66: 	 branch_block_stmt_1083/merge_stmt_1316_PhiAck/dummy
      -- CP-element group 66: 	 branch_block_stmt_1083/return___PhiReq/$entry
      -- CP-element group 66: 	 branch_block_stmt_1083/return___PhiReq/$exit
      -- CP-element group 66: 	 branch_block_stmt_1083/merge_stmt_1318_PhiReqMerge
      -- CP-element group 66: 	 branch_block_stmt_1083/merge_stmt_1318_PhiAck/$entry
      -- CP-element group 66: 	 branch_block_stmt_1083/merge_stmt_1318_PhiAck/$exit
      -- CP-element group 66: 	 branch_block_stmt_1083/merge_stmt_1318_PhiAck/dummy
      -- 
    sendOutput_CP_3122_elements(66) <= OrReduce(sendOutput_CP_3122_elements(9) & sendOutput_CP_3122_elements(58));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_indvar_1191_resized : std_logic_vector(13 downto 0);
    signal R_indvar_1191_scaled : std_logic_vector(13 downto 0);
    signal array_obj_ref_1192_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1192_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1192_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1192_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1192_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1192_root_address : std_logic_vector(13 downto 0);
    signal arrayidx_1194 : std_logic_vector(31 downto 0);
    signal cmp73_1135 : std_logic_vector(0 downto 0);
    signal conv17_1212 : std_logic_vector(7 downto 0);
    signal conv23_1222 : std_logic_vector(7 downto 0);
    signal conv29_1232 : std_logic_vector(7 downto 0);
    signal conv35_1242 : std_logic_vector(7 downto 0);
    signal conv41_1252 : std_logic_vector(7 downto 0);
    signal conv47_1262 : std_logic_vector(7 downto 0);
    signal conv53_1272 : std_logic_vector(7 downto 0);
    signal conv_1202 : std_logic_vector(7 downto 0);
    signal exitcond1_1307 : std_logic_vector(0 downto 0);
    signal iNsTr_0_1091 : std_logic_vector(31 downto 0);
    signal iNsTr_1_1103 : std_logic_vector(31 downto 0);
    signal iNsTr_2_1115 : std_logic_vector(31 downto 0);
    signal iNsTr_4_1164 : std_logic_vector(63 downto 0);
    signal indvar_1180 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_1302 : std_logic_vector(63 downto 0);
    signal mul3_1129 : std_logic_vector(31 downto 0);
    signal mul_1124 : std_logic_vector(31 downto 0);
    signal ptr_deref_1094_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1094_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1094_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1094_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1094_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1106_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1106_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1106_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1106_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1106_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1118_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1118_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1118_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1118_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1118_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1197_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1197_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1197_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1197_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1197_word_offset_0 : std_logic_vector(13 downto 0);
    signal shr14_1208 : std_logic_vector(63 downto 0);
    signal shr20_1218 : std_logic_vector(63 downto 0);
    signal shr26_1228 : std_logic_vector(63 downto 0);
    signal shr32_1238 : std_logic_vector(63 downto 0);
    signal shr38_1248 : std_logic_vector(63 downto 0);
    signal shr44_1258 : std_logic_vector(63 downto 0);
    signal shr50_1268 : std_logic_vector(63 downto 0);
    signal tmp1_1107 : std_logic_vector(31 downto 0);
    signal tmp2_1119 : std_logic_vector(31 downto 0);
    signal tmp77_1148 : std_logic_vector(31 downto 0);
    signal tmp77x_xop_1160 : std_logic_vector(31 downto 0);
    signal tmp78_1154 : std_logic_vector(0 downto 0);
    signal tmp81_1177 : std_logic_vector(63 downto 0);
    signal tmp9_1198 : std_logic_vector(63 downto 0);
    signal tmp_1095 : std_logic_vector(31 downto 0);
    signal type_cast_1133_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1146_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1152_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1158_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1168_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1175_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1184_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1186_wire : std_logic_vector(63 downto 0);
    signal type_cast_1206_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1216_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1226_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1236_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1246_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1256_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1266_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1300_wire_constant : std_logic_vector(63 downto 0);
    signal xx_xop_1170 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    array_obj_ref_1192_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1192_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1192_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1192_resized_base_address <= "00000000000000";
    iNsTr_0_1091 <= "00000000000000000000000000000011";
    iNsTr_1_1103 <= "00000000000000000000000000000100";
    iNsTr_2_1115 <= "00000000000000000000000000000101";
    ptr_deref_1094_word_offset_0 <= "0000000";
    ptr_deref_1106_word_offset_0 <= "0000000";
    ptr_deref_1118_word_offset_0 <= "0000000";
    ptr_deref_1197_word_offset_0 <= "00000000000000";
    type_cast_1133_wire_constant <= "00000000000000000000000000000111";
    type_cast_1146_wire_constant <= "00000000000000000000000000000011";
    type_cast_1152_wire_constant <= "00000000000000000000000000000001";
    type_cast_1158_wire_constant <= "11111111111111111111111111111111";
    type_cast_1168_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1175_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1184_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1206_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1216_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1226_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1236_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1246_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1256_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1266_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1300_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    phi_stmt_1180: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1184_wire_constant & type_cast_1186_wire;
      req <= phi_stmt_1180_req_0 & phi_stmt_1180_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1180",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1180_ack_0,
          idata => idata,
          odata => indvar_1180,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1180
    -- flow-through select operator MUX_1176_inst
    tmp81_1177 <= xx_xop_1170 when (tmp78_1154(0) /=  '0') else type_cast_1175_wire_constant;
    addr_of_1193_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1193_final_reg_req_0;
      addr_of_1193_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1193_final_reg_req_1;
      addr_of_1193_final_reg_ack_1<= rack(0);
      addr_of_1193_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1193_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1192_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_1194,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1163_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1163_inst_req_0;
      type_cast_1163_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1163_inst_req_1;
      type_cast_1163_inst_ack_1<= rack(0);
      type_cast_1163_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1163_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp77x_xop_1160,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_4_1164,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1186_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1186_inst_req_0;
      type_cast_1186_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1186_inst_req_1;
      type_cast_1186_inst_ack_1<= rack(0);
      type_cast_1186_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1186_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1302,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1186_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1201_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1201_inst_req_0;
      type_cast_1201_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1201_inst_req_1;
      type_cast_1201_inst_ack_1<= rack(0);
      type_cast_1201_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1201_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp9_1198,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_1202,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1211_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1211_inst_req_0;
      type_cast_1211_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1211_inst_req_1;
      type_cast_1211_inst_ack_1<= rack(0);
      type_cast_1211_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1211_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr14_1208,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_1212,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1221_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1221_inst_req_0;
      type_cast_1221_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1221_inst_req_1;
      type_cast_1221_inst_ack_1<= rack(0);
      type_cast_1221_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1221_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr20_1218,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv23_1222,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1231_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1231_inst_req_0;
      type_cast_1231_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1231_inst_req_1;
      type_cast_1231_inst_ack_1<= rack(0);
      type_cast_1231_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1231_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr26_1228,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv29_1232,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1241_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1241_inst_req_0;
      type_cast_1241_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1241_inst_req_1;
      type_cast_1241_inst_ack_1<= rack(0);
      type_cast_1241_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1241_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr32_1238,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv35_1242,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1251_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1251_inst_req_0;
      type_cast_1251_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1251_inst_req_1;
      type_cast_1251_inst_ack_1<= rack(0);
      type_cast_1251_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1251_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr38_1248,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv41_1252,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1261_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1261_inst_req_0;
      type_cast_1261_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1261_inst_req_1;
      type_cast_1261_inst_ack_1<= rack(0);
      type_cast_1261_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1261_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr44_1258,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv47_1262,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1271_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1271_inst_req_0;
      type_cast_1271_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1271_inst_req_1;
      type_cast_1271_inst_ack_1<= rack(0);
      type_cast_1271_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1271_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr50_1268,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv53_1272,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1192_index_1_rename
    process(R_indvar_1191_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_1191_resized;
      ov(13 downto 0) := iv;
      R_indvar_1191_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1192_index_1_resize
    process(indvar_1180) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_1180;
      ov := iv(13 downto 0);
      R_indvar_1191_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1192_root_address_inst
    process(array_obj_ref_1192_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1192_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1192_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1094_addr_0
    process(ptr_deref_1094_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1094_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1094_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1094_base_resize
    process(iNsTr_0_1091) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_0_1091;
      ov := iv(6 downto 0);
      ptr_deref_1094_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1094_gather_scatter
    process(ptr_deref_1094_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1094_data_0;
      ov(31 downto 0) := iv;
      tmp_1095 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1094_root_address_inst
    process(ptr_deref_1094_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1094_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1094_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1106_addr_0
    process(ptr_deref_1106_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1106_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1106_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1106_base_resize
    process(iNsTr_1_1103) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_1_1103;
      ov := iv(6 downto 0);
      ptr_deref_1106_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1106_gather_scatter
    process(ptr_deref_1106_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1106_data_0;
      ov(31 downto 0) := iv;
      tmp1_1107 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1106_root_address_inst
    process(ptr_deref_1106_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1106_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1106_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1118_addr_0
    process(ptr_deref_1118_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1118_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1118_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1118_base_resize
    process(iNsTr_2_1115) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_2_1115;
      ov := iv(6 downto 0);
      ptr_deref_1118_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1118_gather_scatter
    process(ptr_deref_1118_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1118_data_0;
      ov(31 downto 0) := iv;
      tmp2_1119 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1118_root_address_inst
    process(ptr_deref_1118_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1118_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1118_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1197_addr_0
    process(ptr_deref_1197_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1197_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1197_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1197_base_resize
    process(arrayidx_1194) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_1194;
      ov := iv(13 downto 0);
      ptr_deref_1197_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1197_gather_scatter
    process(ptr_deref_1197_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1197_data_0;
      ov(63 downto 0) := iv;
      tmp9_1198 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1197_root_address_inst
    process(ptr_deref_1197_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1197_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1197_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1136_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp73_1135;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1136_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1136_branch_req_0,
          ack0 => if_stmt_1136_branch_ack_0,
          ack1 => if_stmt_1136_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1308_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond1_1307;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1308_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1308_branch_req_0,
          ack0 => if_stmt_1308_branch_ack_0,
          ack1 => if_stmt_1308_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u32_u32_1159_inst
    process(tmp77_1148) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp77_1148, type_cast_1158_wire_constant, tmp_var);
      tmp77x_xop_1160 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1169_inst
    process(iNsTr_4_1164) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_4_1164, type_cast_1168_wire_constant, tmp_var);
      xx_xop_1170 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1301_inst
    process(indvar_1180) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1180, type_cast_1300_wire_constant, tmp_var);
      indvarx_xnext_1302 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1306_inst
    process(indvarx_xnext_1302, tmp81_1177) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_1302, tmp81_1177, tmp_var);
      exitcond1_1307 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1147_inst
    process(mul3_1129) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul3_1129, type_cast_1146_wire_constant, tmp_var);
      tmp77_1148 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1207_inst
    process(tmp9_1198) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp9_1198, type_cast_1206_wire_constant, tmp_var);
      shr14_1208 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1217_inst
    process(tmp9_1198) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp9_1198, type_cast_1216_wire_constant, tmp_var);
      shr20_1218 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1227_inst
    process(tmp9_1198) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp9_1198, type_cast_1226_wire_constant, tmp_var);
      shr26_1228 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1237_inst
    process(tmp9_1198) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp9_1198, type_cast_1236_wire_constant, tmp_var);
      shr32_1238 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1247_inst
    process(tmp9_1198) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp9_1198, type_cast_1246_wire_constant, tmp_var);
      shr38_1248 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1257_inst
    process(tmp9_1198) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp9_1198, type_cast_1256_wire_constant, tmp_var);
      shr44_1258 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1267_inst
    process(tmp9_1198) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp9_1198, type_cast_1266_wire_constant, tmp_var);
      shr50_1268 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1123_inst
    process(tmp1_1107, tmp_1095) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp1_1107, tmp_1095, tmp_var);
      mul_1124 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1128_inst
    process(mul_1124, tmp2_1119) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_1124, tmp2_1119, tmp_var);
      mul3_1129 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1134_inst
    process(mul3_1129) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul3_1129, type_cast_1133_wire_constant, tmp_var);
      cmp73_1135 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1153_inst
    process(tmp77_1148) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp77_1148, type_cast_1152_wire_constant, tmp_var);
      tmp78_1154 <= tmp_var; --
    end process;
    -- shared split operator group (16) : array_obj_ref_1192_index_offset 
    ApIntAdd_group_16: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_1191_scaled;
      array_obj_ref_1192_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1192_index_offset_req_0;
      array_obj_ref_1192_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1192_index_offset_req_1;
      array_obj_ref_1192_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_16_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_16_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_16",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 16
    -- shared load operator group (0) : ptr_deref_1094_load_0 ptr_deref_1106_load_0 ptr_deref_1118_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(20 downto 0);
      signal data_out: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_1094_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_1106_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1118_load_0_req_0;
      ptr_deref_1094_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_1106_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1118_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_1094_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_1106_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1118_load_0_req_1;
      ptr_deref_1094_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_1106_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1118_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1094_word_address_0 & ptr_deref_1106_word_address_0 & ptr_deref_1118_word_address_0;
      ptr_deref_1094_data_0 <= data_out(95 downto 64);
      ptr_deref_1106_data_0 <= data_out(63 downto 32);
      ptr_deref_1118_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 7,
        num_reqs => 3,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(6 downto 0),
          mtag => memory_space_3_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 32,
        num_reqs => 3,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(31 downto 0),
          mtag => memory_space_3_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_1197_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1197_load_0_req_0;
      ptr_deref_1197_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1197_load_0_req_1;
      ptr_deref_1197_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1197_word_address_0;
      ptr_deref_1197_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_6_lr_req(0),
          mack => memory_space_6_lr_ack(0),
          maddr => memory_space_6_lr_addr(13 downto 0),
          mtag => memory_space_6_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_6_lc_req(0),
          mack => memory_space_6_lc_ack(0),
          mdata => memory_space_6_lc_data(63 downto 0),
          mtag => memory_space_6_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared outport operator group (0) : WPIPE_ConvTranspose_output_pipe_1273_inst WPIPE_ConvTranspose_output_pipe_1276_inst WPIPE_ConvTranspose_output_pipe_1279_inst WPIPE_ConvTranspose_output_pipe_1282_inst WPIPE_ConvTranspose_output_pipe_1285_inst WPIPE_ConvTranspose_output_pipe_1288_inst WPIPE_ConvTranspose_output_pipe_1291_inst WPIPE_ConvTranspose_output_pipe_1294_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 7 downto 0);
      signal update_req, update_ack : BooleanArray( 7 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 7 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 7 downto 0);
      signal guard_vector : std_logic_vector( 7 downto 0);
      constant inBUFs : IntegerArray(7 downto 0) := (7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(7 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false);
      constant guardBuffering: IntegerArray(7 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2);
      -- 
    begin -- 
      sample_req_unguarded(7) <= WPIPE_ConvTranspose_output_pipe_1273_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_ConvTranspose_output_pipe_1276_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_ConvTranspose_output_pipe_1279_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_ConvTranspose_output_pipe_1282_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_ConvTranspose_output_pipe_1285_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_ConvTranspose_output_pipe_1288_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_ConvTranspose_output_pipe_1291_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_ConvTranspose_output_pipe_1294_inst_req_0;
      WPIPE_ConvTranspose_output_pipe_1273_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_ConvTranspose_output_pipe_1276_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_ConvTranspose_output_pipe_1279_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_ConvTranspose_output_pipe_1282_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_ConvTranspose_output_pipe_1285_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_ConvTranspose_output_pipe_1288_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_ConvTranspose_output_pipe_1291_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_ConvTranspose_output_pipe_1294_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(7) <= WPIPE_ConvTranspose_output_pipe_1273_inst_req_1;
      update_req_unguarded(6) <= WPIPE_ConvTranspose_output_pipe_1276_inst_req_1;
      update_req_unguarded(5) <= WPIPE_ConvTranspose_output_pipe_1279_inst_req_1;
      update_req_unguarded(4) <= WPIPE_ConvTranspose_output_pipe_1282_inst_req_1;
      update_req_unguarded(3) <= WPIPE_ConvTranspose_output_pipe_1285_inst_req_1;
      update_req_unguarded(2) <= WPIPE_ConvTranspose_output_pipe_1288_inst_req_1;
      update_req_unguarded(1) <= WPIPE_ConvTranspose_output_pipe_1291_inst_req_1;
      update_req_unguarded(0) <= WPIPE_ConvTranspose_output_pipe_1294_inst_req_1;
      WPIPE_ConvTranspose_output_pipe_1273_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_ConvTranspose_output_pipe_1276_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_ConvTranspose_output_pipe_1279_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_ConvTranspose_output_pipe_1282_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_ConvTranspose_output_pipe_1285_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_ConvTranspose_output_pipe_1288_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_ConvTranspose_output_pipe_1291_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_ConvTranspose_output_pipe_1294_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      data_in <= conv53_1272 & conv47_1262 & conv41_1252 & conv35_1242 & conv29_1232 & conv23_1222 & conv17_1212 & conv_1202;
      ConvTranspose_output_pipe_write_0_gI: SplitGuardInterface generic map(name => "ConvTranspose_output_pipe_write_0_gI", nreqs => 8, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      ConvTranspose_output_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "ConvTranspose_output_pipe", data_width => 8, num_reqs => 8, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => ConvTranspose_output_pipe_pipe_write_req(0),
          oack => ConvTranspose_output_pipe_pipe_write_ack(0),
          odata => ConvTranspose_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end sendOutput_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity testConfigure is -- 
  generic (tag_length : integer); 
  port ( -- 
    ret_val_x_x : out  std_logic_vector(15 downto 0);
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(6 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sr_addr : out  std_logic_vector(10 downto 0);
    memory_space_5_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_5_sr_tag :  out  std_logic_vector(0 downto 0);
    memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_6_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_6_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_7_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_7_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_7_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_7_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_7_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_7_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(6 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_8_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_8_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_8_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_8_sr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_8_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_8_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_8_sc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(6 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_4_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_4_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_sc_tag :  in  std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity testConfigure;
architecture testConfigure_arch of testConfigure is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 16)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal ret_val_x_x_buffer :  std_logic_vector(15 downto 0);
  signal testConfigure_CP_0_start: Boolean;
  signal testConfigure_CP_0_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal ptr_deref_954_load_0_ack_0 : boolean;
  signal type_cast_1011_inst_req_0 : boolean;
  signal type_cast_829_inst_ack_1 : boolean;
  signal addr_of_1041_final_reg_req_0 : boolean;
  signal type_cast_901_inst_req_1 : boolean;
  signal array_obj_ref_1040_index_offset_ack_1 : boolean;
  signal array_obj_ref_1040_index_offset_req_1 : boolean;
  signal type_cast_1011_inst_ack_0 : boolean;
  signal ptr_deref_471_load_0_req_1 : boolean;
  signal ptr_deref_471_load_0_ack_1 : boolean;
  signal array_obj_ref_49_index_offset_ack_0 : boolean;
  signal array_obj_ref_49_index_offset_req_1 : boolean;
  signal array_obj_ref_49_index_offset_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_356_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_356_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_356_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_356_inst_req_0 : boolean;
  signal type_cast_883_inst_ack_1 : boolean;
  signal array_obj_ref_49_index_offset_req_0 : boolean;
  signal ptr_deref_459_load_0_ack_1 : boolean;
  signal array_obj_ref_119_index_offset_req_0 : boolean;
  signal array_obj_ref_119_index_offset_ack_0 : boolean;
  signal addr_of_1041_final_reg_ack_0 : boolean;
  signal array_obj_ref_119_index_offset_req_1 : boolean;
  signal addr_of_50_final_reg_req_0 : boolean;
  signal addr_of_50_final_reg_ack_0 : boolean;
  signal addr_of_50_final_reg_req_1 : boolean;
  signal addr_of_50_final_reg_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_53_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_53_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_53_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_53_inst_ack_1 : boolean;
  signal ptr_deref_459_load_0_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_843_inst_req_0 : boolean;
  signal type_cast_57_inst_req_0 : boolean;
  signal type_cast_57_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_861_inst_req_0 : boolean;
  signal type_cast_57_inst_req_1 : boolean;
  signal type_cast_57_inst_ack_1 : boolean;
  signal ptr_deref_60_store_0_req_0 : boolean;
  signal ptr_deref_60_store_0_ack_0 : boolean;
  signal ptr_deref_60_store_0_req_1 : boolean;
  signal ptr_deref_60_store_0_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_70_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_70_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_70_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_70_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_861_inst_req_1 : boolean;
  signal type_cast_74_inst_req_0 : boolean;
  signal type_cast_74_inst_ack_0 : boolean;
  signal type_cast_74_inst_req_1 : boolean;
  signal type_cast_74_inst_ack_1 : boolean;
  signal type_cast_883_inst_ack_0 : boolean;
  signal ptr_deref_82_store_0_req_0 : boolean;
  signal ptr_deref_82_store_0_ack_0 : boolean;
  signal ptr_deref_82_store_0_req_1 : boolean;
  signal ptr_deref_82_store_0_ack_1 : boolean;
  signal ptr_deref_471_load_0_ack_0 : boolean;
  signal ptr_deref_413_load_0_ack_1 : boolean;
  signal if_stmt_98_branch_req_0 : boolean;
  signal if_stmt_98_branch_ack_1 : boolean;
  signal ptr_deref_346_store_0_ack_1 : boolean;
  signal if_stmt_98_branch_ack_0 : boolean;
  signal ptr_deref_413_load_0_req_1 : boolean;
  signal ptr_deref_346_store_0_req_1 : boolean;
  signal ptr_deref_401_load_0_req_0 : boolean;
  signal ptr_deref_248_store_0_req_0 : boolean;
  signal ptr_deref_248_store_0_ack_0 : boolean;
  signal ptr_deref_248_store_0_req_1 : boolean;
  signal ptr_deref_248_store_0_ack_1 : boolean;
  signal type_cast_360_inst_ack_1 : boolean;
  signal type_cast_360_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_258_inst_req_0 : boolean;
  signal array_obj_ref_119_index_offset_ack_1 : boolean;
  signal addr_of_120_final_reg_req_0 : boolean;
  signal addr_of_120_final_reg_ack_0 : boolean;
  signal addr_of_120_final_reg_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_861_inst_ack_1 : boolean;
  signal addr_of_120_final_reg_ack_1 : boolean;
  signal ptr_deref_471_load_0_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_123_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_123_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_123_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_123_inst_ack_1 : boolean;
  signal ptr_deref_942_load_0_req_0 : boolean;
  signal type_cast_127_inst_req_0 : boolean;
  signal type_cast_127_inst_ack_0 : boolean;
  signal type_cast_127_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_843_inst_req_1 : boolean;
  signal type_cast_127_inst_ack_1 : boolean;
  signal ptr_deref_376_store_0_req_1 : boolean;
  signal ptr_deref_413_load_0_ack_0 : boolean;
  signal ptr_deref_942_load_0_ack_0 : boolean;
  signal ptr_deref_130_store_0_req_0 : boolean;
  signal ptr_deref_130_store_0_ack_0 : boolean;
  signal ptr_deref_376_store_0_ack_1 : boolean;
  signal ptr_deref_130_store_0_req_1 : boolean;
  signal ptr_deref_130_store_0_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_140_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_140_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_140_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_140_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_843_inst_ack_0 : boolean;
  signal ptr_deref_435_load_0_ack_1 : boolean;
  signal type_cast_144_inst_req_0 : boolean;
  signal type_cast_144_inst_ack_0 : boolean;
  signal type_cast_144_inst_req_1 : boolean;
  signal type_cast_144_inst_ack_1 : boolean;
  signal ptr_deref_413_load_0_req_0 : boolean;
  signal if_stmt_984_branch_req_0 : boolean;
  signal type_cast_883_inst_req_0 : boolean;
  signal type_cast_883_inst_req_1 : boolean;
  signal ptr_deref_435_load_0_req_1 : boolean;
  signal ptr_deref_152_store_0_req_0 : boolean;
  signal ptr_deref_152_store_0_ack_0 : boolean;
  signal ptr_deref_152_store_0_req_1 : boolean;
  signal ptr_deref_152_store_0_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_843_inst_ack_1 : boolean;
  signal if_stmt_167_branch_req_0 : boolean;
  signal if_stmt_167_branch_ack_1 : boolean;
  signal if_stmt_167_branch_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_175_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_175_inst_ack_0 : boolean;
  signal ptr_deref_447_load_0_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_175_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_175_inst_ack_1 : boolean;
  signal ptr_deref_447_load_0_req_1 : boolean;
  signal ptr_deref_954_load_0_req_0 : boolean;
  signal ptr_deref_346_store_0_ack_0 : boolean;
  signal ptr_deref_389_load_0_ack_1 : boolean;
  signal ptr_deref_389_load_0_req_1 : boolean;
  signal addr_of_196_final_reg_req_0 : boolean;
  signal ptr_deref_401_load_0_ack_1 : boolean;
  signal addr_of_196_final_reg_ack_0 : boolean;
  signal addr_of_196_final_reg_req_1 : boolean;
  signal addr_of_196_final_reg_ack_1 : boolean;
  signal ptr_deref_401_load_0_req_1 : boolean;
  signal ptr_deref_199_store_0_req_0 : boolean;
  signal ptr_deref_199_store_0_ack_0 : boolean;
  signal ptr_deref_346_store_0_req_0 : boolean;
  signal ptr_deref_376_store_0_ack_0 : boolean;
  signal ptr_deref_199_store_0_req_1 : boolean;
  signal ptr_deref_199_store_0_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_861_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_203_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_203_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_203_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_203_inst_ack_1 : boolean;
  signal if_stmt_217_branch_req_0 : boolean;
  signal if_stmt_217_branch_ack_1 : boolean;
  signal if_stmt_217_branch_ack_0 : boolean;
  signal ptr_deref_376_store_0_req_0 : boolean;
  signal ptr_deref_435_load_0_ack_0 : boolean;
  signal STORE_padding_229_store_0_req_0 : boolean;
  signal STORE_padding_229_store_0_ack_0 : boolean;
  signal STORE_padding_229_store_0_req_1 : boolean;
  signal STORE_padding_229_store_0_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_233_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_233_inst_ack_0 : boolean;
  signal ptr_deref_447_load_0_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_233_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_233_inst_ack_1 : boolean;
  signal ptr_deref_389_load_0_ack_0 : boolean;
  signal ptr_deref_389_load_0_req_0 : boolean;
  signal type_cast_237_inst_req_0 : boolean;
  signal type_cast_237_inst_ack_0 : boolean;
  signal ptr_deref_435_load_0_req_0 : boolean;
  signal type_cast_237_inst_req_1 : boolean;
  signal type_cast_237_inst_ack_1 : boolean;
  signal if_stmt_984_branch_ack_1 : boolean;
  signal ptr_deref_447_load_0_req_0 : boolean;
  signal ptr_deref_401_load_0_ack_0 : boolean;
  signal ptr_deref_459_load_0_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_258_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_258_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_258_inst_ack_1 : boolean;
  signal type_cast_901_inst_ack_1 : boolean;
  signal type_cast_262_inst_req_0 : boolean;
  signal type_cast_262_inst_ack_0 : boolean;
  signal type_cast_262_inst_req_1 : boolean;
  signal type_cast_262_inst_ack_1 : boolean;
  signal type_cast_360_inst_ack_0 : boolean;
  signal ptr_deref_942_load_0_req_1 : boolean;
  signal type_cast_360_inst_req_0 : boolean;
  signal ptr_deref_459_load_0_req_0 : boolean;
  signal ptr_deref_278_store_0_req_0 : boolean;
  signal ptr_deref_942_load_0_ack_1 : boolean;
  signal ptr_deref_278_store_0_ack_0 : boolean;
  signal ptr_deref_278_store_0_req_1 : boolean;
  signal ptr_deref_278_store_0_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_897_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_282_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_282_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_282_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_282_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_897_inst_ack_0 : boolean;
  signal type_cast_286_inst_req_0 : boolean;
  signal type_cast_286_inst_ack_0 : boolean;
  signal type_cast_286_inst_req_1 : boolean;
  signal type_cast_286_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_897_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_897_inst_ack_1 : boolean;
  signal ptr_deref_966_load_0_req_0 : boolean;
  signal ptr_deref_297_store_0_req_0 : boolean;
  signal ptr_deref_297_store_0_ack_0 : boolean;
  signal ptr_deref_297_store_0_req_1 : boolean;
  signal ptr_deref_297_store_0_ack_1 : boolean;
  signal addr_of_1041_final_reg_req_1 : boolean;
  signal type_cast_847_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_307_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_307_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_307_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_307_inst_ack_1 : boolean;
  signal type_cast_311_inst_req_0 : boolean;
  signal type_cast_311_inst_ack_0 : boolean;
  signal type_cast_311_inst_req_1 : boolean;
  signal type_cast_311_inst_ack_1 : boolean;
  signal ptr_deref_327_store_0_req_0 : boolean;
  signal ptr_deref_327_store_0_ack_0 : boolean;
  signal ptr_deref_327_store_0_req_1 : boolean;
  signal ptr_deref_327_store_0_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_331_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_331_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_331_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_331_inst_ack_1 : boolean;
  signal type_cast_335_inst_req_0 : boolean;
  signal type_cast_335_inst_ack_0 : boolean;
  signal type_cast_335_inst_req_1 : boolean;
  signal type_cast_335_inst_ack_1 : boolean;
  signal if_stmt_494_branch_req_0 : boolean;
  signal if_stmt_494_branch_ack_1 : boolean;
  signal if_stmt_494_branch_ack_0 : boolean;
  signal type_cast_901_inst_ack_0 : boolean;
  signal type_cast_847_inst_ack_1 : boolean;
  signal type_cast_847_inst_req_1 : boolean;
  signal if_stmt_509_branch_req_0 : boolean;
  signal if_stmt_509_branch_ack_1 : boolean;
  signal if_stmt_509_branch_ack_0 : boolean;
  signal type_cast_901_inst_req_0 : boolean;
  signal type_cast_536_inst_req_0 : boolean;
  signal type_cast_536_inst_ack_0 : boolean;
  signal type_cast_536_inst_req_1 : boolean;
  signal type_cast_536_inst_ack_1 : boolean;
  signal type_cast_847_inst_ack_0 : boolean;
  signal if_stmt_923_branch_ack_0 : boolean;
  signal array_obj_ref_1040_index_offset_ack_0 : boolean;
  signal array_obj_ref_565_index_offset_req_0 : boolean;
  signal array_obj_ref_565_index_offset_ack_0 : boolean;
  signal array_obj_ref_565_index_offset_req_1 : boolean;
  signal array_obj_ref_565_index_offset_ack_1 : boolean;
  signal array_obj_ref_1040_index_offset_req_0 : boolean;
  signal if_stmt_923_branch_ack_1 : boolean;
  signal addr_of_566_final_reg_req_0 : boolean;
  signal addr_of_566_final_reg_ack_0 : boolean;
  signal addr_of_566_final_reg_req_1 : boolean;
  signal addr_of_566_final_reg_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_879_inst_ack_1 : boolean;
  signal if_stmt_923_branch_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_569_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_569_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_879_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_569_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_569_inst_ack_1 : boolean;
  signal addr_of_1041_final_reg_ack_1 : boolean;
  signal type_cast_573_inst_req_0 : boolean;
  signal type_cast_573_inst_ack_0 : boolean;
  signal type_cast_573_inst_req_1 : boolean;
  signal type_cast_573_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_582_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_582_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_582_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_582_inst_ack_1 : boolean;
  signal type_cast_586_inst_req_0 : boolean;
  signal type_cast_586_inst_ack_0 : boolean;
  signal type_cast_586_inst_req_1 : boolean;
  signal type_cast_586_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_600_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_600_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_879_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_600_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_600_inst_ack_1 : boolean;
  signal ptr_deref_909_store_0_ack_1 : boolean;
  signal type_cast_604_inst_req_0 : boolean;
  signal type_cast_604_inst_ack_0 : boolean;
  signal type_cast_604_inst_req_1 : boolean;
  signal type_cast_604_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_879_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_618_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_618_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_618_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_618_inst_ack_1 : boolean;
  signal ptr_deref_909_store_0_req_1 : boolean;
  signal type_cast_622_inst_req_0 : boolean;
  signal type_cast_622_inst_ack_0 : boolean;
  signal type_cast_622_inst_req_1 : boolean;
  signal type_cast_622_inst_ack_1 : boolean;
  signal if_stmt_984_branch_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_636_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_636_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_636_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_636_inst_ack_1 : boolean;
  signal type_cast_640_inst_req_0 : boolean;
  signal type_cast_640_inst_ack_0 : boolean;
  signal type_cast_640_inst_req_1 : boolean;
  signal type_cast_640_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_654_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_654_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_654_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_654_inst_ack_1 : boolean;
  signal type_cast_658_inst_req_0 : boolean;
  signal type_cast_658_inst_ack_0 : boolean;
  signal type_cast_658_inst_req_1 : boolean;
  signal type_cast_658_inst_ack_1 : boolean;
  signal type_cast_865_inst_ack_1 : boolean;
  signal ptr_deref_966_load_0_ack_1 : boolean;
  signal ptr_deref_909_store_0_ack_0 : boolean;
  signal ptr_deref_909_store_0_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_672_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_672_inst_ack_0 : boolean;
  signal type_cast_865_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_672_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_672_inst_ack_1 : boolean;
  signal ptr_deref_966_load_0_req_1 : boolean;
  signal type_cast_676_inst_req_0 : boolean;
  signal type_cast_676_inst_ack_0 : boolean;
  signal type_cast_676_inst_req_1 : boolean;
  signal type_cast_676_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_690_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_690_inst_ack_0 : boolean;
  signal type_cast_865_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_690_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_690_inst_ack_1 : boolean;
  signal type_cast_865_inst_req_0 : boolean;
  signal type_cast_694_inst_req_0 : boolean;
  signal type_cast_694_inst_ack_0 : boolean;
  signal type_cast_694_inst_req_1 : boolean;
  signal ptr_deref_954_load_0_ack_1 : boolean;
  signal type_cast_694_inst_ack_1 : boolean;
  signal ptr_deref_966_load_0_ack_0 : boolean;
  signal ptr_deref_954_load_0_req_1 : boolean;
  signal ptr_deref_702_store_0_req_0 : boolean;
  signal ptr_deref_702_store_0_ack_0 : boolean;
  signal type_cast_829_inst_req_1 : boolean;
  signal ptr_deref_702_store_0_req_1 : boolean;
  signal ptr_deref_702_store_0_ack_1 : boolean;
  signal type_cast_1011_inst_ack_1 : boolean;
  signal type_cast_1011_inst_req_1 : boolean;
  signal if_stmt_716_branch_req_0 : boolean;
  signal if_stmt_716_branch_ack_1 : boolean;
  signal if_stmt_716_branch_ack_0 : boolean;
  signal type_cast_743_inst_req_0 : boolean;
  signal type_cast_743_inst_ack_0 : boolean;
  signal type_cast_743_inst_req_1 : boolean;
  signal type_cast_743_inst_ack_1 : boolean;
  signal array_obj_ref_772_index_offset_req_0 : boolean;
  signal array_obj_ref_772_index_offset_ack_0 : boolean;
  signal array_obj_ref_772_index_offset_req_1 : boolean;
  signal array_obj_ref_772_index_offset_ack_1 : boolean;
  signal addr_of_773_final_reg_req_0 : boolean;
  signal addr_of_773_final_reg_ack_0 : boolean;
  signal addr_of_773_final_reg_req_1 : boolean;
  signal addr_of_773_final_reg_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_776_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_776_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_776_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_776_inst_ack_1 : boolean;
  signal type_cast_780_inst_req_0 : boolean;
  signal type_cast_780_inst_ack_0 : boolean;
  signal type_cast_780_inst_req_1 : boolean;
  signal type_cast_780_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_789_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_789_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_789_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_789_inst_ack_1 : boolean;
  signal type_cast_793_inst_req_0 : boolean;
  signal type_cast_793_inst_ack_0 : boolean;
  signal type_cast_793_inst_req_1 : boolean;
  signal type_cast_793_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_807_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_807_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_807_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_807_inst_ack_1 : boolean;
  signal type_cast_811_inst_req_0 : boolean;
  signal type_cast_811_inst_ack_0 : boolean;
  signal type_cast_811_inst_req_1 : boolean;
  signal type_cast_811_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_825_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_825_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_825_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_825_inst_ack_1 : boolean;
  signal type_cast_829_inst_req_0 : boolean;
  signal type_cast_829_inst_ack_0 : boolean;
  signal ptr_deref_1044_store_0_req_0 : boolean;
  signal ptr_deref_1044_store_0_ack_0 : boolean;
  signal ptr_deref_1044_store_0_req_1 : boolean;
  signal ptr_deref_1044_store_0_ack_1 : boolean;
  signal if_stmt_1059_branch_req_0 : boolean;
  signal if_stmt_1059_branch_ack_1 : boolean;
  signal if_stmt_1059_branch_ack_0 : boolean;
  signal phi_stmt_37_req_0 : boolean;
  signal type_cast_43_inst_req_0 : boolean;
  signal type_cast_43_inst_ack_0 : boolean;
  signal type_cast_43_inst_req_1 : boolean;
  signal type_cast_43_inst_ack_1 : boolean;
  signal phi_stmt_37_req_1 : boolean;
  signal phi_stmt_37_ack_0 : boolean;
  signal type_cast_110_inst_req_0 : boolean;
  signal type_cast_110_inst_ack_0 : boolean;
  signal type_cast_110_inst_req_1 : boolean;
  signal type_cast_110_inst_ack_1 : boolean;
  signal phi_stmt_107_req_0 : boolean;
  signal phi_stmt_107_req_1 : boolean;
  signal phi_stmt_107_ack_0 : boolean;
  signal phi_stmt_179_req_0 : boolean;
  signal type_cast_189_inst_req_0 : boolean;
  signal type_cast_189_inst_ack_0 : boolean;
  signal type_cast_189_inst_req_1 : boolean;
  signal type_cast_189_inst_ack_1 : boolean;
  signal phi_stmt_186_req_0 : boolean;
  signal type_cast_185_inst_req_0 : boolean;
  signal type_cast_185_inst_ack_0 : boolean;
  signal type_cast_185_inst_req_1 : boolean;
  signal type_cast_185_inst_ack_1 : boolean;
  signal phi_stmt_179_req_1 : boolean;
  signal type_cast_191_inst_req_0 : boolean;
  signal type_cast_191_inst_ack_0 : boolean;
  signal type_cast_191_inst_req_1 : boolean;
  signal type_cast_191_inst_ack_1 : boolean;
  signal phi_stmt_186_req_1 : boolean;
  signal phi_stmt_179_ack_0 : boolean;
  signal phi_stmt_186_ack_0 : boolean;
  signal type_cast_227_inst_req_0 : boolean;
  signal type_cast_227_inst_ack_0 : boolean;
  signal type_cast_227_inst_req_1 : boolean;
  signal type_cast_227_inst_ack_1 : boolean;
  signal phi_stmt_224_req_0 : boolean;
  signal phi_stmt_224_ack_0 : boolean;
  signal phi_stmt_553_req_0 : boolean;
  signal type_cast_559_inst_req_0 : boolean;
  signal type_cast_559_inst_ack_0 : boolean;
  signal type_cast_559_inst_req_1 : boolean;
  signal type_cast_559_inst_ack_1 : boolean;
  signal phi_stmt_553_req_1 : boolean;
  signal phi_stmt_553_ack_0 : boolean;
  signal phi_stmt_760_req_0 : boolean;
  signal type_cast_766_inst_req_0 : boolean;
  signal type_cast_766_inst_ack_0 : boolean;
  signal type_cast_766_inst_req_1 : boolean;
  signal type_cast_766_inst_ack_1 : boolean;
  signal phi_stmt_760_req_1 : boolean;
  signal phi_stmt_760_ack_0 : boolean;
  signal phi_stmt_1028_req_0 : boolean;
  signal type_cast_1034_inst_req_0 : boolean;
  signal type_cast_1034_inst_ack_0 : boolean;
  signal type_cast_1034_inst_req_1 : boolean;
  signal type_cast_1034_inst_ack_1 : boolean;
  signal phi_stmt_1028_req_1 : boolean;
  signal phi_stmt_1028_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "testConfigure_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  testConfigure_CP_0_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "testConfigure_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 16) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  ret_val_x_x_buffer <= "0000000000000001";
  out_buffer_data_in(15 downto 0) <= ret_val_x_x_buffer;
  ret_val_x_x <= out_buffer_data_out(15 downto 0);
  out_buffer_data_in(tag_length + 15 downto 16) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 15 downto 16);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= testConfigure_CP_0_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= testConfigure_CP_0_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= testConfigure_CP_0_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  testConfigure_CP_0: Block -- control-path 
    signal testConfigure_CP_0_elements: BooleanArray(286 downto 0);
    -- 
  begin -- 
    testConfigure_CP_0_elements(0) <= testConfigure_CP_0_start;
    testConfigure_CP_0_symbol <= testConfigure_CP_0_elements(286);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	233 
    -- CP-element group 0:  members (7) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_34/$entry
      -- CP-element group 0: 	 branch_block_stmt_34/branch_block_stmt_34__entry__
      -- CP-element group 0: 	 branch_block_stmt_34/bbx_xnph246_forx_xbody
      -- CP-element group 0: 	 branch_block_stmt_34/bbx_xnph246_forx_xbody_PhiReq/$entry
      -- CP-element group 0: 	 branch_block_stmt_34/bbx_xnph246_forx_xbody_PhiReq/phi_stmt_37/$entry
      -- CP-element group 0: 	 branch_block_stmt_34/bbx_xnph246_forx_xbody_PhiReq/phi_stmt_37/phi_stmt_37_sources/$entry
      -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	238 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	20 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/array_obj_ref_49_final_index_sum_regn_Sample/ack
      -- CP-element group 1: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/array_obj_ref_49_final_index_sum_regn_sample_complete
      -- CP-element group 1: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/array_obj_ref_49_final_index_sum_regn_Sample/$exit
      -- 
    ack_120_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_49_index_offset_ack_0, ack => testConfigure_CP_0_elements(1)); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	238 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (11) 
      -- CP-element group 2: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/array_obj_ref_49_final_index_sum_regn_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/array_obj_ref_49_final_index_sum_regn_Update/ack
      -- CP-element group 2: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/addr_of_50_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/array_obj_ref_49_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/array_obj_ref_49_offset_calculated
      -- CP-element group 2: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/array_obj_ref_49_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/array_obj_ref_49_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/array_obj_ref_49_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/array_obj_ref_49_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/addr_of_50_request/$entry
      -- CP-element group 2: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/addr_of_50_request/req
      -- 
    ack_125_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_49_index_offset_ack_1, ack => testConfigure_CP_0_elements(2)); -- 
    req_134_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_134_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(2), ack => addr_of_50_final_reg_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/addr_of_50_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/addr_of_50_request/$exit
      -- CP-element group 3: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/addr_of_50_request/ack
      -- 
    ack_135_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_50_final_reg_ack_0, ack => testConfigure_CP_0_elements(3)); -- 
    -- CP-element group 4:  fork  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	238 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	16 
    -- CP-element group 4: 	9 
    -- CP-element group 4:  members (35) 
      -- CP-element group 4: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/addr_of_50_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/addr_of_50_complete/$exit
      -- CP-element group 4: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/addr_of_50_complete/ack
      -- CP-element group 4: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_60_base_address_calculated
      -- CP-element group 4: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_60_word_address_calculated
      -- CP-element group 4: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_60_root_address_calculated
      -- CP-element group 4: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_60_base_address_resized
      -- CP-element group 4: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_60_base_addr_resize/$entry
      -- CP-element group 4: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_60_base_addr_resize/$exit
      -- CP-element group 4: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_60_base_addr_resize/base_resize_req
      -- CP-element group 4: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_60_base_addr_resize/base_resize_ack
      -- CP-element group 4: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_60_base_plus_offset/$entry
      -- CP-element group 4: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_60_base_plus_offset/$exit
      -- CP-element group 4: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_60_base_plus_offset/sum_rename_req
      -- CP-element group 4: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_60_base_plus_offset/sum_rename_ack
      -- CP-element group 4: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_60_word_addrgen/$entry
      -- CP-element group 4: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_60_word_addrgen/$exit
      -- CP-element group 4: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_60_word_addrgen/root_register_req
      -- CP-element group 4: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_60_word_addrgen/root_register_ack
      -- CP-element group 4: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_82_base_address_calculated
      -- CP-element group 4: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_82_word_address_calculated
      -- CP-element group 4: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_82_root_address_calculated
      -- CP-element group 4: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_82_base_address_resized
      -- CP-element group 4: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_82_base_addr_resize/$entry
      -- CP-element group 4: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_82_base_addr_resize/$exit
      -- CP-element group 4: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_82_base_addr_resize/base_resize_req
      -- CP-element group 4: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_82_base_addr_resize/base_resize_ack
      -- CP-element group 4: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_82_base_plus_offset/$entry
      -- CP-element group 4: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_82_base_plus_offset/$exit
      -- CP-element group 4: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_82_base_plus_offset/sum_rename_req
      -- CP-element group 4: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_82_base_plus_offset/sum_rename_ack
      -- CP-element group 4: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_82_word_addrgen/$entry
      -- CP-element group 4: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_82_word_addrgen/$exit
      -- CP-element group 4: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_82_word_addrgen/root_register_req
      -- CP-element group 4: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_82_word_addrgen/root_register_ack
      -- 
    ack_140_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_50_final_reg_ack_1, ack => testConfigure_CP_0_elements(4)); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	238 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/RPIPE_ConvTranspose_input_pipe_53_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/RPIPE_ConvTranspose_input_pipe_53_update_start_
      -- CP-element group 5: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/RPIPE_ConvTranspose_input_pipe_53_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/RPIPE_ConvTranspose_input_pipe_53_Sample/ra
      -- CP-element group 5: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/RPIPE_ConvTranspose_input_pipe_53_Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/RPIPE_ConvTranspose_input_pipe_53_Update/cr
      -- 
    ra_149_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_53_inst_ack_0, ack => testConfigure_CP_0_elements(5)); -- 
    cr_153_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_153_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(5), ack => RPIPE_ConvTranspose_input_pipe_53_inst_req_1); -- 
    -- CP-element group 6:  fork  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	12 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/RPIPE_ConvTranspose_input_pipe_53_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/RPIPE_ConvTranspose_input_pipe_53_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/RPIPE_ConvTranspose_input_pipe_53_Update/ca
      -- CP-element group 6: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/type_cast_57_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/type_cast_57_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/type_cast_57_Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/RPIPE_ConvTranspose_input_pipe_70_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/RPIPE_ConvTranspose_input_pipe_70_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/RPIPE_ConvTranspose_input_pipe_70_Sample/rr
      -- 
    ca_154_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_53_inst_ack_1, ack => testConfigure_CP_0_elements(6)); -- 
    rr_226_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_226_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(6), ack => RPIPE_ConvTranspose_input_pipe_70_inst_req_0); -- 
    rr_162_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_162_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(6), ack => type_cast_57_inst_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/type_cast_57_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/type_cast_57_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/type_cast_57_Sample/ra
      -- 
    ra_163_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_57_inst_ack_0, ack => testConfigure_CP_0_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	238 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/type_cast_57_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/type_cast_57_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/type_cast_57_Update/ca
      -- 
    ca_168_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_57_inst_ack_1, ack => testConfigure_CP_0_elements(8)); -- 
    -- CP-element group 9:  join  transition  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	4 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (9) 
      -- CP-element group 9: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_60_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_60_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_60_Sample/ptr_deref_60_Split/$entry
      -- CP-element group 9: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_60_Sample/ptr_deref_60_Split/$exit
      -- CP-element group 9: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_60_Sample/ptr_deref_60_Split/split_req
      -- CP-element group 9: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_60_Sample/ptr_deref_60_Split/split_ack
      -- CP-element group 9: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_60_Sample/word_access_start/$entry
      -- CP-element group 9: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_60_Sample/word_access_start/word_0/$entry
      -- CP-element group 9: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_60_Sample/word_access_start/word_0/rr
      -- 
    rr_206_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_206_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(9), ack => ptr_deref_60_store_0_req_0); -- 
    testConfigure_cp_element_group_9: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "testConfigure_cp_element_group_9"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(4) & testConfigure_CP_0_elements(8);
      gj_testConfigure_cp_element_group_9 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(9), clk => clk, reset => reset); --
    end block;
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	19 
    -- CP-element group 10:  members (5) 
      -- CP-element group 10: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_60_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_60_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_60_Sample/word_access_start/$exit
      -- CP-element group 10: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_60_Sample/word_access_start/word_0/$exit
      -- CP-element group 10: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_60_Sample/word_access_start/word_0/ra
      -- 
    ra_207_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_60_store_0_ack_0, ack => testConfigure_CP_0_elements(10)); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	238 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	20 
    -- CP-element group 11:  members (5) 
      -- CP-element group 11: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_60_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_60_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_60_Update/word_access_complete/$exit
      -- CP-element group 11: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_60_Update/word_access_complete/word_0/$exit
      -- CP-element group 11: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_60_Update/word_access_complete/word_0/ca
      -- 
    ca_218_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_60_store_0_ack_1, ack => testConfigure_CP_0_elements(11)); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	6 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/RPIPE_ConvTranspose_input_pipe_70_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/RPIPE_ConvTranspose_input_pipe_70_update_start_
      -- CP-element group 12: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/RPIPE_ConvTranspose_input_pipe_70_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/RPIPE_ConvTranspose_input_pipe_70_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/RPIPE_ConvTranspose_input_pipe_70_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/RPIPE_ConvTranspose_input_pipe_70_Update/cr
      -- 
    ra_227_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_70_inst_ack_0, ack => testConfigure_CP_0_elements(12)); -- 
    cr_231_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_231_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(12), ack => RPIPE_ConvTranspose_input_pipe_70_inst_req_1); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/RPIPE_ConvTranspose_input_pipe_70_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/RPIPE_ConvTranspose_input_pipe_70_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/RPIPE_ConvTranspose_input_pipe_70_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/type_cast_74_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/type_cast_74_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/type_cast_74_Sample/rr
      -- 
    ca_232_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_70_inst_ack_1, ack => testConfigure_CP_0_elements(13)); -- 
    rr_240_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_240_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(13), ack => type_cast_74_inst_req_0); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/type_cast_74_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/type_cast_74_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/type_cast_74_Sample/ra
      -- 
    ra_241_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_74_inst_ack_0, ack => testConfigure_CP_0_elements(14)); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	238 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/type_cast_74_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/type_cast_74_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/type_cast_74_Update/ca
      -- 
    ca_246_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_74_inst_ack_1, ack => testConfigure_CP_0_elements(15)); -- 
    -- CP-element group 16:  join  transition  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: 	19 
    -- CP-element group 16: 	4 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (9) 
      -- CP-element group 16: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_82_sample_start_
      -- CP-element group 16: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_82_Sample/$entry
      -- CP-element group 16: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_82_Sample/ptr_deref_82_Split/$entry
      -- CP-element group 16: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_82_Sample/ptr_deref_82_Split/$exit
      -- CP-element group 16: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_82_Sample/ptr_deref_82_Split/split_req
      -- CP-element group 16: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_82_Sample/ptr_deref_82_Split/split_ack
      -- CP-element group 16: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_82_Sample/word_access_start/$entry
      -- CP-element group 16: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_82_Sample/word_access_start/word_0/$entry
      -- CP-element group 16: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_82_Sample/word_access_start/word_0/rr
      -- 
    rr_284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(16), ack => ptr_deref_82_store_0_req_0); -- 
    testConfigure_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(15) & testConfigure_CP_0_elements(19) & testConfigure_CP_0_elements(4);
      gj_testConfigure_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (5) 
      -- CP-element group 17: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_82_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_82_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_82_Sample/word_access_start/$exit
      -- CP-element group 17: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_82_Sample/word_access_start/word_0/$exit
      -- CP-element group 17: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_82_Sample/word_access_start/word_0/ra
      -- 
    ra_285_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_82_store_0_ack_0, ack => testConfigure_CP_0_elements(17)); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	238 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	20 
    -- CP-element group 18:  members (5) 
      -- CP-element group 18: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_82_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_82_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_82_Update/word_access_complete/$exit
      -- CP-element group 18: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_82_Update/word_access_complete/word_0/$exit
      -- CP-element group 18: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_82_Update/word_access_complete/word_0/ca
      -- 
    ca_296_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_82_store_0_ack_1, ack => testConfigure_CP_0_elements(18)); -- 
    -- CP-element group 19:  transition  delay-element  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	10 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	16 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_60_ptr_deref_82_delay
      -- 
    -- Element group testConfigure_CP_0_elements(19) is a control-delay.
    cp_element_19_delay: control_delay_element  generic map(name => " 19_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(10), ack => testConfigure_CP_0_elements(19), clk => clk, reset =>reset);
    -- CP-element group 20:  branch  join  transition  place  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	11 
    -- CP-element group 20: 	18 
    -- CP-element group 20: 	1 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20: 	22 
    -- CP-element group 20:  members (10) 
      -- CP-element group 20: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97__exit__
      -- CP-element group 20: 	 branch_block_stmt_34/if_stmt_98__entry__
      -- CP-element group 20: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/$exit
      -- CP-element group 20: 	 branch_block_stmt_34/if_stmt_98_dead_link/$entry
      -- CP-element group 20: 	 branch_block_stmt_34/if_stmt_98_eval_test/$entry
      -- CP-element group 20: 	 branch_block_stmt_34/if_stmt_98_eval_test/$exit
      -- CP-element group 20: 	 branch_block_stmt_34/if_stmt_98_eval_test/branch_req
      -- CP-element group 20: 	 branch_block_stmt_34/R_exitcond5_99_place
      -- CP-element group 20: 	 branch_block_stmt_34/if_stmt_98_if_link/$entry
      -- CP-element group 20: 	 branch_block_stmt_34/if_stmt_98_else_link/$entry
      -- 
    branch_req_305_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_305_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(20), ack => if_stmt_98_branch_req_0); -- 
    testConfigure_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(11) & testConfigure_CP_0_elements(18) & testConfigure_CP_0_elements(1);
      gj_testConfigure_cp_element_group_20 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  merge  transition  place  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	242 
    -- CP-element group 21:  members (14) 
      -- CP-element group 21: 	 branch_block_stmt_34/merge_stmt_104__exit__
      -- CP-element group 21: 	 branch_block_stmt_34/forx_xbody16x_xpreheader_forx_xbody16
      -- CP-element group 21: 	 branch_block_stmt_34/if_stmt_98_if_link/$exit
      -- CP-element group 21: 	 branch_block_stmt_34/if_stmt_98_if_link/if_choice_transition
      -- CP-element group 21: 	 branch_block_stmt_34/forx_xbody_forx_xbody16x_xpreheader
      -- CP-element group 21: 	 branch_block_stmt_34/forx_xbody_forx_xbody16x_xpreheader_PhiReq/$entry
      -- CP-element group 21: 	 branch_block_stmt_34/forx_xbody_forx_xbody16x_xpreheader_PhiReq/$exit
      -- CP-element group 21: 	 branch_block_stmt_34/merge_stmt_104_PhiReqMerge
      -- CP-element group 21: 	 branch_block_stmt_34/merge_stmt_104_PhiAck/$entry
      -- CP-element group 21: 	 branch_block_stmt_34/merge_stmt_104_PhiAck/$exit
      -- CP-element group 21: 	 branch_block_stmt_34/merge_stmt_104_PhiAck/dummy
      -- CP-element group 21: 	 branch_block_stmt_34/forx_xbody16x_xpreheader_forx_xbody16_PhiReq/$entry
      -- CP-element group 21: 	 branch_block_stmt_34/forx_xbody16x_xpreheader_forx_xbody16_PhiReq/phi_stmt_107/$entry
      -- CP-element group 21: 	 branch_block_stmt_34/forx_xbody16x_xpreheader_forx_xbody16_PhiReq/phi_stmt_107/phi_stmt_107_sources/$entry
      -- 
    if_choice_transition_310_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_98_branch_ack_1, ack => testConfigure_CP_0_elements(21)); -- 
    -- CP-element group 22:  fork  transition  place  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	20 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	234 
    -- CP-element group 22: 	235 
    -- CP-element group 22:  members (12) 
      -- CP-element group 22: 	 branch_block_stmt_34/if_stmt_98_else_link/$exit
      -- CP-element group 22: 	 branch_block_stmt_34/if_stmt_98_else_link/else_choice_transition
      -- CP-element group 22: 	 branch_block_stmt_34/forx_xbody_forx_xbody
      -- CP-element group 22: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 22: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_37/$entry
      -- CP-element group 22: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_37/phi_stmt_37_sources/$entry
      -- CP-element group 22: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_37/phi_stmt_37_sources/type_cast_43/$entry
      -- CP-element group 22: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_37/phi_stmt_37_sources/type_cast_43/SplitProtocol/$entry
      -- CP-element group 22: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_37/phi_stmt_37_sources/type_cast_43/SplitProtocol/Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_37/phi_stmt_37_sources/type_cast_43/SplitProtocol/Sample/rr
      -- CP-element group 22: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_37/phi_stmt_37_sources/type_cast_43/SplitProtocol/Update/$entry
      -- CP-element group 22: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_37/phi_stmt_37_sources/type_cast_43/SplitProtocol/Update/cr
      -- 
    else_choice_transition_314_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_98_branch_ack_0, ack => testConfigure_CP_0_elements(22)); -- 
    rr_2641_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2641_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(22), ack => type_cast_43_inst_req_0); -- 
    cr_2646_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2646_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(22), ack => type_cast_43_inst_req_1); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	244 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	42 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/array_obj_ref_119_final_index_sum_regn_sample_complete
      -- CP-element group 23: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/array_obj_ref_119_final_index_sum_regn_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/array_obj_ref_119_final_index_sum_regn_Sample/ack
      -- 
    ack_345_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_119_index_offset_ack_0, ack => testConfigure_CP_0_elements(23)); -- 
    -- CP-element group 24:  transition  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	244 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (11) 
      -- CP-element group 24: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/array_obj_ref_119_final_index_sum_regn_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/addr_of_120_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/array_obj_ref_119_root_address_calculated
      -- CP-element group 24: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/array_obj_ref_119_offset_calculated
      -- CP-element group 24: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/array_obj_ref_119_final_index_sum_regn_Update/ack
      -- CP-element group 24: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/array_obj_ref_119_base_plus_offset/$entry
      -- CP-element group 24: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/array_obj_ref_119_base_plus_offset/$exit
      -- CP-element group 24: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/array_obj_ref_119_base_plus_offset/sum_rename_req
      -- CP-element group 24: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/array_obj_ref_119_base_plus_offset/sum_rename_ack
      -- CP-element group 24: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/addr_of_120_request/$entry
      -- CP-element group 24: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/addr_of_120_request/req
      -- 
    ack_350_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_119_index_offset_ack_1, ack => testConfigure_CP_0_elements(24)); -- 
    req_359_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_359_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(24), ack => addr_of_120_final_reg_req_0); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/addr_of_120_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/addr_of_120_request/$exit
      -- CP-element group 25: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/addr_of_120_request/ack
      -- 
    ack_360_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_120_final_reg_ack_0, ack => testConfigure_CP_0_elements(25)); -- 
    -- CP-element group 26:  fork  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	244 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	31 
    -- CP-element group 26: 	38 
    -- CP-element group 26:  members (35) 
      -- CP-element group 26: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/addr_of_120_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/addr_of_120_complete/$exit
      -- CP-element group 26: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/addr_of_120_complete/ack
      -- CP-element group 26: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_130_base_address_calculated
      -- CP-element group 26: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_130_word_address_calculated
      -- CP-element group 26: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_130_root_address_calculated
      -- CP-element group 26: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_130_base_address_resized
      -- CP-element group 26: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_130_base_addr_resize/$entry
      -- CP-element group 26: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_130_base_addr_resize/$exit
      -- CP-element group 26: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_130_base_addr_resize/base_resize_req
      -- CP-element group 26: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_130_base_addr_resize/base_resize_ack
      -- CP-element group 26: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_130_base_plus_offset/$entry
      -- CP-element group 26: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_130_base_plus_offset/$exit
      -- CP-element group 26: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_130_base_plus_offset/sum_rename_req
      -- CP-element group 26: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_130_base_plus_offset/sum_rename_ack
      -- CP-element group 26: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_130_word_addrgen/$entry
      -- CP-element group 26: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_130_word_addrgen/$exit
      -- CP-element group 26: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_130_word_addrgen/root_register_req
      -- CP-element group 26: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_130_word_addrgen/root_register_ack
      -- CP-element group 26: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_152_base_address_calculated
      -- CP-element group 26: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_152_word_address_calculated
      -- CP-element group 26: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_152_root_address_calculated
      -- CP-element group 26: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_152_base_address_resized
      -- CP-element group 26: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_152_base_addr_resize/$entry
      -- CP-element group 26: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_152_base_addr_resize/$exit
      -- CP-element group 26: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_152_base_addr_resize/base_resize_req
      -- CP-element group 26: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_152_base_addr_resize/base_resize_ack
      -- CP-element group 26: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_152_base_plus_offset/$entry
      -- CP-element group 26: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_152_base_plus_offset/$exit
      -- CP-element group 26: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_152_base_plus_offset/sum_rename_req
      -- CP-element group 26: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_152_base_plus_offset/sum_rename_ack
      -- CP-element group 26: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_152_word_addrgen/$entry
      -- CP-element group 26: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_152_word_addrgen/$exit
      -- CP-element group 26: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_152_word_addrgen/root_register_req
      -- CP-element group 26: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_152_word_addrgen/root_register_ack
      -- 
    ack_365_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_120_final_reg_ack_1, ack => testConfigure_CP_0_elements(26)); -- 
    -- CP-element group 27:  transition  input  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	244 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27:  members (6) 
      -- CP-element group 27: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/RPIPE_ConvTranspose_input_pipe_123_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/RPIPE_ConvTranspose_input_pipe_123_update_start_
      -- CP-element group 27: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/RPIPE_ConvTranspose_input_pipe_123_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/RPIPE_ConvTranspose_input_pipe_123_Sample/ra
      -- CP-element group 27: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/RPIPE_ConvTranspose_input_pipe_123_Update/$entry
      -- CP-element group 27: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/RPIPE_ConvTranspose_input_pipe_123_Update/cr
      -- 
    ra_374_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_123_inst_ack_0, ack => testConfigure_CP_0_elements(27)); -- 
    cr_378_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_378_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(27), ack => RPIPE_ConvTranspose_input_pipe_123_inst_req_1); -- 
    -- CP-element group 28:  fork  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28: 	34 
    -- CP-element group 28:  members (9) 
      -- CP-element group 28: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/RPIPE_ConvTranspose_input_pipe_123_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/RPIPE_ConvTranspose_input_pipe_123_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/RPIPE_ConvTranspose_input_pipe_123_Update/ca
      -- CP-element group 28: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/type_cast_127_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/type_cast_127_Sample/$entry
      -- CP-element group 28: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/type_cast_127_Sample/rr
      -- CP-element group 28: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/RPIPE_ConvTranspose_input_pipe_140_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/RPIPE_ConvTranspose_input_pipe_140_Sample/$entry
      -- CP-element group 28: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/RPIPE_ConvTranspose_input_pipe_140_Sample/rr
      -- 
    ca_379_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_123_inst_ack_1, ack => testConfigure_CP_0_elements(28)); -- 
    rr_387_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_387_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(28), ack => type_cast_127_inst_req_0); -- 
    rr_451_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_451_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(28), ack => RPIPE_ConvTranspose_input_pipe_140_inst_req_0); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/type_cast_127_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/type_cast_127_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/type_cast_127_Sample/ra
      -- 
    ra_388_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_127_inst_ack_0, ack => testConfigure_CP_0_elements(29)); -- 
    -- CP-element group 30:  fork  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	244 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30: 	38 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/type_cast_127_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/type_cast_127_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/type_cast_127_Update/ca
      -- 
    ca_393_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_127_inst_ack_1, ack => testConfigure_CP_0_elements(30)); -- 
    -- CP-element group 31:  join  transition  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: 	26 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (9) 
      -- CP-element group 31: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_130_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_130_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_130_Sample/ptr_deref_130_Split/$entry
      -- CP-element group 31: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_130_Sample/ptr_deref_130_Split/$exit
      -- CP-element group 31: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_130_Sample/ptr_deref_130_Split/split_req
      -- CP-element group 31: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_130_Sample/ptr_deref_130_Split/split_ack
      -- CP-element group 31: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_130_Sample/word_access_start/$entry
      -- CP-element group 31: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_130_Sample/word_access_start/word_0/$entry
      -- CP-element group 31: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_130_Sample/word_access_start/word_0/rr
      -- 
    rr_431_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_431_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(31), ack => ptr_deref_130_store_0_req_0); -- 
    testConfigure_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(30) & testConfigure_CP_0_elements(26);
      gj_testConfigure_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	41 
    -- CP-element group 32:  members (5) 
      -- CP-element group 32: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_130_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_130_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_130_Sample/word_access_start/$exit
      -- CP-element group 32: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_130_Sample/word_access_start/word_0/$exit
      -- CP-element group 32: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_130_Sample/word_access_start/word_0/ra
      -- 
    ra_432_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_130_store_0_ack_0, ack => testConfigure_CP_0_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	244 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	42 
    -- CP-element group 33:  members (5) 
      -- CP-element group 33: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_130_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_130_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_130_Update/word_access_complete/$exit
      -- CP-element group 33: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_130_Update/word_access_complete/word_0/$exit
      -- CP-element group 33: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_130_Update/word_access_complete/word_0/ca
      -- 
    ca_443_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_130_store_0_ack_1, ack => testConfigure_CP_0_elements(33)); -- 
    -- CP-element group 34:  transition  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	28 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34:  members (6) 
      -- CP-element group 34: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/RPIPE_ConvTranspose_input_pipe_140_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/RPIPE_ConvTranspose_input_pipe_140_update_start_
      -- CP-element group 34: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/RPIPE_ConvTranspose_input_pipe_140_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/RPIPE_ConvTranspose_input_pipe_140_Sample/ra
      -- CP-element group 34: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/RPIPE_ConvTranspose_input_pipe_140_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/RPIPE_ConvTranspose_input_pipe_140_Update/cr
      -- 
    ra_452_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_140_inst_ack_0, ack => testConfigure_CP_0_elements(34)); -- 
    cr_456_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_456_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(34), ack => RPIPE_ConvTranspose_input_pipe_140_inst_req_1); -- 
    -- CP-element group 35:  transition  input  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (6) 
      -- CP-element group 35: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/RPIPE_ConvTranspose_input_pipe_140_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/RPIPE_ConvTranspose_input_pipe_140_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/RPIPE_ConvTranspose_input_pipe_140_Update/ca
      -- CP-element group 35: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/type_cast_144_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/type_cast_144_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/type_cast_144_Sample/rr
      -- 
    ca_457_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_140_inst_ack_1, ack => testConfigure_CP_0_elements(35)); -- 
    rr_465_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_465_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(35), ack => type_cast_144_inst_req_0); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/type_cast_144_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/type_cast_144_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/type_cast_144_Sample/ra
      -- 
    ra_466_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_144_inst_ack_0, ack => testConfigure_CP_0_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	244 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/type_cast_144_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/type_cast_144_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/type_cast_144_Update/ca
      -- 
    ca_471_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_144_inst_ack_1, ack => testConfigure_CP_0_elements(37)); -- 
    -- CP-element group 38:  join  transition  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	30 
    -- CP-element group 38: 	37 
    -- CP-element group 38: 	41 
    -- CP-element group 38: 	26 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (9) 
      -- CP-element group 38: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_152_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_152_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_152_Sample/ptr_deref_152_Split/$entry
      -- CP-element group 38: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_152_Sample/ptr_deref_152_Split/$exit
      -- CP-element group 38: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_152_Sample/ptr_deref_152_Split/split_req
      -- CP-element group 38: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_152_Sample/ptr_deref_152_Split/split_ack
      -- CP-element group 38: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_152_Sample/word_access_start/$entry
      -- CP-element group 38: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_152_Sample/word_access_start/word_0/$entry
      -- CP-element group 38: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_152_Sample/word_access_start/word_0/rr
      -- 
    rr_509_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_509_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(38), ack => ptr_deref_152_store_0_req_0); -- 
    testConfigure_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(30) & testConfigure_CP_0_elements(37) & testConfigure_CP_0_elements(41) & testConfigure_CP_0_elements(26);
      gj_testConfigure_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (5) 
      -- CP-element group 39: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_152_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_152_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_152_Sample/word_access_start/$exit
      -- CP-element group 39: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_152_Sample/word_access_start/word_0/$exit
      -- CP-element group 39: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_152_Sample/word_access_start/word_0/ra
      -- 
    ra_510_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_152_store_0_ack_0, ack => testConfigure_CP_0_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	244 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	42 
    -- CP-element group 40:  members (5) 
      -- CP-element group 40: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_152_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_152_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_152_Update/word_access_complete/$exit
      -- CP-element group 40: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_152_Update/word_access_complete/word_0/$exit
      -- CP-element group 40: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_152_Update/word_access_complete/word_0/ca
      -- 
    ca_521_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_152_store_0_ack_1, ack => testConfigure_CP_0_elements(40)); -- 
    -- CP-element group 41:  transition  delay-element  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	32 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	38 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_130_ptr_deref_152_delay
      -- 
    -- Element group testConfigure_CP_0_elements(41) is a control-delay.
    cp_element_41_delay: control_delay_element  generic map(name => " 41_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(32), ack => testConfigure_CP_0_elements(41), clk => clk, reset =>reset);
    -- CP-element group 42:  branch  join  transition  place  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	33 
    -- CP-element group 42: 	40 
    -- CP-element group 42: 	23 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42: 	44 
    -- CP-element group 42:  members (10) 
      -- CP-element group 42: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166__exit__
      -- CP-element group 42: 	 branch_block_stmt_34/if_stmt_167__entry__
      -- CP-element group 42: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/$exit
      -- CP-element group 42: 	 branch_block_stmt_34/if_stmt_167_dead_link/$entry
      -- CP-element group 42: 	 branch_block_stmt_34/if_stmt_167_eval_test/$entry
      -- CP-element group 42: 	 branch_block_stmt_34/if_stmt_167_eval_test/$exit
      -- CP-element group 42: 	 branch_block_stmt_34/if_stmt_167_eval_test/branch_req
      -- CP-element group 42: 	 branch_block_stmt_34/R_exitcond4_168_place
      -- CP-element group 42: 	 branch_block_stmt_34/if_stmt_167_if_link/$entry
      -- CP-element group 42: 	 branch_block_stmt_34/if_stmt_167_else_link/$entry
      -- 
    branch_req_530_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_530_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(42), ack => if_stmt_167_branch_req_0); -- 
    testConfigure_cp_element_group_42: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_42"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(33) & testConfigure_CP_0_elements(40) & testConfigure_CP_0_elements(23);
      gj_testConfigure_cp_element_group_42 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(42), clk => clk, reset => reset); --
    end block;
    -- CP-element group 43:  merge  transition  place  input  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	45 
    -- CP-element group 43:  members (15) 
      -- CP-element group 43: 	 branch_block_stmt_34/merge_stmt_173__exit__
      -- CP-element group 43: 	 branch_block_stmt_34/assign_stmt_176__entry__
      -- CP-element group 43: 	 branch_block_stmt_34/if_stmt_167_if_link/$exit
      -- CP-element group 43: 	 branch_block_stmt_34/if_stmt_167_if_link/if_choice_transition
      -- CP-element group 43: 	 branch_block_stmt_34/forx_xbody16_bbx_xnph240
      -- CP-element group 43: 	 branch_block_stmt_34/assign_stmt_176/$entry
      -- CP-element group 43: 	 branch_block_stmt_34/assign_stmt_176/RPIPE_ConvTranspose_input_pipe_175_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_34/assign_stmt_176/RPIPE_ConvTranspose_input_pipe_175_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_34/assign_stmt_176/RPIPE_ConvTranspose_input_pipe_175_Sample/rr
      -- CP-element group 43: 	 branch_block_stmt_34/forx_xbody16_bbx_xnph240_PhiReq/$entry
      -- CP-element group 43: 	 branch_block_stmt_34/forx_xbody16_bbx_xnph240_PhiReq/$exit
      -- CP-element group 43: 	 branch_block_stmt_34/merge_stmt_173_PhiReqMerge
      -- CP-element group 43: 	 branch_block_stmt_34/merge_stmt_173_PhiAck/$entry
      -- CP-element group 43: 	 branch_block_stmt_34/merge_stmt_173_PhiAck/$exit
      -- CP-element group 43: 	 branch_block_stmt_34/merge_stmt_173_PhiAck/dummy
      -- 
    if_choice_transition_535_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_167_branch_ack_1, ack => testConfigure_CP_0_elements(43)); -- 
    rr_552_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_552_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(43), ack => RPIPE_ConvTranspose_input_pipe_175_inst_req_0); -- 
    -- CP-element group 44:  fork  transition  place  input  output  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	42 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	239 
    -- CP-element group 44: 	240 
    -- CP-element group 44:  members (12) 
      -- CP-element group 44: 	 branch_block_stmt_34/if_stmt_167_else_link/$exit
      -- CP-element group 44: 	 branch_block_stmt_34/if_stmt_167_else_link/else_choice_transition
      -- CP-element group 44: 	 branch_block_stmt_34/forx_xbody16_forx_xbody16
      -- CP-element group 44: 	 branch_block_stmt_34/forx_xbody16_forx_xbody16_PhiReq/$entry
      -- CP-element group 44: 	 branch_block_stmt_34/forx_xbody16_forx_xbody16_PhiReq/phi_stmt_107/$entry
      -- CP-element group 44: 	 branch_block_stmt_34/forx_xbody16_forx_xbody16_PhiReq/phi_stmt_107/phi_stmt_107_sources/$entry
      -- CP-element group 44: 	 branch_block_stmt_34/forx_xbody16_forx_xbody16_PhiReq/phi_stmt_107/phi_stmt_107_sources/type_cast_110/$entry
      -- CP-element group 44: 	 branch_block_stmt_34/forx_xbody16_forx_xbody16_PhiReq/phi_stmt_107/phi_stmt_107_sources/type_cast_110/SplitProtocol/$entry
      -- CP-element group 44: 	 branch_block_stmt_34/forx_xbody16_forx_xbody16_PhiReq/phi_stmt_107/phi_stmt_107_sources/type_cast_110/SplitProtocol/Sample/$entry
      -- CP-element group 44: 	 branch_block_stmt_34/forx_xbody16_forx_xbody16_PhiReq/phi_stmt_107/phi_stmt_107_sources/type_cast_110/SplitProtocol/Sample/rr
      -- CP-element group 44: 	 branch_block_stmt_34/forx_xbody16_forx_xbody16_PhiReq/phi_stmt_107/phi_stmt_107_sources/type_cast_110/SplitProtocol/Update/$entry
      -- CP-element group 44: 	 branch_block_stmt_34/forx_xbody16_forx_xbody16_PhiReq/phi_stmt_107/phi_stmt_107_sources/type_cast_110/SplitProtocol/Update/cr
      -- 
    else_choice_transition_539_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_167_branch_ack_0, ack => testConfigure_CP_0_elements(44)); -- 
    rr_2684_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2684_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(44), ack => type_cast_110_inst_req_0); -- 
    cr_2689_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2689_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(44), ack => type_cast_110_inst_req_1); -- 
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	43 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (6) 
      -- CP-element group 45: 	 branch_block_stmt_34/assign_stmt_176/RPIPE_ConvTranspose_input_pipe_175_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_34/assign_stmt_176/RPIPE_ConvTranspose_input_pipe_175_update_start_
      -- CP-element group 45: 	 branch_block_stmt_34/assign_stmt_176/RPIPE_ConvTranspose_input_pipe_175_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_34/assign_stmt_176/RPIPE_ConvTranspose_input_pipe_175_Sample/ra
      -- CP-element group 45: 	 branch_block_stmt_34/assign_stmt_176/RPIPE_ConvTranspose_input_pipe_175_Update/$entry
      -- CP-element group 45: 	 branch_block_stmt_34/assign_stmt_176/RPIPE_ConvTranspose_input_pipe_175_Update/cr
      -- 
    ra_553_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_175_inst_ack_0, ack => testConfigure_CP_0_elements(45)); -- 
    cr_557_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_557_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(45), ack => RPIPE_ConvTranspose_input_pipe_175_inst_req_1); -- 
    -- CP-element group 46:  fork  transition  place  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	245 
    -- CP-element group 46: 	246 
    -- CP-element group 46: 	247 
    -- CP-element group 46:  members (17) 
      -- CP-element group 46: 	 branch_block_stmt_34/assign_stmt_176__exit__
      -- CP-element group 46: 	 branch_block_stmt_34/bbx_xnph240_forx_xbody41
      -- CP-element group 46: 	 branch_block_stmt_34/assign_stmt_176/$exit
      -- CP-element group 46: 	 branch_block_stmt_34/assign_stmt_176/RPIPE_ConvTranspose_input_pipe_175_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_34/assign_stmt_176/RPIPE_ConvTranspose_input_pipe_175_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_34/assign_stmt_176/RPIPE_ConvTranspose_input_pipe_175_Update/ca
      -- CP-element group 46: 	 branch_block_stmt_34/bbx_xnph240_forx_xbody41_PhiReq/$entry
      -- CP-element group 46: 	 branch_block_stmt_34/bbx_xnph240_forx_xbody41_PhiReq/phi_stmt_179/$entry
      -- CP-element group 46: 	 branch_block_stmt_34/bbx_xnph240_forx_xbody41_PhiReq/phi_stmt_179/phi_stmt_179_sources/$entry
      -- CP-element group 46: 	 branch_block_stmt_34/bbx_xnph240_forx_xbody41_PhiReq/phi_stmt_186/$entry
      -- CP-element group 46: 	 branch_block_stmt_34/bbx_xnph240_forx_xbody41_PhiReq/phi_stmt_186/phi_stmt_186_sources/$entry
      -- CP-element group 46: 	 branch_block_stmt_34/bbx_xnph240_forx_xbody41_PhiReq/phi_stmt_186/phi_stmt_186_sources/type_cast_189/$entry
      -- CP-element group 46: 	 branch_block_stmt_34/bbx_xnph240_forx_xbody41_PhiReq/phi_stmt_186/phi_stmt_186_sources/type_cast_189/SplitProtocol/$entry
      -- CP-element group 46: 	 branch_block_stmt_34/bbx_xnph240_forx_xbody41_PhiReq/phi_stmt_186/phi_stmt_186_sources/type_cast_189/SplitProtocol/Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_34/bbx_xnph240_forx_xbody41_PhiReq/phi_stmt_186/phi_stmt_186_sources/type_cast_189/SplitProtocol/Sample/rr
      -- CP-element group 46: 	 branch_block_stmt_34/bbx_xnph240_forx_xbody41_PhiReq/phi_stmt_186/phi_stmt_186_sources/type_cast_189/SplitProtocol/Update/$entry
      -- CP-element group 46: 	 branch_block_stmt_34/bbx_xnph240_forx_xbody41_PhiReq/phi_stmt_186/phi_stmt_186_sources/type_cast_189/SplitProtocol/Update/cr
      -- 
    ca_558_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_175_inst_ack_1, ack => testConfigure_CP_0_elements(46)); -- 
    rr_2746_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2746_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(46), ack => type_cast_189_inst_req_0); -- 
    cr_2751_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2751_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(46), ack => type_cast_189_inst_req_1); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	260 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/addr_of_196_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/addr_of_196_request/$exit
      -- CP-element group 47: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/addr_of_196_request/ack
      -- 
    ack_595_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_196_final_reg_ack_0, ack => testConfigure_CP_0_elements(47)); -- 
    -- CP-element group 48:  join  fork  transition  input  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	260 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (28) 
      -- CP-element group 48: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/addr_of_196_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/addr_of_196_complete/$exit
      -- CP-element group 48: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/addr_of_196_complete/ack
      -- CP-element group 48: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/ptr_deref_199_sample_start_
      -- CP-element group 48: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/ptr_deref_199_base_address_calculated
      -- CP-element group 48: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/ptr_deref_199_word_address_calculated
      -- CP-element group 48: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/ptr_deref_199_root_address_calculated
      -- CP-element group 48: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/ptr_deref_199_base_address_resized
      -- CP-element group 48: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/ptr_deref_199_base_addr_resize/$entry
      -- CP-element group 48: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/ptr_deref_199_base_addr_resize/$exit
      -- CP-element group 48: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/ptr_deref_199_base_addr_resize/base_resize_req
      -- CP-element group 48: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/ptr_deref_199_base_addr_resize/base_resize_ack
      -- CP-element group 48: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/ptr_deref_199_base_plus_offset/$entry
      -- CP-element group 48: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/ptr_deref_199_base_plus_offset/$exit
      -- CP-element group 48: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/ptr_deref_199_base_plus_offset/sum_rename_req
      -- CP-element group 48: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/ptr_deref_199_base_plus_offset/sum_rename_ack
      -- CP-element group 48: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/ptr_deref_199_word_addrgen/$entry
      -- CP-element group 48: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/ptr_deref_199_word_addrgen/$exit
      -- CP-element group 48: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/ptr_deref_199_word_addrgen/root_register_req
      -- CP-element group 48: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/ptr_deref_199_word_addrgen/root_register_ack
      -- CP-element group 48: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/ptr_deref_199_Sample/$entry
      -- CP-element group 48: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/ptr_deref_199_Sample/ptr_deref_199_Split/$entry
      -- CP-element group 48: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/ptr_deref_199_Sample/ptr_deref_199_Split/$exit
      -- CP-element group 48: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/ptr_deref_199_Sample/ptr_deref_199_Split/split_req
      -- CP-element group 48: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/ptr_deref_199_Sample/ptr_deref_199_Split/split_ack
      -- CP-element group 48: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/ptr_deref_199_Sample/word_access_start/$entry
      -- CP-element group 48: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/ptr_deref_199_Sample/word_access_start/word_0/$entry
      -- CP-element group 48: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/ptr_deref_199_Sample/word_access_start/word_0/rr
      -- 
    ack_600_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_196_final_reg_ack_1, ack => testConfigure_CP_0_elements(48)); -- 
    rr_638_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_638_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(48), ack => ptr_deref_199_store_0_req_0); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (5) 
      -- CP-element group 49: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/ptr_deref_199_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/ptr_deref_199_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/ptr_deref_199_Sample/word_access_start/$exit
      -- CP-element group 49: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/ptr_deref_199_Sample/word_access_start/word_0/$exit
      -- CP-element group 49: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/ptr_deref_199_Sample/word_access_start/word_0/ra
      -- 
    ra_639_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_199_store_0_ack_0, ack => testConfigure_CP_0_elements(49)); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	260 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	53 
    -- CP-element group 50:  members (5) 
      -- CP-element group 50: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/ptr_deref_199_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/ptr_deref_199_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/ptr_deref_199_Update/word_access_complete/$exit
      -- CP-element group 50: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/ptr_deref_199_Update/word_access_complete/word_0/$exit
      -- CP-element group 50: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/ptr_deref_199_Update/word_access_complete/word_0/ca
      -- 
    ca_650_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_199_store_0_ack_1, ack => testConfigure_CP_0_elements(50)); -- 
    -- CP-element group 51:  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	260 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (6) 
      -- CP-element group 51: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/RPIPE_ConvTranspose_input_pipe_203_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/RPIPE_ConvTranspose_input_pipe_203_update_start_
      -- CP-element group 51: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/RPIPE_ConvTranspose_input_pipe_203_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/RPIPE_ConvTranspose_input_pipe_203_Sample/ra
      -- CP-element group 51: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/RPIPE_ConvTranspose_input_pipe_203_Update/$entry
      -- CP-element group 51: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/RPIPE_ConvTranspose_input_pipe_203_Update/cr
      -- 
    ra_659_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_203_inst_ack_0, ack => testConfigure_CP_0_elements(51)); -- 
    cr_663_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_663_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(51), ack => RPIPE_ConvTranspose_input_pipe_203_inst_req_1); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	53 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/RPIPE_ConvTranspose_input_pipe_203_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/RPIPE_ConvTranspose_input_pipe_203_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/RPIPE_ConvTranspose_input_pipe_203_Update/ca
      -- 
    ca_664_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_203_inst_ack_1, ack => testConfigure_CP_0_elements(52)); -- 
    -- CP-element group 53:  branch  join  transition  place  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	52 
    -- CP-element group 53: 	50 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (10) 
      -- CP-element group 53: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216__exit__
      -- CP-element group 53: 	 branch_block_stmt_34/if_stmt_217__entry__
      -- CP-element group 53: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/$exit
      -- CP-element group 53: 	 branch_block_stmt_34/if_stmt_217_dead_link/$entry
      -- CP-element group 53: 	 branch_block_stmt_34/if_stmt_217_eval_test/$entry
      -- CP-element group 53: 	 branch_block_stmt_34/if_stmt_217_eval_test/$exit
      -- CP-element group 53: 	 branch_block_stmt_34/if_stmt_217_eval_test/branch_req
      -- CP-element group 53: 	 branch_block_stmt_34/R_exitcond3_218_place
      -- CP-element group 53: 	 branch_block_stmt_34/if_stmt_217_if_link/$entry
      -- CP-element group 53: 	 branch_block_stmt_34/if_stmt_217_else_link/$entry
      -- 
    branch_req_672_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_672_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(53), ack => if_stmt_217_branch_req_0); -- 
    testConfigure_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(52) & testConfigure_CP_0_elements(50);
      gj_testConfigure_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  fork  transition  place  input  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	261 
    -- CP-element group 54: 	262 
    -- CP-element group 54:  members (12) 
      -- CP-element group 54: 	 branch_block_stmt_34/if_stmt_217_if_link/$exit
      -- CP-element group 54: 	 branch_block_stmt_34/if_stmt_217_if_link/if_choice_transition
      -- CP-element group 54: 	 branch_block_stmt_34/forx_xbody41_forx_xend49
      -- CP-element group 54: 	 branch_block_stmt_34/forx_xbody41_forx_xend49_PhiReq/$entry
      -- CP-element group 54: 	 branch_block_stmt_34/forx_xbody41_forx_xend49_PhiReq/phi_stmt_224/$entry
      -- CP-element group 54: 	 branch_block_stmt_34/forx_xbody41_forx_xend49_PhiReq/phi_stmt_224/phi_stmt_224_sources/$entry
      -- CP-element group 54: 	 branch_block_stmt_34/forx_xbody41_forx_xend49_PhiReq/phi_stmt_224/phi_stmt_224_sources/type_cast_227/$entry
      -- CP-element group 54: 	 branch_block_stmt_34/forx_xbody41_forx_xend49_PhiReq/phi_stmt_224/phi_stmt_224_sources/type_cast_227/SplitProtocol/$entry
      -- CP-element group 54: 	 branch_block_stmt_34/forx_xbody41_forx_xend49_PhiReq/phi_stmt_224/phi_stmt_224_sources/type_cast_227/SplitProtocol/Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_34/forx_xbody41_forx_xend49_PhiReq/phi_stmt_224/phi_stmt_224_sources/type_cast_227/SplitProtocol/Sample/rr
      -- CP-element group 54: 	 branch_block_stmt_34/forx_xbody41_forx_xend49_PhiReq/phi_stmt_224/phi_stmt_224_sources/type_cast_227/SplitProtocol/Update/$entry
      -- CP-element group 54: 	 branch_block_stmt_34/forx_xbody41_forx_xend49_PhiReq/phi_stmt_224/phi_stmt_224_sources/type_cast_227/SplitProtocol/Update/cr
      -- 
    if_choice_transition_677_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_217_branch_ack_1, ack => testConfigure_CP_0_elements(54)); -- 
    rr_2831_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2831_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(54), ack => type_cast_227_inst_req_0); -- 
    cr_2836_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2836_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(54), ack => type_cast_227_inst_req_1); -- 
    -- CP-element group 55:  fork  transition  place  input  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	250 
    -- CP-element group 55: 	251 
    -- CP-element group 55: 	253 
    -- CP-element group 55: 	254 
    -- CP-element group 55:  members (20) 
      -- CP-element group 55: 	 branch_block_stmt_34/if_stmt_217_else_link/$exit
      -- CP-element group 55: 	 branch_block_stmt_34/if_stmt_217_else_link/else_choice_transition
      -- CP-element group 55: 	 branch_block_stmt_34/forx_xbody41_forx_xbody41
      -- CP-element group 55: 	 branch_block_stmt_34/forx_xbody41_forx_xbody41_PhiReq/$entry
      -- CP-element group 55: 	 branch_block_stmt_34/forx_xbody41_forx_xbody41_PhiReq/phi_stmt_179/$entry
      -- CP-element group 55: 	 branch_block_stmt_34/forx_xbody41_forx_xbody41_PhiReq/phi_stmt_179/phi_stmt_179_sources/$entry
      -- CP-element group 55: 	 branch_block_stmt_34/forx_xbody41_forx_xbody41_PhiReq/phi_stmt_179/phi_stmt_179_sources/type_cast_185/$entry
      -- CP-element group 55: 	 branch_block_stmt_34/forx_xbody41_forx_xbody41_PhiReq/phi_stmt_179/phi_stmt_179_sources/type_cast_185/SplitProtocol/$entry
      -- CP-element group 55: 	 branch_block_stmt_34/forx_xbody41_forx_xbody41_PhiReq/phi_stmt_179/phi_stmt_179_sources/type_cast_185/SplitProtocol/Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_34/forx_xbody41_forx_xbody41_PhiReq/phi_stmt_179/phi_stmt_179_sources/type_cast_185/SplitProtocol/Sample/rr
      -- CP-element group 55: 	 branch_block_stmt_34/forx_xbody41_forx_xbody41_PhiReq/phi_stmt_179/phi_stmt_179_sources/type_cast_185/SplitProtocol/Update/$entry
      -- CP-element group 55: 	 branch_block_stmt_34/forx_xbody41_forx_xbody41_PhiReq/phi_stmt_179/phi_stmt_179_sources/type_cast_185/SplitProtocol/Update/cr
      -- CP-element group 55: 	 branch_block_stmt_34/forx_xbody41_forx_xbody41_PhiReq/phi_stmt_186/$entry
      -- CP-element group 55: 	 branch_block_stmt_34/forx_xbody41_forx_xbody41_PhiReq/phi_stmt_186/phi_stmt_186_sources/$entry
      -- CP-element group 55: 	 branch_block_stmt_34/forx_xbody41_forx_xbody41_PhiReq/phi_stmt_186/phi_stmt_186_sources/type_cast_191/$entry
      -- CP-element group 55: 	 branch_block_stmt_34/forx_xbody41_forx_xbody41_PhiReq/phi_stmt_186/phi_stmt_186_sources/type_cast_191/SplitProtocol/$entry
      -- CP-element group 55: 	 branch_block_stmt_34/forx_xbody41_forx_xbody41_PhiReq/phi_stmt_186/phi_stmt_186_sources/type_cast_191/SplitProtocol/Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_34/forx_xbody41_forx_xbody41_PhiReq/phi_stmt_186/phi_stmt_186_sources/type_cast_191/SplitProtocol/Sample/rr
      -- CP-element group 55: 	 branch_block_stmt_34/forx_xbody41_forx_xbody41_PhiReq/phi_stmt_186/phi_stmt_186_sources/type_cast_191/SplitProtocol/Update/$entry
      -- CP-element group 55: 	 branch_block_stmt_34/forx_xbody41_forx_xbody41_PhiReq/phi_stmt_186/phi_stmt_186_sources/type_cast_191/SplitProtocol/Update/cr
      -- 
    else_choice_transition_681_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_217_branch_ack_0, ack => testConfigure_CP_0_elements(55)); -- 
    rr_2772_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2772_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(55), ack => type_cast_185_inst_req_0); -- 
    cr_2777_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2777_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(55), ack => type_cast_185_inst_req_1); -- 
    rr_2795_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2795_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(55), ack => type_cast_191_inst_req_0); -- 
    cr_2800_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2800_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(55), ack => type_cast_191_inst_req_1); -- 
    -- CP-element group 56:  join  fork  transition  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	264 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56: 	58 
    -- CP-element group 56: 	59 
    -- CP-element group 56: 	62 
    -- CP-element group 56: 	63 
    -- CP-element group 56: 	65 
    -- CP-element group 56: 	69 
    -- CP-element group 56: 	70 
    -- CP-element group 56: 	72 
    -- CP-element group 56: 	76 
    -- CP-element group 56: 	77 
    -- CP-element group 56: 	79 
    -- CP-element group 56: 	83 
    -- CP-element group 56: 	84 
    -- CP-element group 56: 	86 
    -- CP-element group 56: 	90 
    -- CP-element group 56: 	91 
    -- CP-element group 56: 	93 
    -- CP-element group 56: 	97 
    -- CP-element group 56: 	98 
    -- CP-element group 56: 	100 
    -- CP-element group 56: 	101 
    -- CP-element group 56: 	102 
    -- CP-element group 56: 	103 
    -- CP-element group 56: 	104 
    -- CP-element group 56: 	105 
    -- CP-element group 56: 	106 
    -- CP-element group 56: 	107 
    -- CP-element group 56: 	108 
    -- CP-element group 56: 	109 
    -- CP-element group 56: 	110 
    -- CP-element group 56: 	111 
    -- CP-element group 56: 	112 
    -- CP-element group 56: 	113 
    -- CP-element group 56: 	114 
    -- CP-element group 56:  members (346) 
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_471_base_plus_offset/sum_rename_req
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_471_word_addrgen/$exit
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_471_base_addr_resize/base_resize_ack
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_471_base_addr_resize/base_resize_req
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_471_word_addrgen/root_register_ack
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_471_word_addrgen/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_471_base_addr_resize/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_471_base_addr_resize/$exit
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_389_base_plus_offset/$exit
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_435_word_addrgen/root_register_ack
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_401_base_addr_resize/base_resize_req
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_401_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_471_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_401_base_addr_resize/$exit
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_401_base_addr_resize/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_471_Update/word_access_complete/word_0/cr
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_459_base_addr_resize/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_471_base_plus_offset/sum_rename_ack
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_447_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_447_base_addr_resize/base_resize_ack
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_413_base_plus_offset/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_389_base_plus_offset/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_360_update_start_
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_435_word_addrgen/root_register_req
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_389_base_addr_resize/base_resize_ack
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_389_base_addr_resize/base_resize_req
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_389_base_addr_resize/$exit
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_459_base_addr_resize/base_resize_req
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_435_Sample/word_access_start/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_435_word_addrgen/$exit
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_401_base_address_resized
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_435_word_addrgen/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_459_base_addr_resize/$exit
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_459_Update/word_access_complete/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_401_word_addrgen/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_376_base_plus_offset/sum_rename_req
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_413_update_start_
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_401_root_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_376_word_addrgen/root_register_ack
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_447_Sample/word_access_start/word_0/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_376_word_addrgen/root_register_req
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_435_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_413_base_addr_resize/base_resize_ack
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_376_word_addrgen/$exit
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_459_base_address_resized
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_471_base_address_resized
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_459_Sample/word_access_start/word_0/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_447_base_addr_resize/base_resize_req
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_459_Update/word_access_complete/word_0/cr
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_401_word_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_413_base_addr_resize/base_resize_req
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_471_Update/word_access_complete/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_459_root_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_413_base_addr_resize/$exit
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_413_base_addr_resize/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_401_base_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_389_base_addr_resize/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_413_base_address_resized
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_389_base_address_resized
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_459_word_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_389_root_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_459_base_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_447_Sample/word_access_start/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_447_base_addr_resize/$exit
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_435_base_plus_offset/sum_rename_ack
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_435_base_plus_offset/sum_rename_req
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_413_root_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_376_word_addrgen/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_459_Sample/word_access_start/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_459_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_459_Update/word_access_complete/word_0/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_413_word_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_447_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_471_Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_401_update_start_
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_459_update_start_
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_413_base_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_389_word_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_389_base_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_401_word_addrgen/root_register_ack
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_376_base_plus_offset/sum_rename_ack
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_401_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_471_word_addrgen/root_register_req
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_435_base_plus_offset/$exit
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_447_base_addr_resize/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_401_word_addrgen/root_register_req
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_471_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_346_word_addrgen/root_register_ack
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_389_update_start_
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_459_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_435_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_435_base_plus_offset/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_413_Update/word_access_complete/word_0/cr
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_346_Update/word_access_complete/word_0/cr
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_401_word_addrgen/$exit
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_401_Sample/word_access_start/word_0/rr
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_346_base_plus_offset/sum_rename_req
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_248_Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_248_Update/word_access_complete/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_248_Update/word_access_complete/word_0/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_248_Update/word_access_complete/word_0/cr
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_413_base_plus_offset/sum_rename_req
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_346_base_plus_offset/$exit
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_360_Update/cr
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_435_update_start_
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_376_base_plus_offset/$exit
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_447_base_address_resized
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_471_Sample/word_access_start/word_0/rr
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_376_base_plus_offset/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_413_Update/word_access_complete/word_0/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_413_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_376_base_addr_resize/base_resize_ack
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_471_root_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_459_word_addrgen/root_register_ack
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_459_word_addrgen/root_register_req
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_447_root_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_447_word_addrgen/root_register_ack
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_413_Update/word_access_complete/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_413_Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_376_Update/word_access_complete/word_0/cr
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_389_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_447_word_addrgen/root_register_req
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_471_Sample/word_access_start/word_0/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_435_base_addr_resize/base_resize_ack
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_435_base_addr_resize/base_resize_req
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_376_base_addr_resize/base_resize_req
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_471_word_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_459_word_addrgen/$exit
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_447_word_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_459_Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_346_word_addrgen/root_register_req
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_447_word_addrgen/$exit
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_447_word_addrgen/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_413_Sample/word_access_start/word_0/rr
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_413_Sample/word_access_start/word_0/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_413_Sample/word_access_start/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_413_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_435_Update/word_access_complete/word_0/cr
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_376_Update/word_access_complete/word_0/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_346_Update/word_access_complete/word_0/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_459_word_addrgen/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_471_Sample/word_access_start/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_447_base_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_435_base_addr_resize/$exit
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_346_Update/word_access_complete/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_401_base_plus_offset/sum_rename_ack
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_346_Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_376_Update/word_access_complete/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_401_base_plus_offset/sum_rename_req
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_435_Update/word_access_complete/word_0/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_435_base_addr_resize/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_376_base_addr_resize/$exit
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_471_base_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_401_base_plus_offset/$exit
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_447_Update/word_access_complete/word_0/cr
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_413_word_addrgen/root_register_ack
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_401_base_plus_offset/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_389_Update/word_access_complete/word_0/cr
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_447_Update/word_access_complete/word_0/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_376_base_addr_resize/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_471_base_plus_offset/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_471_base_plus_offset/$exit
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_435_Update/word_access_complete/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_447_base_plus_offset/sum_rename_ack
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_413_word_addrgen/root_register_req
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_413_word_addrgen/$exit
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_413_word_addrgen/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_401_Update/word_access_complete/word_0/cr
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_435_base_address_resized
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_401_Update/word_access_complete/word_0/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_376_Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_447_Update/word_access_complete/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_389_Update/word_access_complete/word_0/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_459_base_plus_offset/sum_rename_ack
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_447_base_plus_offset/sum_rename_req
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_471_Update/word_access_complete/word_0/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_346_word_addrgen/$exit
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_435_root_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_447_Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_459_base_plus_offset/sum_rename_req
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_459_base_plus_offset/$exit
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_459_base_plus_offset/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_389_Update/word_access_complete/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_435_word_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_435_Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_401_base_addr_resize/base_resize_ack
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_346_word_addrgen/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/STORE_padding_229_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/STORE_padding_229_update_start_
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_447_base_plus_offset/$exit
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/STORE_padding_229_word_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/STORE_padding_229_root_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_447_base_plus_offset/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/STORE_padding_229_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/STORE_padding_229_Sample/STORE_padding_229_Split/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/STORE_padding_229_Sample/STORE_padding_229_Split/$exit
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/STORE_padding_229_Sample/STORE_padding_229_Split/split_req
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_401_Update/word_access_complete/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/STORE_padding_229_Sample/STORE_padding_229_Split/split_ack
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/STORE_padding_229_Sample/word_access_start/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/STORE_padding_229_Sample/word_access_start/word_0/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/STORE_padding_229_Sample/word_access_start/word_0/rr
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_376_base_address_resized
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/STORE_padding_229_Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/STORE_padding_229_Update/word_access_complete/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/STORE_padding_229_Update/word_access_complete/word_0/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/STORE_padding_229_Update/word_access_complete/word_0/cr
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_389_Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_447_update_start_
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_233_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_435_base_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_233_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_233_Sample/rr
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_376_root_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_237_update_start_
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_389_Sample/word_access_start/word_0/rr
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_401_Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_237_Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_435_Sample/word_access_start/word_0/rr
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_237_Update/cr
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_376_word_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_413_base_plus_offset/sum_rename_ack
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_376_base_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_389_Sample/word_access_start/word_0/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_248_update_start_
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_248_base_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_389_Sample/word_access_start/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_248_word_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_248_root_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_248_base_address_resized
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_248_base_addr_resize/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_248_base_addr_resize/$exit
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_447_Sample/word_access_start/word_0/rr
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_248_base_addr_resize/base_resize_req
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_248_base_addr_resize/base_resize_ack
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_389_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_248_base_plus_offset/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_248_base_plus_offset/$exit
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_248_base_plus_offset/sum_rename_req
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_248_base_plus_offset/sum_rename_ack
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_376_update_start_
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_248_word_addrgen/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_248_word_addrgen/$exit
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_248_word_addrgen/root_register_req
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_248_word_addrgen/root_register_ack
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_346_base_plus_offset/sum_rename_ack
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_401_Sample/word_access_start/word_0/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_471_update_start_
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_459_base_addr_resize/base_resize_ack
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_389_word_addrgen/root_register_ack
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_262_update_start_
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_389_word_addrgen/root_register_req
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_262_Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_262_Update/cr
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_360_Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_413_base_plus_offset/$exit
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_389_word_addrgen/$exit
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_278_update_start_
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_389_word_addrgen/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_278_base_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_278_word_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_278_root_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_278_base_address_resized
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_278_base_addr_resize/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_278_base_addr_resize/$exit
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_278_base_addr_resize/base_resize_req
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_401_Sample/word_access_start/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_278_base_addr_resize/base_resize_ack
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_389_base_plus_offset/sum_rename_ack
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_278_base_plus_offset/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_278_base_plus_offset/$exit
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_278_base_plus_offset/sum_rename_req
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_278_base_plus_offset/sum_rename_ack
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_278_word_addrgen/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_278_word_addrgen/$exit
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_459_Sample/word_access_start/word_0/rr
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_278_word_addrgen/root_register_req
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_278_word_addrgen/root_register_ack
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_346_base_plus_offset/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_389_base_plus_offset/sum_rename_req
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_435_Sample/word_access_start/word_0/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_278_Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_278_Update/word_access_complete/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_278_Update/word_access_complete/word_0/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_278_Update/word_access_complete/word_0/cr
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_286_update_start_
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_286_Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_286_Update/cr
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_297_update_start_
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_297_base_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_297_word_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_297_root_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_297_base_address_resized
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_297_base_addr_resize/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_297_base_addr_resize/$exit
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_297_base_addr_resize/base_resize_req
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_297_base_addr_resize/base_resize_ack
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_297_base_plus_offset/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_297_base_plus_offset/$exit
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_297_base_plus_offset/sum_rename_req
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_297_base_plus_offset/sum_rename_ack
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_297_word_addrgen/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_297_word_addrgen/$exit
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_297_word_addrgen/root_register_req
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_297_word_addrgen/root_register_ack
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_297_Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_297_Update/word_access_complete/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_297_Update/word_access_complete/word_0/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_297_Update/word_access_complete/word_0/cr
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_311_update_start_
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_311_Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_311_Update/cr
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_327_update_start_
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_327_base_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_327_word_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_327_root_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_327_base_address_resized
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_327_base_addr_resize/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_327_base_addr_resize/$exit
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_327_base_addr_resize/base_resize_req
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_327_base_addr_resize/base_resize_ack
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_327_base_plus_offset/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_327_base_plus_offset/$exit
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_327_base_plus_offset/sum_rename_req
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_327_base_plus_offset/sum_rename_ack
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_327_word_addrgen/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_327_word_addrgen/$exit
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_327_word_addrgen/root_register_req
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_327_word_addrgen/root_register_ack
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_327_Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_327_Update/word_access_complete/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_327_Update/word_access_complete/word_0/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_327_Update/word_access_complete/word_0/cr
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_335_update_start_
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_335_Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_335_Update/cr
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_346_update_start_
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_346_base_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_346_word_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_346_root_address_calculated
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_346_base_address_resized
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_346_base_addr_resize/$entry
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_346_base_addr_resize/$exit
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_346_base_addr_resize/base_resize_req
      -- CP-element group 56: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_346_base_addr_resize/base_resize_ack
      -- 
    cr_718_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_718_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(56), ack => STORE_padding_229_store_0_req_1); -- 
    rr_707_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_707_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(56), ack => STORE_padding_229_store_0_req_0); -- 
    rr_727_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_727_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(56), ack => RPIPE_ConvTranspose_input_pipe_233_inst_req_0); -- 
    cr_746_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_746_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(56), ack => type_cast_237_inst_req_1); -- 
    cr_796_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_796_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(56), ack => ptr_deref_248_store_0_req_1); -- 
    cr_824_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_824_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(56), ack => type_cast_262_inst_req_1); -- 
    cr_874_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_874_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(56), ack => ptr_deref_278_store_0_req_1); -- 
    cr_902_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_902_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(56), ack => type_cast_286_inst_req_1); -- 
    cr_952_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_952_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(56), ack => ptr_deref_297_store_0_req_1); -- 
    cr_980_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_980_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(56), ack => type_cast_311_inst_req_1); -- 
    cr_1030_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1030_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(56), ack => ptr_deref_327_store_0_req_1); -- 
    cr_1058_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1058_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(56), ack => type_cast_335_inst_req_1); -- 
    cr_1108_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1108_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(56), ack => ptr_deref_346_store_0_req_1); -- 
    cr_1136_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1136_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(56), ack => type_cast_360_inst_req_1); -- 
    cr_1186_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1186_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(56), ack => ptr_deref_376_store_0_req_1); -- 
    cr_1231_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1231_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(56), ack => ptr_deref_389_load_0_req_1); -- 
    rr_1220_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1220_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(56), ack => ptr_deref_389_load_0_req_0); -- 
    cr_1281_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1281_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(56), ack => ptr_deref_401_load_0_req_1); -- 
    rr_1270_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1270_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(56), ack => ptr_deref_401_load_0_req_0); -- 
    cr_1331_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1331_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(56), ack => ptr_deref_413_load_0_req_1); -- 
    rr_1320_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1320_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(56), ack => ptr_deref_413_load_0_req_0); -- 
    cr_1381_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1381_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(56), ack => ptr_deref_435_load_0_req_1); -- 
    rr_1370_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1370_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(56), ack => ptr_deref_435_load_0_req_0); -- 
    cr_1431_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1431_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(56), ack => ptr_deref_447_load_0_req_1); -- 
    rr_1420_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1420_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(56), ack => ptr_deref_447_load_0_req_0); -- 
    cr_1481_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1481_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(56), ack => ptr_deref_459_load_0_req_1); -- 
    rr_1470_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1470_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(56), ack => ptr_deref_459_load_0_req_0); -- 
    cr_1531_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1531_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(56), ack => ptr_deref_471_load_0_req_1); -- 
    rr_1520_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1520_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(56), ack => ptr_deref_471_load_0_req_0); -- 
    testConfigure_CP_0_elements(56) <= testConfigure_CP_0_elements(264);
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (5) 
      -- CP-element group 57: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/STORE_padding_229_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/STORE_padding_229_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/STORE_padding_229_Sample/word_access_start/$exit
      -- CP-element group 57: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/STORE_padding_229_Sample/word_access_start/word_0/$exit
      -- CP-element group 57: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/STORE_padding_229_Sample/word_access_start/word_0/ra
      -- 
    ra_708_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_padding_229_store_0_ack_0, ack => testConfigure_CP_0_elements(57)); -- 
    -- CP-element group 58:  transition  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	56 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	120 
    -- CP-element group 58:  members (5) 
      -- CP-element group 58: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/STORE_padding_229_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/STORE_padding_229_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/STORE_padding_229_Update/word_access_complete/$exit
      -- CP-element group 58: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/STORE_padding_229_Update/word_access_complete/word_0/$exit
      -- CP-element group 58: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/STORE_padding_229_Update/word_access_complete/word_0/ca
      -- 
    ca_719_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_padding_229_store_0_ack_1, ack => testConfigure_CP_0_elements(58)); -- 
    -- CP-element group 59:  transition  input  output  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	56 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59:  members (6) 
      -- CP-element group 59: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_233_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_233_update_start_
      -- CP-element group 59: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_233_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_233_Sample/ra
      -- CP-element group 59: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_233_Update/$entry
      -- CP-element group 59: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_233_Update/cr
      -- 
    ra_728_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_233_inst_ack_0, ack => testConfigure_CP_0_elements(59)); -- 
    cr_732_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_732_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(59), ack => RPIPE_ConvTranspose_input_pipe_233_inst_req_1); -- 
    -- CP-element group 60:  fork  transition  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60: 	66 
    -- CP-element group 60:  members (9) 
      -- CP-element group 60: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_258_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_258_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_258_Sample/rr
      -- CP-element group 60: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_233_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_233_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_233_Update/ca
      -- CP-element group 60: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_237_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_237_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_237_Sample/rr
      -- 
    ca_733_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_233_inst_ack_1, ack => testConfigure_CP_0_elements(60)); -- 
    rr_741_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_741_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(60), ack => type_cast_237_inst_req_0); -- 
    rr_805_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_805_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(60), ack => RPIPE_ConvTranspose_input_pipe_258_inst_req_0); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_237_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_237_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_237_Sample/ra
      -- 
    ra_742_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_237_inst_ack_0, ack => testConfigure_CP_0_elements(61)); -- 
    -- CP-element group 62:  fork  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	56 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62: 	70 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_237_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_237_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_237_Update/ca
      -- 
    ca_747_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_237_inst_ack_1, ack => testConfigure_CP_0_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	56 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (9) 
      -- CP-element group 63: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_248_Sample/ptr_deref_248_Split/split_req
      -- CP-element group 63: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_248_Sample/ptr_deref_248_Split/split_ack
      -- CP-element group 63: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_248_Sample/word_access_start/$entry
      -- CP-element group 63: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_248_Sample/word_access_start/word_0/$entry
      -- CP-element group 63: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_248_Sample/word_access_start/word_0/rr
      -- CP-element group 63: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_248_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_248_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_248_Sample/ptr_deref_248_Split/$entry
      -- CP-element group 63: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_248_Sample/ptr_deref_248_Split/$exit
      -- 
    rr_785_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_785_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(63), ack => ptr_deref_248_store_0_req_0); -- 
    testConfigure_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(56) & testConfigure_CP_0_elements(62);
      gj_testConfigure_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	115 
    -- CP-element group 64:  members (5) 
      -- CP-element group 64: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_248_Sample/word_access_start/$exit
      -- CP-element group 64: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_248_Sample/word_access_start/word_0/$exit
      -- CP-element group 64: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_248_Sample/word_access_start/word_0/ra
      -- CP-element group 64: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_248_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_248_Sample/$exit
      -- 
    ra_786_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_248_store_0_ack_0, ack => testConfigure_CP_0_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	56 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	120 
    -- CP-element group 65:  members (5) 
      -- CP-element group 65: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_248_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_248_Update/word_access_complete/$exit
      -- CP-element group 65: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_248_Update/word_access_complete/word_0/$exit
      -- CP-element group 65: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_248_Update/word_access_complete/word_0/ca
      -- CP-element group 65: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_248_update_completed_
      -- 
    ca_797_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_248_store_0_ack_1, ack => testConfigure_CP_0_elements(65)); -- 
    -- CP-element group 66:  transition  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	60 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (6) 
      -- CP-element group 66: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_258_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_258_update_start_
      -- CP-element group 66: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_258_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_258_Sample/ra
      -- CP-element group 66: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_258_Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_258_Update/cr
      -- 
    ra_806_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_258_inst_ack_0, ack => testConfigure_CP_0_elements(66)); -- 
    cr_810_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_810_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(66), ack => RPIPE_ConvTranspose_input_pipe_258_inst_req_1); -- 
    -- CP-element group 67:  fork  transition  input  output  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67: 	73 
    -- CP-element group 67:  members (9) 
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_258_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_258_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_258_Update/ca
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_262_sample_start_
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_262_Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_262_Sample/rr
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_282_sample_start_
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_282_Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_282_Sample/rr
      -- 
    ca_811_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_258_inst_ack_1, ack => testConfigure_CP_0_elements(67)); -- 
    rr_819_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_819_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(67), ack => type_cast_262_inst_req_0); -- 
    rr_883_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_883_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(67), ack => RPIPE_ConvTranspose_input_pipe_282_inst_req_0); -- 
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_262_sample_completed_
      -- CP-element group 68: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_262_Sample/$exit
      -- CP-element group 68: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_262_Sample/ra
      -- 
    ra_820_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_262_inst_ack_0, ack => testConfigure_CP_0_elements(68)); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	56 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_262_update_completed_
      -- CP-element group 69: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_262_Update/$exit
      -- CP-element group 69: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_262_Update/ca
      -- 
    ca_825_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_262_inst_ack_1, ack => testConfigure_CP_0_elements(69)); -- 
    -- CP-element group 70:  join  transition  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	56 
    -- CP-element group 70: 	62 
    -- CP-element group 70: 	69 
    -- CP-element group 70: 	115 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70:  members (9) 
      -- CP-element group 70: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_278_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_278_Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_278_Sample/ptr_deref_278_Split/$entry
      -- CP-element group 70: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_278_Sample/ptr_deref_278_Split/$exit
      -- CP-element group 70: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_278_Sample/ptr_deref_278_Split/split_req
      -- CP-element group 70: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_278_Sample/ptr_deref_278_Split/split_ack
      -- CP-element group 70: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_278_Sample/word_access_start/$entry
      -- CP-element group 70: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_278_Sample/word_access_start/word_0/$entry
      -- CP-element group 70: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_278_Sample/word_access_start/word_0/rr
      -- 
    rr_863_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_863_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(70), ack => ptr_deref_278_store_0_req_0); -- 
    testConfigure_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(56) & testConfigure_CP_0_elements(62) & testConfigure_CP_0_elements(69) & testConfigure_CP_0_elements(115);
      gj_testConfigure_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	116 
    -- CP-element group 71:  members (5) 
      -- CP-element group 71: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_278_sample_completed_
      -- CP-element group 71: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_278_Sample/$exit
      -- CP-element group 71: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_278_Sample/word_access_start/$exit
      -- CP-element group 71: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_278_Sample/word_access_start/word_0/$exit
      -- CP-element group 71: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_278_Sample/word_access_start/word_0/ra
      -- 
    ra_864_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_278_store_0_ack_0, ack => testConfigure_CP_0_elements(71)); -- 
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	56 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	120 
    -- CP-element group 72:  members (5) 
      -- CP-element group 72: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_278_update_completed_
      -- CP-element group 72: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_278_Update/$exit
      -- CP-element group 72: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_278_Update/word_access_complete/$exit
      -- CP-element group 72: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_278_Update/word_access_complete/word_0/$exit
      -- CP-element group 72: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_278_Update/word_access_complete/word_0/ca
      -- 
    ca_875_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_278_store_0_ack_1, ack => testConfigure_CP_0_elements(72)); -- 
    -- CP-element group 73:  transition  input  output  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	67 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (6) 
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_282_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_282_update_start_
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_282_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_282_Sample/ra
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_282_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_282_Update/cr
      -- 
    ra_884_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_282_inst_ack_0, ack => testConfigure_CP_0_elements(73)); -- 
    cr_888_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_888_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => RPIPE_ConvTranspose_input_pipe_282_inst_req_1); -- 
    -- CP-element group 74:  fork  transition  input  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74: 	80 
    -- CP-element group 74:  members (9) 
      -- CP-element group 74: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_282_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_282_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_282_Update/ca
      -- CP-element group 74: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_286_sample_start_
      -- CP-element group 74: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_286_Sample/$entry
      -- CP-element group 74: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_286_Sample/rr
      -- CP-element group 74: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_307_sample_start_
      -- CP-element group 74: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_307_Sample/$entry
      -- CP-element group 74: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_307_Sample/rr
      -- 
    ca_889_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_282_inst_ack_1, ack => testConfigure_CP_0_elements(74)); -- 
    rr_897_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_897_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(74), ack => type_cast_286_inst_req_0); -- 
    rr_961_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_961_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(74), ack => RPIPE_ConvTranspose_input_pipe_307_inst_req_0); -- 
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_286_sample_completed_
      -- CP-element group 75: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_286_Sample/$exit
      -- CP-element group 75: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_286_Sample/ra
      -- 
    ra_898_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_286_inst_ack_0, ack => testConfigure_CP_0_elements(75)); -- 
    -- CP-element group 76:  fork  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	56 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76: 	84 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_286_update_completed_
      -- CP-element group 76: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_286_Update/$exit
      -- CP-element group 76: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_286_Update/ca
      -- 
    ca_903_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_286_inst_ack_1, ack => testConfigure_CP_0_elements(76)); -- 
    -- CP-element group 77:  join  transition  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	56 
    -- CP-element group 77: 	76 
    -- CP-element group 77: 	116 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (9) 
      -- CP-element group 77: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_297_sample_start_
      -- CP-element group 77: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_297_Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_297_Sample/ptr_deref_297_Split/$entry
      -- CP-element group 77: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_297_Sample/ptr_deref_297_Split/$exit
      -- CP-element group 77: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_297_Sample/ptr_deref_297_Split/split_req
      -- CP-element group 77: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_297_Sample/ptr_deref_297_Split/split_ack
      -- CP-element group 77: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_297_Sample/word_access_start/$entry
      -- CP-element group 77: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_297_Sample/word_access_start/word_0/$entry
      -- CP-element group 77: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_297_Sample/word_access_start/word_0/rr
      -- 
    rr_941_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_941_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => ptr_deref_297_store_0_req_0); -- 
    testConfigure_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(56) & testConfigure_CP_0_elements(76) & testConfigure_CP_0_elements(116);
      gj_testConfigure_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	117 
    -- CP-element group 78:  members (5) 
      -- CP-element group 78: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_297_sample_completed_
      -- CP-element group 78: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_297_Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_297_Sample/word_access_start/$exit
      -- CP-element group 78: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_297_Sample/word_access_start/word_0/$exit
      -- CP-element group 78: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_297_Sample/word_access_start/word_0/ra
      -- 
    ra_942_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_297_store_0_ack_0, ack => testConfigure_CP_0_elements(78)); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	56 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	120 
    -- CP-element group 79:  members (5) 
      -- CP-element group 79: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_297_update_completed_
      -- CP-element group 79: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_297_Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_297_Update/word_access_complete/$exit
      -- CP-element group 79: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_297_Update/word_access_complete/word_0/$exit
      -- CP-element group 79: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_297_Update/word_access_complete/word_0/ca
      -- 
    ca_953_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_297_store_0_ack_1, ack => testConfigure_CP_0_elements(79)); -- 
    -- CP-element group 80:  transition  input  output  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	74 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (6) 
      -- CP-element group 80: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_307_sample_completed_
      -- CP-element group 80: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_307_update_start_
      -- CP-element group 80: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_307_Sample/$exit
      -- CP-element group 80: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_307_Sample/ra
      -- CP-element group 80: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_307_Update/$entry
      -- CP-element group 80: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_307_Update/cr
      -- 
    ra_962_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_307_inst_ack_0, ack => testConfigure_CP_0_elements(80)); -- 
    cr_966_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_966_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(80), ack => RPIPE_ConvTranspose_input_pipe_307_inst_req_1); -- 
    -- CP-element group 81:  fork  transition  input  output  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	82 
    -- CP-element group 81: 	87 
    -- CP-element group 81:  members (9) 
      -- CP-element group 81: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_307_update_completed_
      -- CP-element group 81: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_307_Update/$exit
      -- CP-element group 81: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_307_Update/ca
      -- CP-element group 81: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_311_sample_start_
      -- CP-element group 81: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_311_Sample/$entry
      -- CP-element group 81: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_311_Sample/rr
      -- CP-element group 81: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_331_sample_start_
      -- CP-element group 81: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_331_Sample/$entry
      -- CP-element group 81: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_331_Sample/rr
      -- 
    ca_967_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_307_inst_ack_1, ack => testConfigure_CP_0_elements(81)); -- 
    rr_975_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_975_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(81), ack => type_cast_311_inst_req_0); -- 
    rr_1039_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1039_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(81), ack => RPIPE_ConvTranspose_input_pipe_331_inst_req_0); -- 
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	81 
    -- CP-element group 82: successors 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_311_sample_completed_
      -- CP-element group 82: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_311_Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_311_Sample/ra
      -- 
    ra_976_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_311_inst_ack_0, ack => testConfigure_CP_0_elements(82)); -- 
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	56 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_311_update_completed_
      -- CP-element group 83: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_311_Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_311_Update/ca
      -- 
    ca_981_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_311_inst_ack_1, ack => testConfigure_CP_0_elements(83)); -- 
    -- CP-element group 84:  join  transition  output  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	56 
    -- CP-element group 84: 	76 
    -- CP-element group 84: 	83 
    -- CP-element group 84: 	117 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84:  members (9) 
      -- CP-element group 84: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_327_sample_start_
      -- CP-element group 84: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_327_Sample/$entry
      -- CP-element group 84: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_327_Sample/ptr_deref_327_Split/$entry
      -- CP-element group 84: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_327_Sample/ptr_deref_327_Split/$exit
      -- CP-element group 84: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_327_Sample/ptr_deref_327_Split/split_req
      -- CP-element group 84: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_327_Sample/ptr_deref_327_Split/split_ack
      -- CP-element group 84: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_327_Sample/word_access_start/$entry
      -- CP-element group 84: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_327_Sample/word_access_start/word_0/$entry
      -- CP-element group 84: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_327_Sample/word_access_start/word_0/rr
      -- 
    rr_1019_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1019_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(84), ack => ptr_deref_327_store_0_req_0); -- 
    testConfigure_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(56) & testConfigure_CP_0_elements(76) & testConfigure_CP_0_elements(83) & testConfigure_CP_0_elements(117);
      gj_testConfigure_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	118 
    -- CP-element group 85:  members (5) 
      -- CP-element group 85: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_327_sample_completed_
      -- CP-element group 85: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_327_Sample/$exit
      -- CP-element group 85: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_327_Sample/word_access_start/$exit
      -- CP-element group 85: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_327_Sample/word_access_start/word_0/$exit
      -- CP-element group 85: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_327_Sample/word_access_start/word_0/ra
      -- 
    ra_1020_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_327_store_0_ack_0, ack => testConfigure_CP_0_elements(85)); -- 
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	56 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	120 
    -- CP-element group 86:  members (5) 
      -- CP-element group 86: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_327_update_completed_
      -- CP-element group 86: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_327_Update/$exit
      -- CP-element group 86: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_327_Update/word_access_complete/$exit
      -- CP-element group 86: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_327_Update/word_access_complete/word_0/$exit
      -- CP-element group 86: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_327_Update/word_access_complete/word_0/ca
      -- 
    ca_1031_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_327_store_0_ack_1, ack => testConfigure_CP_0_elements(86)); -- 
    -- CP-element group 87:  transition  input  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	81 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (6) 
      -- CP-element group 87: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_331_sample_completed_
      -- CP-element group 87: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_331_update_start_
      -- CP-element group 87: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_331_Sample/$exit
      -- CP-element group 87: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_331_Sample/ra
      -- CP-element group 87: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_331_Update/$entry
      -- CP-element group 87: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_331_Update/cr
      -- 
    ra_1040_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_331_inst_ack_0, ack => testConfigure_CP_0_elements(87)); -- 
    cr_1044_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1044_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(87), ack => RPIPE_ConvTranspose_input_pipe_331_inst_req_1); -- 
    -- CP-element group 88:  fork  transition  input  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	89 
    -- CP-element group 88: 	94 
    -- CP-element group 88:  members (9) 
      -- CP-element group 88: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_356_Sample/rr
      -- CP-element group 88: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_356_Sample/$entry
      -- CP-element group 88: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_356_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_331_update_completed_
      -- CP-element group 88: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_331_Update/$exit
      -- CP-element group 88: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_331_Update/ca
      -- CP-element group 88: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_335_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_335_Sample/$entry
      -- CP-element group 88: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_335_Sample/rr
      -- 
    ca_1045_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_331_inst_ack_1, ack => testConfigure_CP_0_elements(88)); -- 
    rr_1053_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1053_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(88), ack => type_cast_335_inst_req_0); -- 
    rr_1117_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1117_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(88), ack => RPIPE_ConvTranspose_input_pipe_356_inst_req_0); -- 
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	88 
    -- CP-element group 89: successors 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_335_sample_completed_
      -- CP-element group 89: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_335_Sample/$exit
      -- CP-element group 89: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_335_Sample/ra
      -- 
    ra_1054_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_335_inst_ack_0, ack => testConfigure_CP_0_elements(89)); -- 
    -- CP-element group 90:  fork  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	56 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90: 	98 
    -- CP-element group 90:  members (3) 
      -- CP-element group 90: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_335_update_completed_
      -- CP-element group 90: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_335_Update/$exit
      -- CP-element group 90: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_335_Update/ca
      -- 
    ca_1059_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_335_inst_ack_1, ack => testConfigure_CP_0_elements(90)); -- 
    -- CP-element group 91:  join  transition  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	56 
    -- CP-element group 91: 	90 
    -- CP-element group 91: 	118 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (9) 
      -- CP-element group 91: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_346_Sample/ptr_deref_346_Split/split_req
      -- CP-element group 91: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_346_Sample/ptr_deref_346_Split/$exit
      -- CP-element group 91: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_346_Sample/ptr_deref_346_Split/$entry
      -- CP-element group 91: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_346_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_346_Sample/word_access_start/word_0/rr
      -- CP-element group 91: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_346_Sample/word_access_start/word_0/$entry
      -- CP-element group 91: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_346_Sample/word_access_start/$entry
      -- CP-element group 91: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_346_Sample/ptr_deref_346_Split/split_ack
      -- CP-element group 91: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_346_sample_start_
      -- 
    rr_1097_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1097_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(91), ack => ptr_deref_346_store_0_req_0); -- 
    testConfigure_cp_element_group_91: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_91"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(56) & testConfigure_CP_0_elements(90) & testConfigure_CP_0_elements(118);
      gj_testConfigure_cp_element_group_91 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(91), clk => clk, reset => reset); --
    end block;
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	119 
    -- CP-element group 92:  members (5) 
      -- CP-element group 92: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_346_Sample/$exit
      -- CP-element group 92: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_346_Sample/word_access_start/word_0/ra
      -- CP-element group 92: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_346_Sample/word_access_start/word_0/$exit
      -- CP-element group 92: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_346_Sample/word_access_start/$exit
      -- CP-element group 92: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_346_sample_completed_
      -- 
    ra_1098_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_346_store_0_ack_0, ack => testConfigure_CP_0_elements(92)); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	56 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	120 
    -- CP-element group 93:  members (5) 
      -- CP-element group 93: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_346_Update/word_access_complete/word_0/ca
      -- CP-element group 93: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_346_Update/word_access_complete/word_0/$exit
      -- CP-element group 93: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_346_Update/word_access_complete/$exit
      -- CP-element group 93: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_346_Update/$exit
      -- CP-element group 93: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_346_update_completed_
      -- 
    ca_1109_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_346_store_0_ack_1, ack => testConfigure_CP_0_elements(93)); -- 
    -- CP-element group 94:  transition  input  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	88 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94:  members (6) 
      -- CP-element group 94: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_356_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_356_Update/cr
      -- CP-element group 94: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_356_Sample/ra
      -- CP-element group 94: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_356_Sample/$exit
      -- CP-element group 94: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_356_update_start_
      -- CP-element group 94: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_356_sample_completed_
      -- 
    ra_1118_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_356_inst_ack_0, ack => testConfigure_CP_0_elements(94)); -- 
    cr_1122_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1122_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(94), ack => RPIPE_ConvTranspose_input_pipe_356_inst_req_1); -- 
    -- CP-element group 95:  transition  input  output  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95:  members (6) 
      -- CP-element group 95: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_360_Sample/$entry
      -- CP-element group 95: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_360_sample_start_
      -- CP-element group 95: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_356_Update/ca
      -- CP-element group 95: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_356_Update/$exit
      -- CP-element group 95: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/RPIPE_ConvTranspose_input_pipe_356_update_completed_
      -- CP-element group 95: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_360_Sample/rr
      -- 
    ca_1123_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_356_inst_ack_1, ack => testConfigure_CP_0_elements(95)); -- 
    rr_1131_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1131_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(95), ack => type_cast_360_inst_req_0); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_360_Sample/$exit
      -- CP-element group 96: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_360_sample_completed_
      -- CP-element group 96: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_360_Sample/ra
      -- 
    ra_1132_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_360_inst_ack_0, ack => testConfigure_CP_0_elements(96)); -- 
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	56 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_360_update_completed_
      -- CP-element group 97: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_360_Update/ca
      -- CP-element group 97: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/type_cast_360_Update/$exit
      -- 
    ca_1137_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_360_inst_ack_1, ack => testConfigure_CP_0_elements(97)); -- 
    -- CP-element group 98:  join  transition  output  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	56 
    -- CP-element group 98: 	90 
    -- CP-element group 98: 	97 
    -- CP-element group 98: 	119 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (9) 
      -- CP-element group 98: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_376_Sample/ptr_deref_376_Split/$exit
      -- CP-element group 98: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_376_Sample/ptr_deref_376_Split/$entry
      -- CP-element group 98: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_376_Sample/$entry
      -- CP-element group 98: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_376_Sample/word_access_start/$entry
      -- CP-element group 98: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_376_Sample/ptr_deref_376_Split/split_ack
      -- CP-element group 98: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_376_sample_start_
      -- CP-element group 98: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_376_Sample/word_access_start/word_0/rr
      -- CP-element group 98: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_376_Sample/word_access_start/word_0/$entry
      -- CP-element group 98: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_376_Sample/ptr_deref_376_Split/split_req
      -- 
    rr_1175_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1175_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(98), ack => ptr_deref_376_store_0_req_0); -- 
    testConfigure_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(56) & testConfigure_CP_0_elements(90) & testConfigure_CP_0_elements(97) & testConfigure_CP_0_elements(119);
      gj_testConfigure_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99:  members (5) 
      -- CP-element group 99: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_376_Sample/$exit
      -- CP-element group 99: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_376_sample_completed_
      -- CP-element group 99: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_376_Sample/word_access_start/word_0/ra
      -- CP-element group 99: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_376_Sample/word_access_start/word_0/$exit
      -- CP-element group 99: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_376_Sample/word_access_start/$exit
      -- 
    ra_1176_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_376_store_0_ack_0, ack => testConfigure_CP_0_elements(99)); -- 
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	56 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	120 
    -- CP-element group 100:  members (5) 
      -- CP-element group 100: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_376_Update/word_access_complete/word_0/ca
      -- CP-element group 100: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_376_Update/word_access_complete/word_0/$exit
      -- CP-element group 100: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_376_Update/word_access_complete/$exit
      -- CP-element group 100: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_376_Update/$exit
      -- CP-element group 100: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_376_update_completed_
      -- 
    ca_1187_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_376_store_0_ack_1, ack => testConfigure_CP_0_elements(100)); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	56 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (5) 
      -- CP-element group 101: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_389_sample_completed_
      -- CP-element group 101: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_389_Sample/word_access_start/word_0/ra
      -- CP-element group 101: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_389_Sample/word_access_start/word_0/$exit
      -- CP-element group 101: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_389_Sample/word_access_start/$exit
      -- CP-element group 101: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_389_Sample/$exit
      -- 
    ra_1221_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_389_load_0_ack_0, ack => testConfigure_CP_0_elements(101)); -- 
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	56 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	120 
    -- CP-element group 102:  members (9) 
      -- CP-element group 102: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_389_update_completed_
      -- CP-element group 102: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_389_Update/ptr_deref_389_Merge/merge_ack
      -- CP-element group 102: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_389_Update/ptr_deref_389_Merge/merge_req
      -- CP-element group 102: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_389_Update/ptr_deref_389_Merge/$exit
      -- CP-element group 102: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_389_Update/ptr_deref_389_Merge/$entry
      -- CP-element group 102: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_389_Update/word_access_complete/word_0/ca
      -- CP-element group 102: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_389_Update/word_access_complete/word_0/$exit
      -- CP-element group 102: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_389_Update/word_access_complete/$exit
      -- CP-element group 102: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_389_Update/$exit
      -- 
    ca_1232_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_389_load_0_ack_1, ack => testConfigure_CP_0_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	56 
    -- CP-element group 103: successors 
    -- CP-element group 103:  members (5) 
      -- CP-element group 103: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_401_sample_completed_
      -- CP-element group 103: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_401_Sample/word_access_start/word_0/$exit
      -- CP-element group 103: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_401_Sample/word_access_start/word_0/ra
      -- CP-element group 103: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_401_Sample/word_access_start/$exit
      -- CP-element group 103: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_401_Sample/$exit
      -- 
    ra_1271_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_401_load_0_ack_0, ack => testConfigure_CP_0_elements(103)); -- 
    -- CP-element group 104:  transition  input  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	56 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	120 
    -- CP-element group 104:  members (9) 
      -- CP-element group 104: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_401_update_completed_
      -- CP-element group 104: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_401_Update/ptr_deref_401_Merge/merge_ack
      -- CP-element group 104: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_401_Update/ptr_deref_401_Merge/merge_req
      -- CP-element group 104: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_401_Update/ptr_deref_401_Merge/$exit
      -- CP-element group 104: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_401_Update/ptr_deref_401_Merge/$entry
      -- CP-element group 104: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_401_Update/word_access_complete/word_0/ca
      -- CP-element group 104: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_401_Update/word_access_complete/word_0/$exit
      -- CP-element group 104: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_401_Update/word_access_complete/$exit
      -- CP-element group 104: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_401_Update/$exit
      -- 
    ca_1282_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_401_load_0_ack_1, ack => testConfigure_CP_0_elements(104)); -- 
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	56 
    -- CP-element group 105: successors 
    -- CP-element group 105:  members (5) 
      -- CP-element group 105: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_413_sample_completed_
      -- CP-element group 105: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_413_Sample/word_access_start/word_0/ra
      -- CP-element group 105: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_413_Sample/word_access_start/word_0/$exit
      -- CP-element group 105: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_413_Sample/word_access_start/$exit
      -- CP-element group 105: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_413_Sample/$exit
      -- 
    ra_1321_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_413_load_0_ack_0, ack => testConfigure_CP_0_elements(105)); -- 
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	56 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	120 
    -- CP-element group 106:  members (9) 
      -- CP-element group 106: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_413_Update/ptr_deref_413_Merge/merge_ack
      -- CP-element group 106: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_413_Update/ptr_deref_413_Merge/merge_req
      -- CP-element group 106: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_413_Update/ptr_deref_413_Merge/$exit
      -- CP-element group 106: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_413_Update/ptr_deref_413_Merge/$entry
      -- CP-element group 106: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_413_update_completed_
      -- CP-element group 106: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_413_Update/word_access_complete/word_0/ca
      -- CP-element group 106: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_413_Update/word_access_complete/word_0/$exit
      -- CP-element group 106: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_413_Update/word_access_complete/$exit
      -- CP-element group 106: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_413_Update/$exit
      -- 
    ca_1332_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_413_load_0_ack_1, ack => testConfigure_CP_0_elements(106)); -- 
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	56 
    -- CP-element group 107: successors 
    -- CP-element group 107:  members (5) 
      -- CP-element group 107: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_435_Sample/$exit
      -- CP-element group 107: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_435_Sample/word_access_start/$exit
      -- CP-element group 107: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_435_sample_completed_
      -- CP-element group 107: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_435_Sample/word_access_start/word_0/ra
      -- CP-element group 107: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_435_Sample/word_access_start/word_0/$exit
      -- 
    ra_1371_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_435_load_0_ack_0, ack => testConfigure_CP_0_elements(107)); -- 
    -- CP-element group 108:  transition  input  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	56 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	120 
    -- CP-element group 108:  members (9) 
      -- CP-element group 108: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_435_Update/ptr_deref_435_Merge/merge_ack
      -- CP-element group 108: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_435_update_completed_
      -- CP-element group 108: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_435_Update/ptr_deref_435_Merge/merge_req
      -- CP-element group 108: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_435_Update/ptr_deref_435_Merge/$exit
      -- CP-element group 108: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_435_Update/ptr_deref_435_Merge/$entry
      -- CP-element group 108: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_435_Update/word_access_complete/word_0/ca
      -- CP-element group 108: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_435_Update/word_access_complete/word_0/$exit
      -- CP-element group 108: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_435_Update/word_access_complete/$exit
      -- CP-element group 108: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_435_Update/$exit
      -- 
    ca_1382_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_435_load_0_ack_1, ack => testConfigure_CP_0_elements(108)); -- 
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	56 
    -- CP-element group 109: successors 
    -- CP-element group 109:  members (5) 
      -- CP-element group 109: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_447_Sample/word_access_start/$exit
      -- CP-element group 109: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_447_Sample/$exit
      -- CP-element group 109: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_447_sample_completed_
      -- CP-element group 109: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_447_Sample/word_access_start/word_0/ra
      -- CP-element group 109: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_447_Sample/word_access_start/word_0/$exit
      -- 
    ra_1421_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_447_load_0_ack_0, ack => testConfigure_CP_0_elements(109)); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	56 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	120 
    -- CP-element group 110:  members (9) 
      -- CP-element group 110: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_447_Update/ptr_deref_447_Merge/merge_ack
      -- CP-element group 110: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_447_Update/ptr_deref_447_Merge/merge_req
      -- CP-element group 110: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_447_Update/ptr_deref_447_Merge/$exit
      -- CP-element group 110: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_447_Update/ptr_deref_447_Merge/$entry
      -- CP-element group 110: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_447_Update/word_access_complete/word_0/ca
      -- CP-element group 110: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_447_update_completed_
      -- CP-element group 110: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_447_Update/word_access_complete/word_0/$exit
      -- CP-element group 110: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_447_Update/word_access_complete/$exit
      -- CP-element group 110: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_447_Update/$exit
      -- 
    ca_1432_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_447_load_0_ack_1, ack => testConfigure_CP_0_elements(110)); -- 
    -- CP-element group 111:  transition  input  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	56 
    -- CP-element group 111: successors 
    -- CP-element group 111:  members (5) 
      -- CP-element group 111: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_459_Sample/word_access_start/word_0/$exit
      -- CP-element group 111: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_459_Sample/word_access_start/$exit
      -- CP-element group 111: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_459_Sample/$exit
      -- CP-element group 111: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_459_sample_completed_
      -- CP-element group 111: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_459_Sample/word_access_start/word_0/ra
      -- 
    ra_1471_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_459_load_0_ack_0, ack => testConfigure_CP_0_elements(111)); -- 
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	56 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	120 
    -- CP-element group 112:  members (9) 
      -- CP-element group 112: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_459_Update/word_access_complete/word_0/ca
      -- CP-element group 112: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_459_Update/ptr_deref_459_Merge/merge_ack
      -- CP-element group 112: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_459_Update/word_access_complete/word_0/$exit
      -- CP-element group 112: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_459_update_completed_
      -- CP-element group 112: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_459_Update/ptr_deref_459_Merge/merge_req
      -- CP-element group 112: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_459_Update/word_access_complete/$exit
      -- CP-element group 112: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_459_Update/ptr_deref_459_Merge/$exit
      -- CP-element group 112: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_459_Update/$exit
      -- CP-element group 112: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_459_Update/ptr_deref_459_Merge/$entry
      -- 
    ca_1482_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_459_load_0_ack_1, ack => testConfigure_CP_0_elements(112)); -- 
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	56 
    -- CP-element group 113: successors 
    -- CP-element group 113:  members (5) 
      -- CP-element group 113: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_471_sample_completed_
      -- CP-element group 113: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_471_Sample/word_access_start/word_0/ra
      -- CP-element group 113: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_471_Sample/word_access_start/word_0/$exit
      -- CP-element group 113: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_471_Sample/word_access_start/$exit
      -- CP-element group 113: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_471_Sample/$exit
      -- 
    ra_1521_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_471_load_0_ack_0, ack => testConfigure_CP_0_elements(113)); -- 
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	56 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	120 
    -- CP-element group 114:  members (9) 
      -- CP-element group 114: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_471_Update/word_access_complete/word_0/$exit
      -- CP-element group 114: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_471_Update/ptr_deref_471_Merge/$entry
      -- CP-element group 114: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_471_Update/ptr_deref_471_Merge/$exit
      -- CP-element group 114: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_471_Update/ptr_deref_471_Merge/merge_req
      -- CP-element group 114: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_471_Update/ptr_deref_471_Merge/merge_ack
      -- CP-element group 114: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_471_Update/word_access_complete/word_0/ca
      -- CP-element group 114: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_471_Update/word_access_complete/$exit
      -- CP-element group 114: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_471_Update/$exit
      -- CP-element group 114: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_471_update_completed_
      -- 
    ca_1532_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_471_load_0_ack_1, ack => testConfigure_CP_0_elements(114)); -- 
    -- CP-element group 115:  transition  delay-element  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	64 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	70 
    -- CP-element group 115:  members (1) 
      -- CP-element group 115: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_248_ptr_deref_278_delay
      -- 
    -- Element group testConfigure_CP_0_elements(115) is a control-delay.
    cp_element_115_delay: control_delay_element  generic map(name => " 115_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(64), ack => testConfigure_CP_0_elements(115), clk => clk, reset =>reset);
    -- CP-element group 116:  transition  delay-element  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	71 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	77 
    -- CP-element group 116:  members (1) 
      -- CP-element group 116: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_278_ptr_deref_297_delay
      -- 
    -- Element group testConfigure_CP_0_elements(116) is a control-delay.
    cp_element_116_delay: control_delay_element  generic map(name => " 116_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(71), ack => testConfigure_CP_0_elements(116), clk => clk, reset =>reset);
    -- CP-element group 117:  transition  delay-element  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	78 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	84 
    -- CP-element group 117:  members (1) 
      -- CP-element group 117: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_297_ptr_deref_327_delay
      -- 
    -- Element group testConfigure_CP_0_elements(117) is a control-delay.
    cp_element_117_delay: control_delay_element  generic map(name => " 117_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(78), ack => testConfigure_CP_0_elements(117), clk => clk, reset =>reset);
    -- CP-element group 118:  transition  delay-element  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	85 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	91 
    -- CP-element group 118:  members (1) 
      -- CP-element group 118: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_327_ptr_deref_346_delay
      -- 
    -- Element group testConfigure_CP_0_elements(118) is a control-delay.
    cp_element_118_delay: control_delay_element  generic map(name => " 118_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(85), ack => testConfigure_CP_0_elements(118), clk => clk, reset =>reset);
    -- CP-element group 119:  transition  delay-element  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	92 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	98 
    -- CP-element group 119:  members (1) 
      -- CP-element group 119: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/ptr_deref_346_ptr_deref_376_delay
      -- 
    -- Element group testConfigure_CP_0_elements(119) is a control-delay.
    cp_element_119_delay: control_delay_element  generic map(name => " 119_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(92), ack => testConfigure_CP_0_elements(119), clk => clk, reset =>reset);
    -- CP-element group 120:  branch  join  transition  place  output  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	58 
    -- CP-element group 120: 	65 
    -- CP-element group 120: 	72 
    -- CP-element group 120: 	79 
    -- CP-element group 120: 	86 
    -- CP-element group 120: 	93 
    -- CP-element group 120: 	100 
    -- CP-element group 120: 	102 
    -- CP-element group 120: 	104 
    -- CP-element group 120: 	106 
    -- CP-element group 120: 	108 
    -- CP-element group 120: 	110 
    -- CP-element group 120: 	112 
    -- CP-element group 120: 	114 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120: 	122 
    -- CP-element group 120:  members (10) 
      -- CP-element group 120: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493__exit__
      -- CP-element group 120: 	 branch_block_stmt_34/if_stmt_494__entry__
      -- CP-element group 120: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493/$exit
      -- CP-element group 120: 	 branch_block_stmt_34/if_stmt_494_dead_link/$entry
      -- CP-element group 120: 	 branch_block_stmt_34/if_stmt_494_eval_test/$entry
      -- CP-element group 120: 	 branch_block_stmt_34/if_stmt_494_eval_test/$exit
      -- CP-element group 120: 	 branch_block_stmt_34/if_stmt_494_eval_test/branch_req
      -- CP-element group 120: 	 branch_block_stmt_34/R_cmp88233_495_place
      -- CP-element group 120: 	 branch_block_stmt_34/if_stmt_494_if_link/$entry
      -- CP-element group 120: 	 branch_block_stmt_34/if_stmt_494_else_link/$entry
      -- 
    branch_req_1550_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1550_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(120), ack => if_stmt_494_branch_req_0); -- 
    testConfigure_cp_element_group_120: block -- 
      constant place_capacities: IntegerArray(0 to 13) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1);
      constant place_markings: IntegerArray(0 to 13)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0);
      constant place_delays: IntegerArray(0 to 13) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_120"; 
      signal preds: BooleanArray(1 to 14); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(58) & testConfigure_CP_0_elements(65) & testConfigure_CP_0_elements(72) & testConfigure_CP_0_elements(79) & testConfigure_CP_0_elements(86) & testConfigure_CP_0_elements(93) & testConfigure_CP_0_elements(100) & testConfigure_CP_0_elements(102) & testConfigure_CP_0_elements(104) & testConfigure_CP_0_elements(106) & testConfigure_CP_0_elements(108) & testConfigure_CP_0_elements(110) & testConfigure_CP_0_elements(112) & testConfigure_CP_0_elements(114);
      gj_testConfigure_cp_element_group_120 : generic_join generic map(name => joinName, number_of_predecessors => 14, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(120), clk => clk, reset => reset); --
    end block;
    -- CP-element group 121:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	125 
    -- CP-element group 121: 	126 
    -- CP-element group 121:  members (18) 
      -- CP-element group 121: 	 branch_block_stmt_34/merge_stmt_515__exit__
      -- CP-element group 121: 	 branch_block_stmt_34/assign_stmt_521_to_assign_stmt_550__entry__
      -- CP-element group 121: 	 branch_block_stmt_34/if_stmt_494_if_link/$exit
      -- CP-element group 121: 	 branch_block_stmt_34/if_stmt_494_if_link/if_choice_transition
      -- CP-element group 121: 	 branch_block_stmt_34/forx_xend49_bbx_xnph235
      -- CP-element group 121: 	 branch_block_stmt_34/assign_stmt_521_to_assign_stmt_550/$entry
      -- CP-element group 121: 	 branch_block_stmt_34/assign_stmt_521_to_assign_stmt_550/type_cast_536_sample_start_
      -- CP-element group 121: 	 branch_block_stmt_34/assign_stmt_521_to_assign_stmt_550/type_cast_536_update_start_
      -- CP-element group 121: 	 branch_block_stmt_34/assign_stmt_521_to_assign_stmt_550/type_cast_536_Sample/$entry
      -- CP-element group 121: 	 branch_block_stmt_34/assign_stmt_521_to_assign_stmt_550/type_cast_536_Sample/rr
      -- CP-element group 121: 	 branch_block_stmt_34/assign_stmt_521_to_assign_stmt_550/type_cast_536_Update/$entry
      -- CP-element group 121: 	 branch_block_stmt_34/assign_stmt_521_to_assign_stmt_550/type_cast_536_Update/cr
      -- CP-element group 121: 	 branch_block_stmt_34/forx_xend49_bbx_xnph235_PhiReq/$entry
      -- CP-element group 121: 	 branch_block_stmt_34/forx_xend49_bbx_xnph235_PhiReq/$exit
      -- CP-element group 121: 	 branch_block_stmt_34/merge_stmt_515_PhiReqMerge
      -- CP-element group 121: 	 branch_block_stmt_34/merge_stmt_515_PhiAck/$entry
      -- CP-element group 121: 	 branch_block_stmt_34/merge_stmt_515_PhiAck/$exit
      -- CP-element group 121: 	 branch_block_stmt_34/merge_stmt_515_PhiAck/dummy
      -- 
    if_choice_transition_1555_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_494_branch_ack_1, ack => testConfigure_CP_0_elements(121)); -- 
    rr_1594_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1594_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(121), ack => type_cast_536_inst_req_0); -- 
    cr_1599_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1599_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(121), ack => type_cast_536_inst_req_1); -- 
    -- CP-element group 122:  transition  place  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	120 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	265 
    -- CP-element group 122:  members (5) 
      -- CP-element group 122: 	 branch_block_stmt_34/if_stmt_494_else_link/$exit
      -- CP-element group 122: 	 branch_block_stmt_34/if_stmt_494_else_link/else_choice_transition
      -- CP-element group 122: 	 branch_block_stmt_34/forx_xend49_forx_xcond144x_xpreheader
      -- CP-element group 122: 	 branch_block_stmt_34/forx_xend49_forx_xcond144x_xpreheader_PhiReq/$entry
      -- CP-element group 122: 	 branch_block_stmt_34/forx_xend49_forx_xcond144x_xpreheader_PhiReq/$exit
      -- 
    else_choice_transition_1559_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_494_branch_ack_0, ack => testConfigure_CP_0_elements(122)); -- 
    -- CP-element group 123:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	265 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	169 
    -- CP-element group 123: 	170 
    -- CP-element group 123:  members (18) 
      -- CP-element group 123: 	 branch_block_stmt_34/merge_stmt_722__exit__
      -- CP-element group 123: 	 branch_block_stmt_34/assign_stmt_728_to_assign_stmt_757__entry__
      -- CP-element group 123: 	 branch_block_stmt_34/if_stmt_509_if_link/$exit
      -- CP-element group 123: 	 branch_block_stmt_34/if_stmt_509_if_link/if_choice_transition
      -- CP-element group 123: 	 branch_block_stmt_34/forx_xcond144x_xpreheader_bbx_xnph231
      -- CP-element group 123: 	 branch_block_stmt_34/assign_stmt_728_to_assign_stmt_757/$entry
      -- CP-element group 123: 	 branch_block_stmt_34/assign_stmt_728_to_assign_stmt_757/type_cast_743_sample_start_
      -- CP-element group 123: 	 branch_block_stmt_34/assign_stmt_728_to_assign_stmt_757/type_cast_743_update_start_
      -- CP-element group 123: 	 branch_block_stmt_34/assign_stmt_728_to_assign_stmt_757/type_cast_743_Sample/$entry
      -- CP-element group 123: 	 branch_block_stmt_34/assign_stmt_728_to_assign_stmt_757/type_cast_743_Sample/rr
      -- CP-element group 123: 	 branch_block_stmt_34/assign_stmt_728_to_assign_stmt_757/type_cast_743_Update/$entry
      -- CP-element group 123: 	 branch_block_stmt_34/assign_stmt_728_to_assign_stmt_757/type_cast_743_Update/cr
      -- CP-element group 123: 	 branch_block_stmt_34/forx_xcond144x_xpreheader_bbx_xnph231_PhiReq/$entry
      -- CP-element group 123: 	 branch_block_stmt_34/forx_xcond144x_xpreheader_bbx_xnph231_PhiReq/$exit
      -- CP-element group 123: 	 branch_block_stmt_34/merge_stmt_722_PhiReqMerge
      -- CP-element group 123: 	 branch_block_stmt_34/merge_stmt_722_PhiAck/$entry
      -- CP-element group 123: 	 branch_block_stmt_34/merge_stmt_722_PhiAck/$exit
      -- CP-element group 123: 	 branch_block_stmt_34/merge_stmt_722_PhiAck/dummy
      -- 
    if_choice_transition_1577_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_509_branch_ack_1, ack => testConfigure_CP_0_elements(123)); -- 
    rr_1953_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1953_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(123), ack => type_cast_743_inst_req_0); -- 
    cr_1958_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1958_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(123), ack => type_cast_743_inst_req_1); -- 
    -- CP-element group 124:  transition  place  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	265 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	278 
    -- CP-element group 124:  members (5) 
      -- CP-element group 124: 	 branch_block_stmt_34/if_stmt_509_else_link/$exit
      -- CP-element group 124: 	 branch_block_stmt_34/if_stmt_509_else_link/else_choice_transition
      -- CP-element group 124: 	 branch_block_stmt_34/forx_xcond144x_xpreheader_forx_xend204
      -- CP-element group 124: 	 branch_block_stmt_34/forx_xcond144x_xpreheader_forx_xend204_PhiReq/$entry
      -- CP-element group 124: 	 branch_block_stmt_34/forx_xcond144x_xpreheader_forx_xend204_PhiReq/$exit
      -- 
    else_choice_transition_1581_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_509_branch_ack_0, ack => testConfigure_CP_0_elements(124)); -- 
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	121 
    -- CP-element group 125: successors 
    -- CP-element group 125:  members (3) 
      -- CP-element group 125: 	 branch_block_stmt_34/assign_stmt_521_to_assign_stmt_550/type_cast_536_sample_completed_
      -- CP-element group 125: 	 branch_block_stmt_34/assign_stmt_521_to_assign_stmt_550/type_cast_536_Sample/$exit
      -- CP-element group 125: 	 branch_block_stmt_34/assign_stmt_521_to_assign_stmt_550/type_cast_536_Sample/ra
      -- 
    ra_1595_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_536_inst_ack_0, ack => testConfigure_CP_0_elements(125)); -- 
    -- CP-element group 126:  transition  place  input  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	121 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	266 
    -- CP-element group 126:  members (9) 
      -- CP-element group 126: 	 branch_block_stmt_34/assign_stmt_521_to_assign_stmt_550__exit__
      -- CP-element group 126: 	 branch_block_stmt_34/bbx_xnph235_forx_xbody90
      -- CP-element group 126: 	 branch_block_stmt_34/assign_stmt_521_to_assign_stmt_550/$exit
      -- CP-element group 126: 	 branch_block_stmt_34/assign_stmt_521_to_assign_stmt_550/type_cast_536_update_completed_
      -- CP-element group 126: 	 branch_block_stmt_34/assign_stmt_521_to_assign_stmt_550/type_cast_536_Update/$exit
      -- CP-element group 126: 	 branch_block_stmt_34/assign_stmt_521_to_assign_stmt_550/type_cast_536_Update/ca
      -- CP-element group 126: 	 branch_block_stmt_34/bbx_xnph235_forx_xbody90_PhiReq/$entry
      -- CP-element group 126: 	 branch_block_stmt_34/bbx_xnph235_forx_xbody90_PhiReq/phi_stmt_553/$entry
      -- CP-element group 126: 	 branch_block_stmt_34/bbx_xnph235_forx_xbody90_PhiReq/phi_stmt_553/phi_stmt_553_sources/$entry
      -- 
    ca_1600_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_536_inst_ack_1, ack => testConfigure_CP_0_elements(126)); -- 
    -- CP-element group 127:  transition  input  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	271 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	166 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/array_obj_ref_565_final_index_sum_regn_sample_complete
      -- CP-element group 127: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/array_obj_ref_565_final_index_sum_regn_Sample/$exit
      -- CP-element group 127: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/array_obj_ref_565_final_index_sum_regn_Sample/ack
      -- 
    ack_1629_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_565_index_offset_ack_0, ack => testConfigure_CP_0_elements(127)); -- 
    -- CP-element group 128:  transition  input  output  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	271 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	129 
    -- CP-element group 128:  members (11) 
      -- CP-element group 128: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/addr_of_566_sample_start_
      -- CP-element group 128: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/array_obj_ref_565_root_address_calculated
      -- CP-element group 128: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/array_obj_ref_565_offset_calculated
      -- CP-element group 128: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/array_obj_ref_565_final_index_sum_regn_Update/$exit
      -- CP-element group 128: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/array_obj_ref_565_final_index_sum_regn_Update/ack
      -- CP-element group 128: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/array_obj_ref_565_base_plus_offset/$entry
      -- CP-element group 128: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/array_obj_ref_565_base_plus_offset/$exit
      -- CP-element group 128: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/array_obj_ref_565_base_plus_offset/sum_rename_req
      -- CP-element group 128: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/array_obj_ref_565_base_plus_offset/sum_rename_ack
      -- CP-element group 128: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/addr_of_566_request/$entry
      -- CP-element group 128: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/addr_of_566_request/req
      -- 
    ack_1634_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_565_index_offset_ack_1, ack => testConfigure_CP_0_elements(128)); -- 
    req_1643_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1643_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(128), ack => addr_of_566_final_reg_req_0); -- 
    -- CP-element group 129:  transition  input  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	128 
    -- CP-element group 129: successors 
    -- CP-element group 129:  members (3) 
      -- CP-element group 129: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/addr_of_566_sample_completed_
      -- CP-element group 129: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/addr_of_566_request/$exit
      -- CP-element group 129: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/addr_of_566_request/ack
      -- 
    ack_1644_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_566_final_reg_ack_0, ack => testConfigure_CP_0_elements(129)); -- 
    -- CP-element group 130:  fork  transition  input  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	271 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	163 
    -- CP-element group 130:  members (19) 
      -- CP-element group 130: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/addr_of_566_update_completed_
      -- CP-element group 130: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/addr_of_566_complete/$exit
      -- CP-element group 130: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/addr_of_566_complete/ack
      -- CP-element group 130: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/ptr_deref_702_base_address_calculated
      -- CP-element group 130: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/ptr_deref_702_word_address_calculated
      -- CP-element group 130: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/ptr_deref_702_root_address_calculated
      -- CP-element group 130: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/ptr_deref_702_base_address_resized
      -- CP-element group 130: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/ptr_deref_702_base_addr_resize/$entry
      -- CP-element group 130: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/ptr_deref_702_base_addr_resize/$exit
      -- CP-element group 130: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/ptr_deref_702_base_addr_resize/base_resize_req
      -- CP-element group 130: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/ptr_deref_702_base_addr_resize/base_resize_ack
      -- CP-element group 130: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/ptr_deref_702_base_plus_offset/$entry
      -- CP-element group 130: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/ptr_deref_702_base_plus_offset/$exit
      -- CP-element group 130: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/ptr_deref_702_base_plus_offset/sum_rename_req
      -- CP-element group 130: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/ptr_deref_702_base_plus_offset/sum_rename_ack
      -- CP-element group 130: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/ptr_deref_702_word_addrgen/$entry
      -- CP-element group 130: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/ptr_deref_702_word_addrgen/$exit
      -- CP-element group 130: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/ptr_deref_702_word_addrgen/root_register_req
      -- CP-element group 130: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/ptr_deref_702_word_addrgen/root_register_ack
      -- 
    ack_1649_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_566_final_reg_ack_1, ack => testConfigure_CP_0_elements(130)); -- 
    -- CP-element group 131:  transition  input  output  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	271 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	132 
    -- CP-element group 131:  members (6) 
      -- CP-element group 131: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_569_sample_completed_
      -- CP-element group 131: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_569_update_start_
      -- CP-element group 131: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_569_Sample/$exit
      -- CP-element group 131: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_569_Sample/ra
      -- CP-element group 131: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_569_Update/$entry
      -- CP-element group 131: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_569_Update/cr
      -- 
    ra_1658_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_569_inst_ack_0, ack => testConfigure_CP_0_elements(131)); -- 
    cr_1662_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1662_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(131), ack => RPIPE_ConvTranspose_input_pipe_569_inst_req_1); -- 
    -- CP-element group 132:  fork  transition  input  output  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	131 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	133 
    -- CP-element group 132: 	135 
    -- CP-element group 132:  members (9) 
      -- CP-element group 132: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_569_update_completed_
      -- CP-element group 132: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_569_Update/$exit
      -- CP-element group 132: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_569_Update/ca
      -- CP-element group 132: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_573_sample_start_
      -- CP-element group 132: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_573_Sample/$entry
      -- CP-element group 132: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_573_Sample/rr
      -- CP-element group 132: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_582_sample_start_
      -- CP-element group 132: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_582_Sample/$entry
      -- CP-element group 132: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_582_Sample/rr
      -- 
    ca_1663_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_569_inst_ack_1, ack => testConfigure_CP_0_elements(132)); -- 
    rr_1671_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1671_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(132), ack => type_cast_573_inst_req_0); -- 
    rr_1685_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1685_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(132), ack => RPIPE_ConvTranspose_input_pipe_582_inst_req_0); -- 
    -- CP-element group 133:  transition  input  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	132 
    -- CP-element group 133: successors 
    -- CP-element group 133:  members (3) 
      -- CP-element group 133: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_573_sample_completed_
      -- CP-element group 133: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_573_Sample/$exit
      -- CP-element group 133: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_573_Sample/ra
      -- 
    ra_1672_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_573_inst_ack_0, ack => testConfigure_CP_0_elements(133)); -- 
    -- CP-element group 134:  transition  input  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	271 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	163 
    -- CP-element group 134:  members (3) 
      -- CP-element group 134: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_573_update_completed_
      -- CP-element group 134: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_573_Update/$exit
      -- CP-element group 134: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_573_Update/ca
      -- 
    ca_1677_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_573_inst_ack_1, ack => testConfigure_CP_0_elements(134)); -- 
    -- CP-element group 135:  transition  input  output  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	132 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	136 
    -- CP-element group 135:  members (6) 
      -- CP-element group 135: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_582_sample_completed_
      -- CP-element group 135: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_582_update_start_
      -- CP-element group 135: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_582_Sample/$exit
      -- CP-element group 135: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_582_Sample/ra
      -- CP-element group 135: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_582_Update/$entry
      -- CP-element group 135: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_582_Update/cr
      -- 
    ra_1686_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_582_inst_ack_0, ack => testConfigure_CP_0_elements(135)); -- 
    cr_1690_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1690_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(135), ack => RPIPE_ConvTranspose_input_pipe_582_inst_req_1); -- 
    -- CP-element group 136:  fork  transition  input  output  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	135 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	137 
    -- CP-element group 136: 	139 
    -- CP-element group 136:  members (9) 
      -- CP-element group 136: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_582_update_completed_
      -- CP-element group 136: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_582_Update/$exit
      -- CP-element group 136: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_582_Update/ca
      -- CP-element group 136: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_586_sample_start_
      -- CP-element group 136: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_586_Sample/$entry
      -- CP-element group 136: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_586_Sample/rr
      -- CP-element group 136: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_600_sample_start_
      -- CP-element group 136: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_600_Sample/$entry
      -- CP-element group 136: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_600_Sample/rr
      -- 
    ca_1691_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_582_inst_ack_1, ack => testConfigure_CP_0_elements(136)); -- 
    rr_1699_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1699_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(136), ack => type_cast_586_inst_req_0); -- 
    rr_1713_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1713_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(136), ack => RPIPE_ConvTranspose_input_pipe_600_inst_req_0); -- 
    -- CP-element group 137:  transition  input  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	136 
    -- CP-element group 137: successors 
    -- CP-element group 137:  members (3) 
      -- CP-element group 137: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_586_sample_completed_
      -- CP-element group 137: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_586_Sample/$exit
      -- CP-element group 137: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_586_Sample/ra
      -- 
    ra_1700_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_586_inst_ack_0, ack => testConfigure_CP_0_elements(137)); -- 
    -- CP-element group 138:  transition  input  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	271 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	163 
    -- CP-element group 138:  members (3) 
      -- CP-element group 138: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_586_update_completed_
      -- CP-element group 138: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_586_Update/$exit
      -- CP-element group 138: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_586_Update/ca
      -- 
    ca_1705_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_586_inst_ack_1, ack => testConfigure_CP_0_elements(138)); -- 
    -- CP-element group 139:  transition  input  output  bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	136 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	140 
    -- CP-element group 139:  members (6) 
      -- CP-element group 139: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_600_sample_completed_
      -- CP-element group 139: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_600_update_start_
      -- CP-element group 139: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_600_Sample/$exit
      -- CP-element group 139: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_600_Sample/ra
      -- CP-element group 139: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_600_Update/$entry
      -- CP-element group 139: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_600_Update/cr
      -- 
    ra_1714_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_600_inst_ack_0, ack => testConfigure_CP_0_elements(139)); -- 
    cr_1718_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1718_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(139), ack => RPIPE_ConvTranspose_input_pipe_600_inst_req_1); -- 
    -- CP-element group 140:  fork  transition  input  output  bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	139 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	141 
    -- CP-element group 140: 	143 
    -- CP-element group 140:  members (9) 
      -- CP-element group 140: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_600_update_completed_
      -- CP-element group 140: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_600_Update/$exit
      -- CP-element group 140: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_600_Update/ca
      -- CP-element group 140: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_604_sample_start_
      -- CP-element group 140: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_604_Sample/$entry
      -- CP-element group 140: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_604_Sample/rr
      -- CP-element group 140: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_618_sample_start_
      -- CP-element group 140: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_618_Sample/$entry
      -- CP-element group 140: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_618_Sample/rr
      -- 
    ca_1719_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_600_inst_ack_1, ack => testConfigure_CP_0_elements(140)); -- 
    rr_1727_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1727_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(140), ack => type_cast_604_inst_req_0); -- 
    rr_1741_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1741_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(140), ack => RPIPE_ConvTranspose_input_pipe_618_inst_req_0); -- 
    -- CP-element group 141:  transition  input  bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	140 
    -- CP-element group 141: successors 
    -- CP-element group 141:  members (3) 
      -- CP-element group 141: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_604_sample_completed_
      -- CP-element group 141: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_604_Sample/$exit
      -- CP-element group 141: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_604_Sample/ra
      -- 
    ra_1728_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_604_inst_ack_0, ack => testConfigure_CP_0_elements(141)); -- 
    -- CP-element group 142:  transition  input  bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	271 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	163 
    -- CP-element group 142:  members (3) 
      -- CP-element group 142: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_604_update_completed_
      -- CP-element group 142: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_604_Update/$exit
      -- CP-element group 142: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_604_Update/ca
      -- 
    ca_1733_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_604_inst_ack_1, ack => testConfigure_CP_0_elements(142)); -- 
    -- CP-element group 143:  transition  input  output  bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	140 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	144 
    -- CP-element group 143:  members (6) 
      -- CP-element group 143: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_618_sample_completed_
      -- CP-element group 143: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_618_update_start_
      -- CP-element group 143: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_618_Sample/$exit
      -- CP-element group 143: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_618_Sample/ra
      -- CP-element group 143: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_618_Update/$entry
      -- CP-element group 143: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_618_Update/cr
      -- 
    ra_1742_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_618_inst_ack_0, ack => testConfigure_CP_0_elements(143)); -- 
    cr_1746_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1746_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(143), ack => RPIPE_ConvTranspose_input_pipe_618_inst_req_1); -- 
    -- CP-element group 144:  fork  transition  input  output  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	143 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	145 
    -- CP-element group 144: 	147 
    -- CP-element group 144:  members (9) 
      -- CP-element group 144: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_618_update_completed_
      -- CP-element group 144: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_618_Update/$exit
      -- CP-element group 144: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_618_Update/ca
      -- CP-element group 144: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_622_sample_start_
      -- CP-element group 144: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_622_Sample/$entry
      -- CP-element group 144: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_622_Sample/rr
      -- CP-element group 144: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_636_sample_start_
      -- CP-element group 144: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_636_Sample/$entry
      -- CP-element group 144: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_636_Sample/rr
      -- 
    ca_1747_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_618_inst_ack_1, ack => testConfigure_CP_0_elements(144)); -- 
    rr_1755_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1755_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(144), ack => type_cast_622_inst_req_0); -- 
    rr_1769_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1769_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(144), ack => RPIPE_ConvTranspose_input_pipe_636_inst_req_0); -- 
    -- CP-element group 145:  transition  input  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	144 
    -- CP-element group 145: successors 
    -- CP-element group 145:  members (3) 
      -- CP-element group 145: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_622_sample_completed_
      -- CP-element group 145: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_622_Sample/$exit
      -- CP-element group 145: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_622_Sample/ra
      -- 
    ra_1756_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_622_inst_ack_0, ack => testConfigure_CP_0_elements(145)); -- 
    -- CP-element group 146:  transition  input  bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	271 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	163 
    -- CP-element group 146:  members (3) 
      -- CP-element group 146: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_622_update_completed_
      -- CP-element group 146: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_622_Update/$exit
      -- CP-element group 146: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_622_Update/ca
      -- 
    ca_1761_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_622_inst_ack_1, ack => testConfigure_CP_0_elements(146)); -- 
    -- CP-element group 147:  transition  input  output  bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	144 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	148 
    -- CP-element group 147:  members (6) 
      -- CP-element group 147: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_636_sample_completed_
      -- CP-element group 147: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_636_update_start_
      -- CP-element group 147: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_636_Sample/$exit
      -- CP-element group 147: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_636_Sample/ra
      -- CP-element group 147: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_636_Update/$entry
      -- CP-element group 147: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_636_Update/cr
      -- 
    ra_1770_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_636_inst_ack_0, ack => testConfigure_CP_0_elements(147)); -- 
    cr_1774_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1774_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(147), ack => RPIPE_ConvTranspose_input_pipe_636_inst_req_1); -- 
    -- CP-element group 148:  fork  transition  input  output  bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	147 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	149 
    -- CP-element group 148: 	151 
    -- CP-element group 148:  members (9) 
      -- CP-element group 148: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_636_update_completed_
      -- CP-element group 148: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_636_Update/$exit
      -- CP-element group 148: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_636_Update/ca
      -- CP-element group 148: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_640_sample_start_
      -- CP-element group 148: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_640_Sample/$entry
      -- CP-element group 148: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_640_Sample/rr
      -- CP-element group 148: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_654_sample_start_
      -- CP-element group 148: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_654_Sample/$entry
      -- CP-element group 148: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_654_Sample/rr
      -- 
    ca_1775_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_636_inst_ack_1, ack => testConfigure_CP_0_elements(148)); -- 
    rr_1783_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1783_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(148), ack => type_cast_640_inst_req_0); -- 
    rr_1797_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1797_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(148), ack => RPIPE_ConvTranspose_input_pipe_654_inst_req_0); -- 
    -- CP-element group 149:  transition  input  bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	148 
    -- CP-element group 149: successors 
    -- CP-element group 149:  members (3) 
      -- CP-element group 149: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_640_sample_completed_
      -- CP-element group 149: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_640_Sample/$exit
      -- CP-element group 149: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_640_Sample/ra
      -- 
    ra_1784_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_640_inst_ack_0, ack => testConfigure_CP_0_elements(149)); -- 
    -- CP-element group 150:  transition  input  bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	271 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	163 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_640_update_completed_
      -- CP-element group 150: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_640_Update/$exit
      -- CP-element group 150: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_640_Update/ca
      -- 
    ca_1789_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_640_inst_ack_1, ack => testConfigure_CP_0_elements(150)); -- 
    -- CP-element group 151:  transition  input  output  bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	148 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	152 
    -- CP-element group 151:  members (6) 
      -- CP-element group 151: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_654_sample_completed_
      -- CP-element group 151: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_654_update_start_
      -- CP-element group 151: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_654_Sample/$exit
      -- CP-element group 151: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_654_Sample/ra
      -- CP-element group 151: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_654_Update/$entry
      -- CP-element group 151: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_654_Update/cr
      -- 
    ra_1798_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_654_inst_ack_0, ack => testConfigure_CP_0_elements(151)); -- 
    cr_1802_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1802_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(151), ack => RPIPE_ConvTranspose_input_pipe_654_inst_req_1); -- 
    -- CP-element group 152:  fork  transition  input  output  bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	151 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	153 
    -- CP-element group 152: 	155 
    -- CP-element group 152:  members (9) 
      -- CP-element group 152: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_654_update_completed_
      -- CP-element group 152: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_654_Update/$exit
      -- CP-element group 152: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_654_Update/ca
      -- CP-element group 152: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_658_sample_start_
      -- CP-element group 152: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_658_Sample/$entry
      -- CP-element group 152: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_658_Sample/rr
      -- CP-element group 152: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_672_sample_start_
      -- CP-element group 152: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_672_Sample/$entry
      -- CP-element group 152: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_672_Sample/rr
      -- 
    ca_1803_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_654_inst_ack_1, ack => testConfigure_CP_0_elements(152)); -- 
    rr_1811_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1811_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(152), ack => type_cast_658_inst_req_0); -- 
    rr_1825_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1825_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(152), ack => RPIPE_ConvTranspose_input_pipe_672_inst_req_0); -- 
    -- CP-element group 153:  transition  input  bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	152 
    -- CP-element group 153: successors 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_658_sample_completed_
      -- CP-element group 153: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_658_Sample/$exit
      -- CP-element group 153: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_658_Sample/ra
      -- 
    ra_1812_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_658_inst_ack_0, ack => testConfigure_CP_0_elements(153)); -- 
    -- CP-element group 154:  transition  input  bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	271 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	163 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_658_update_completed_
      -- CP-element group 154: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_658_Update/$exit
      -- CP-element group 154: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_658_Update/ca
      -- 
    ca_1817_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_658_inst_ack_1, ack => testConfigure_CP_0_elements(154)); -- 
    -- CP-element group 155:  transition  input  output  bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	152 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	156 
    -- CP-element group 155:  members (6) 
      -- CP-element group 155: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_672_sample_completed_
      -- CP-element group 155: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_672_update_start_
      -- CP-element group 155: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_672_Sample/$exit
      -- CP-element group 155: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_672_Sample/ra
      -- CP-element group 155: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_672_Update/$entry
      -- CP-element group 155: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_672_Update/cr
      -- 
    ra_1826_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_672_inst_ack_0, ack => testConfigure_CP_0_elements(155)); -- 
    cr_1830_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1830_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(155), ack => RPIPE_ConvTranspose_input_pipe_672_inst_req_1); -- 
    -- CP-element group 156:  fork  transition  input  output  bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	155 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	157 
    -- CP-element group 156: 	159 
    -- CP-element group 156:  members (9) 
      -- CP-element group 156: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_672_update_completed_
      -- CP-element group 156: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_672_Update/$exit
      -- CP-element group 156: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_672_Update/ca
      -- CP-element group 156: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_676_sample_start_
      -- CP-element group 156: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_676_Sample/$entry
      -- CP-element group 156: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_676_Sample/rr
      -- CP-element group 156: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_690_sample_start_
      -- CP-element group 156: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_690_Sample/$entry
      -- CP-element group 156: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_690_Sample/rr
      -- 
    ca_1831_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_672_inst_ack_1, ack => testConfigure_CP_0_elements(156)); -- 
    rr_1839_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1839_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(156), ack => type_cast_676_inst_req_0); -- 
    rr_1853_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1853_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(156), ack => RPIPE_ConvTranspose_input_pipe_690_inst_req_0); -- 
    -- CP-element group 157:  transition  input  bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	156 
    -- CP-element group 157: successors 
    -- CP-element group 157:  members (3) 
      -- CP-element group 157: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_676_sample_completed_
      -- CP-element group 157: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_676_Sample/$exit
      -- CP-element group 157: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_676_Sample/ra
      -- 
    ra_1840_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_676_inst_ack_0, ack => testConfigure_CP_0_elements(157)); -- 
    -- CP-element group 158:  transition  input  bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	271 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	163 
    -- CP-element group 158:  members (3) 
      -- CP-element group 158: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_676_update_completed_
      -- CP-element group 158: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_676_Update/$exit
      -- CP-element group 158: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_676_Update/ca
      -- 
    ca_1845_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_676_inst_ack_1, ack => testConfigure_CP_0_elements(158)); -- 
    -- CP-element group 159:  transition  input  output  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	156 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	160 
    -- CP-element group 159:  members (6) 
      -- CP-element group 159: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_690_sample_completed_
      -- CP-element group 159: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_690_update_start_
      -- CP-element group 159: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_690_Sample/$exit
      -- CP-element group 159: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_690_Sample/ra
      -- CP-element group 159: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_690_Update/$entry
      -- CP-element group 159: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_690_Update/cr
      -- 
    ra_1854_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_690_inst_ack_0, ack => testConfigure_CP_0_elements(159)); -- 
    cr_1858_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1858_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(159), ack => RPIPE_ConvTranspose_input_pipe_690_inst_req_1); -- 
    -- CP-element group 160:  transition  input  output  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	159 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	161 
    -- CP-element group 160:  members (6) 
      -- CP-element group 160: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_690_update_completed_
      -- CP-element group 160: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_690_Update/$exit
      -- CP-element group 160: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_690_Update/ca
      -- CP-element group 160: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_694_sample_start_
      -- CP-element group 160: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_694_Sample/$entry
      -- CP-element group 160: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_694_Sample/rr
      -- 
    ca_1859_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_690_inst_ack_1, ack => testConfigure_CP_0_elements(160)); -- 
    rr_1867_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1867_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(160), ack => type_cast_694_inst_req_0); -- 
    -- CP-element group 161:  transition  input  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	160 
    -- CP-element group 161: successors 
    -- CP-element group 161:  members (3) 
      -- CP-element group 161: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_694_sample_completed_
      -- CP-element group 161: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_694_Sample/$exit
      -- CP-element group 161: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_694_Sample/ra
      -- 
    ra_1868_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_694_inst_ack_0, ack => testConfigure_CP_0_elements(161)); -- 
    -- CP-element group 162:  transition  input  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	271 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	163 
    -- CP-element group 162:  members (3) 
      -- CP-element group 162: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_694_update_completed_
      -- CP-element group 162: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_694_Update/$exit
      -- CP-element group 162: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_694_Update/ca
      -- 
    ca_1873_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_694_inst_ack_1, ack => testConfigure_CP_0_elements(162)); -- 
    -- CP-element group 163:  join  transition  output  bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	130 
    -- CP-element group 163: 	134 
    -- CP-element group 163: 	138 
    -- CP-element group 163: 	142 
    -- CP-element group 163: 	146 
    -- CP-element group 163: 	150 
    -- CP-element group 163: 	154 
    -- CP-element group 163: 	158 
    -- CP-element group 163: 	162 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	164 
    -- CP-element group 163:  members (9) 
      -- CP-element group 163: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/ptr_deref_702_sample_start_
      -- CP-element group 163: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/ptr_deref_702_Sample/$entry
      -- CP-element group 163: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/ptr_deref_702_Sample/ptr_deref_702_Split/$entry
      -- CP-element group 163: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/ptr_deref_702_Sample/ptr_deref_702_Split/$exit
      -- CP-element group 163: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/ptr_deref_702_Sample/ptr_deref_702_Split/split_req
      -- CP-element group 163: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/ptr_deref_702_Sample/ptr_deref_702_Split/split_ack
      -- CP-element group 163: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/ptr_deref_702_Sample/word_access_start/$entry
      -- CP-element group 163: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/ptr_deref_702_Sample/word_access_start/word_0/$entry
      -- CP-element group 163: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/ptr_deref_702_Sample/word_access_start/word_0/rr
      -- 
    rr_1911_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1911_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(163), ack => ptr_deref_702_store_0_req_0); -- 
    testConfigure_cp_element_group_163: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_163"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(130) & testConfigure_CP_0_elements(134) & testConfigure_CP_0_elements(138) & testConfigure_CP_0_elements(142) & testConfigure_CP_0_elements(146) & testConfigure_CP_0_elements(150) & testConfigure_CP_0_elements(154) & testConfigure_CP_0_elements(158) & testConfigure_CP_0_elements(162);
      gj_testConfigure_cp_element_group_163 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(163), clk => clk, reset => reset); --
    end block;
    -- CP-element group 164:  transition  input  bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	163 
    -- CP-element group 164: successors 
    -- CP-element group 164:  members (5) 
      -- CP-element group 164: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/ptr_deref_702_sample_completed_
      -- CP-element group 164: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/ptr_deref_702_Sample/$exit
      -- CP-element group 164: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/ptr_deref_702_Sample/word_access_start/$exit
      -- CP-element group 164: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/ptr_deref_702_Sample/word_access_start/word_0/$exit
      -- CP-element group 164: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/ptr_deref_702_Sample/word_access_start/word_0/ra
      -- 
    ra_1912_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_702_store_0_ack_0, ack => testConfigure_CP_0_elements(164)); -- 
    -- CP-element group 165:  transition  input  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	271 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	166 
    -- CP-element group 165:  members (5) 
      -- CP-element group 165: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/ptr_deref_702_update_completed_
      -- CP-element group 165: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/ptr_deref_702_Update/$exit
      -- CP-element group 165: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/ptr_deref_702_Update/word_access_complete/$exit
      -- CP-element group 165: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/ptr_deref_702_Update/word_access_complete/word_0/$exit
      -- CP-element group 165: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/ptr_deref_702_Update/word_access_complete/word_0/ca
      -- 
    ca_1923_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_702_store_0_ack_1, ack => testConfigure_CP_0_elements(165)); -- 
    -- CP-element group 166:  branch  join  transition  place  output  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	127 
    -- CP-element group 166: 	165 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	167 
    -- CP-element group 166: 	168 
    -- CP-element group 166:  members (10) 
      -- CP-element group 166: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715__exit__
      -- CP-element group 166: 	 branch_block_stmt_34/if_stmt_716__entry__
      -- CP-element group 166: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/$exit
      -- CP-element group 166: 	 branch_block_stmt_34/if_stmt_716_dead_link/$entry
      -- CP-element group 166: 	 branch_block_stmt_34/if_stmt_716_eval_test/$entry
      -- CP-element group 166: 	 branch_block_stmt_34/if_stmt_716_eval_test/$exit
      -- CP-element group 166: 	 branch_block_stmt_34/if_stmt_716_eval_test/branch_req
      -- CP-element group 166: 	 branch_block_stmt_34/R_exitcond2_717_place
      -- CP-element group 166: 	 branch_block_stmt_34/if_stmt_716_if_link/$entry
      -- CP-element group 166: 	 branch_block_stmt_34/if_stmt_716_else_link/$entry
      -- 
    branch_req_1931_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1931_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(166), ack => if_stmt_716_branch_req_0); -- 
    testConfigure_cp_element_group_166: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_166"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(127) & testConfigure_CP_0_elements(165);
      gj_testConfigure_cp_element_group_166 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(166), clk => clk, reset => reset); --
    end block;
    -- CP-element group 167:  merge  transition  place  input  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	166 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	265 
    -- CP-element group 167:  members (13) 
      -- CP-element group 167: 	 branch_block_stmt_34/merge_stmt_500__exit__
      -- CP-element group 167: 	 branch_block_stmt_34/forx_xcond144x_xpreheaderx_xloopexit_forx_xcond144x_xpreheader
      -- CP-element group 167: 	 branch_block_stmt_34/if_stmt_716_if_link/$exit
      -- CP-element group 167: 	 branch_block_stmt_34/if_stmt_716_if_link/if_choice_transition
      -- CP-element group 167: 	 branch_block_stmt_34/forx_xbody90_forx_xcond144x_xpreheaderx_xloopexit
      -- CP-element group 167: 	 branch_block_stmt_34/forx_xbody90_forx_xcond144x_xpreheaderx_xloopexit_PhiReq/$entry
      -- CP-element group 167: 	 branch_block_stmt_34/forx_xbody90_forx_xcond144x_xpreheaderx_xloopexit_PhiReq/$exit
      -- CP-element group 167: 	 branch_block_stmt_34/merge_stmt_500_PhiReqMerge
      -- CP-element group 167: 	 branch_block_stmt_34/merge_stmt_500_PhiAck/$entry
      -- CP-element group 167: 	 branch_block_stmt_34/merge_stmt_500_PhiAck/$exit
      -- CP-element group 167: 	 branch_block_stmt_34/merge_stmt_500_PhiAck/dummy
      -- CP-element group 167: 	 branch_block_stmt_34/forx_xcond144x_xpreheaderx_xloopexit_forx_xcond144x_xpreheader_PhiReq/$entry
      -- CP-element group 167: 	 branch_block_stmt_34/forx_xcond144x_xpreheaderx_xloopexit_forx_xcond144x_xpreheader_PhiReq/$exit
      -- 
    if_choice_transition_1936_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_716_branch_ack_1, ack => testConfigure_CP_0_elements(167)); -- 
    -- CP-element group 168:  fork  transition  place  input  output  bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	166 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	267 
    -- CP-element group 168: 	268 
    -- CP-element group 168:  members (12) 
      -- CP-element group 168: 	 branch_block_stmt_34/if_stmt_716_else_link/$exit
      -- CP-element group 168: 	 branch_block_stmt_34/if_stmt_716_else_link/else_choice_transition
      -- CP-element group 168: 	 branch_block_stmt_34/forx_xbody90_forx_xbody90
      -- CP-element group 168: 	 branch_block_stmt_34/forx_xbody90_forx_xbody90_PhiReq/$entry
      -- CP-element group 168: 	 branch_block_stmt_34/forx_xbody90_forx_xbody90_PhiReq/phi_stmt_553/$entry
      -- CP-element group 168: 	 branch_block_stmt_34/forx_xbody90_forx_xbody90_PhiReq/phi_stmt_553/phi_stmt_553_sources/$entry
      -- CP-element group 168: 	 branch_block_stmt_34/forx_xbody90_forx_xbody90_PhiReq/phi_stmt_553/phi_stmt_553_sources/type_cast_559/$entry
      -- CP-element group 168: 	 branch_block_stmt_34/forx_xbody90_forx_xbody90_PhiReq/phi_stmt_553/phi_stmt_553_sources/type_cast_559/SplitProtocol/$entry
      -- CP-element group 168: 	 branch_block_stmt_34/forx_xbody90_forx_xbody90_PhiReq/phi_stmt_553/phi_stmt_553_sources/type_cast_559/SplitProtocol/Sample/$entry
      -- CP-element group 168: 	 branch_block_stmt_34/forx_xbody90_forx_xbody90_PhiReq/phi_stmt_553/phi_stmt_553_sources/type_cast_559/SplitProtocol/Sample/rr
      -- CP-element group 168: 	 branch_block_stmt_34/forx_xbody90_forx_xbody90_PhiReq/phi_stmt_553/phi_stmt_553_sources/type_cast_559/SplitProtocol/Update/$entry
      -- CP-element group 168: 	 branch_block_stmt_34/forx_xbody90_forx_xbody90_PhiReq/phi_stmt_553/phi_stmt_553_sources/type_cast_559/SplitProtocol/Update/cr
      -- 
    else_choice_transition_1940_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_716_branch_ack_0, ack => testConfigure_CP_0_elements(168)); -- 
    rr_2908_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2908_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(168), ack => type_cast_559_inst_req_0); -- 
    cr_2913_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2913_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(168), ack => type_cast_559_inst_req_1); -- 
    -- CP-element group 169:  transition  input  bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	123 
    -- CP-element group 169: successors 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_34/assign_stmt_728_to_assign_stmt_757/type_cast_743_sample_completed_
      -- CP-element group 169: 	 branch_block_stmt_34/assign_stmt_728_to_assign_stmt_757/type_cast_743_Sample/$exit
      -- CP-element group 169: 	 branch_block_stmt_34/assign_stmt_728_to_assign_stmt_757/type_cast_743_Sample/ra
      -- 
    ra_1954_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_743_inst_ack_0, ack => testConfigure_CP_0_elements(169)); -- 
    -- CP-element group 170:  transition  place  input  bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	123 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	272 
    -- CP-element group 170:  members (9) 
      -- CP-element group 170: 	 branch_block_stmt_34/assign_stmt_728_to_assign_stmt_757__exit__
      -- CP-element group 170: 	 branch_block_stmt_34/bbx_xnph231_forx_xbody150
      -- CP-element group 170: 	 branch_block_stmt_34/assign_stmt_728_to_assign_stmt_757/$exit
      -- CP-element group 170: 	 branch_block_stmt_34/assign_stmt_728_to_assign_stmt_757/type_cast_743_update_completed_
      -- CP-element group 170: 	 branch_block_stmt_34/assign_stmt_728_to_assign_stmt_757/type_cast_743_Update/$exit
      -- CP-element group 170: 	 branch_block_stmt_34/assign_stmt_728_to_assign_stmt_757/type_cast_743_Update/ca
      -- CP-element group 170: 	 branch_block_stmt_34/bbx_xnph231_forx_xbody150_PhiReq/$entry
      -- CP-element group 170: 	 branch_block_stmt_34/bbx_xnph231_forx_xbody150_PhiReq/phi_stmt_760/$entry
      -- CP-element group 170: 	 branch_block_stmt_34/bbx_xnph231_forx_xbody150_PhiReq/phi_stmt_760/phi_stmt_760_sources/$entry
      -- 
    ca_1959_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_743_inst_ack_1, ack => testConfigure_CP_0_elements(170)); -- 
    -- CP-element group 171:  transition  input  bypass 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	277 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	210 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/array_obj_ref_772_final_index_sum_regn_sample_complete
      -- CP-element group 171: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/array_obj_ref_772_final_index_sum_regn_Sample/$exit
      -- CP-element group 171: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/array_obj_ref_772_final_index_sum_regn_Sample/ack
      -- 
    ack_1988_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_772_index_offset_ack_0, ack => testConfigure_CP_0_elements(171)); -- 
    -- CP-element group 172:  transition  input  output  bypass 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	277 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	173 
    -- CP-element group 172:  members (11) 
      -- CP-element group 172: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/addr_of_773_sample_start_
      -- CP-element group 172: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/array_obj_ref_772_root_address_calculated
      -- CP-element group 172: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/array_obj_ref_772_offset_calculated
      -- CP-element group 172: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/array_obj_ref_772_final_index_sum_regn_Update/$exit
      -- CP-element group 172: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/array_obj_ref_772_final_index_sum_regn_Update/ack
      -- CP-element group 172: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/array_obj_ref_772_base_plus_offset/$entry
      -- CP-element group 172: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/array_obj_ref_772_base_plus_offset/$exit
      -- CP-element group 172: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/array_obj_ref_772_base_plus_offset/sum_rename_req
      -- CP-element group 172: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/array_obj_ref_772_base_plus_offset/sum_rename_ack
      -- CP-element group 172: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/addr_of_773_request/$entry
      -- CP-element group 172: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/addr_of_773_request/req
      -- 
    ack_1993_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_772_index_offset_ack_1, ack => testConfigure_CP_0_elements(172)); -- 
    req_2002_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2002_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(172), ack => addr_of_773_final_reg_req_0); -- 
    -- CP-element group 173:  transition  input  bypass 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	172 
    -- CP-element group 173: successors 
    -- CP-element group 173:  members (3) 
      -- CP-element group 173: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/addr_of_773_sample_completed_
      -- CP-element group 173: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/addr_of_773_request/$exit
      -- CP-element group 173: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/addr_of_773_request/ack
      -- 
    ack_2003_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_773_final_reg_ack_0, ack => testConfigure_CP_0_elements(173)); -- 
    -- CP-element group 174:  fork  transition  input  bypass 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	277 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	207 
    -- CP-element group 174:  members (19) 
      -- CP-element group 174: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/ptr_deref_909_root_address_calculated
      -- CP-element group 174: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/ptr_deref_909_base_address_resized
      -- CP-element group 174: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/ptr_deref_909_base_addr_resize/$entry
      -- CP-element group 174: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/ptr_deref_909_base_address_calculated
      -- CP-element group 174: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/ptr_deref_909_word_address_calculated
      -- CP-element group 174: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/ptr_deref_909_word_addrgen/root_register_ack
      -- CP-element group 174: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/ptr_deref_909_word_addrgen/root_register_req
      -- CP-element group 174: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/ptr_deref_909_word_addrgen/$exit
      -- CP-element group 174: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/ptr_deref_909_word_addrgen/$entry
      -- CP-element group 174: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/ptr_deref_909_base_plus_offset/sum_rename_ack
      -- CP-element group 174: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/ptr_deref_909_base_plus_offset/sum_rename_req
      -- CP-element group 174: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/ptr_deref_909_base_plus_offset/$exit
      -- CP-element group 174: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/ptr_deref_909_base_plus_offset/$entry
      -- CP-element group 174: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/ptr_deref_909_base_addr_resize/base_resize_ack
      -- CP-element group 174: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/ptr_deref_909_base_addr_resize/base_resize_req
      -- CP-element group 174: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/ptr_deref_909_base_addr_resize/$exit
      -- CP-element group 174: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/addr_of_773_update_completed_
      -- CP-element group 174: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/addr_of_773_complete/$exit
      -- CP-element group 174: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/addr_of_773_complete/ack
      -- 
    ack_2008_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_773_final_reg_ack_1, ack => testConfigure_CP_0_elements(174)); -- 
    -- CP-element group 175:  transition  input  output  bypass 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	277 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	176 
    -- CP-element group 175:  members (6) 
      -- CP-element group 175: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_776_sample_completed_
      -- CP-element group 175: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_776_update_start_
      -- CP-element group 175: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_776_Sample/$exit
      -- CP-element group 175: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_776_Sample/ra
      -- CP-element group 175: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_776_Update/$entry
      -- CP-element group 175: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_776_Update/cr
      -- 
    ra_2017_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_776_inst_ack_0, ack => testConfigure_CP_0_elements(175)); -- 
    cr_2021_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2021_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(175), ack => RPIPE_ConvTranspose_input_pipe_776_inst_req_1); -- 
    -- CP-element group 176:  fork  transition  input  output  bypass 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	175 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	177 
    -- CP-element group 176: 	179 
    -- CP-element group 176:  members (9) 
      -- CP-element group 176: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_776_update_completed_
      -- CP-element group 176: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_776_Update/$exit
      -- CP-element group 176: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_776_Update/ca
      -- CP-element group 176: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_780_sample_start_
      -- CP-element group 176: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_780_Sample/$entry
      -- CP-element group 176: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_780_Sample/rr
      -- CP-element group 176: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_789_sample_start_
      -- CP-element group 176: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_789_Sample/$entry
      -- CP-element group 176: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_789_Sample/rr
      -- 
    ca_2022_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_776_inst_ack_1, ack => testConfigure_CP_0_elements(176)); -- 
    rr_2030_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2030_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(176), ack => type_cast_780_inst_req_0); -- 
    rr_2044_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2044_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(176), ack => RPIPE_ConvTranspose_input_pipe_789_inst_req_0); -- 
    -- CP-element group 177:  transition  input  bypass 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	176 
    -- CP-element group 177: successors 
    -- CP-element group 177:  members (3) 
      -- CP-element group 177: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_780_sample_completed_
      -- CP-element group 177: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_780_Sample/$exit
      -- CP-element group 177: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_780_Sample/ra
      -- 
    ra_2031_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_780_inst_ack_0, ack => testConfigure_CP_0_elements(177)); -- 
    -- CP-element group 178:  transition  input  bypass 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	277 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	207 
    -- CP-element group 178:  members (3) 
      -- CP-element group 178: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_780_update_completed_
      -- CP-element group 178: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_780_Update/$exit
      -- CP-element group 178: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_780_Update/ca
      -- 
    ca_2036_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_780_inst_ack_1, ack => testConfigure_CP_0_elements(178)); -- 
    -- CP-element group 179:  transition  input  output  bypass 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	176 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	180 
    -- CP-element group 179:  members (6) 
      -- CP-element group 179: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_789_sample_completed_
      -- CP-element group 179: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_789_update_start_
      -- CP-element group 179: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_789_Sample/$exit
      -- CP-element group 179: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_789_Sample/ra
      -- CP-element group 179: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_789_Update/$entry
      -- CP-element group 179: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_789_Update/cr
      -- 
    ra_2045_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_789_inst_ack_0, ack => testConfigure_CP_0_elements(179)); -- 
    cr_2049_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2049_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(179), ack => RPIPE_ConvTranspose_input_pipe_789_inst_req_1); -- 
    -- CP-element group 180:  fork  transition  input  output  bypass 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	179 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	181 
    -- CP-element group 180: 	183 
    -- CP-element group 180:  members (9) 
      -- CP-element group 180: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_789_update_completed_
      -- CP-element group 180: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_789_Update/$exit
      -- CP-element group 180: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_789_Update/ca
      -- CP-element group 180: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_793_sample_start_
      -- CP-element group 180: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_793_Sample/$entry
      -- CP-element group 180: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_793_Sample/rr
      -- CP-element group 180: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_807_sample_start_
      -- CP-element group 180: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_807_Sample/$entry
      -- CP-element group 180: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_807_Sample/rr
      -- 
    ca_2050_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_789_inst_ack_1, ack => testConfigure_CP_0_elements(180)); -- 
    rr_2058_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2058_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(180), ack => type_cast_793_inst_req_0); -- 
    rr_2072_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2072_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(180), ack => RPIPE_ConvTranspose_input_pipe_807_inst_req_0); -- 
    -- CP-element group 181:  transition  input  bypass 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	180 
    -- CP-element group 181: successors 
    -- CP-element group 181:  members (3) 
      -- CP-element group 181: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_793_sample_completed_
      -- CP-element group 181: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_793_Sample/$exit
      -- CP-element group 181: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_793_Sample/ra
      -- 
    ra_2059_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_793_inst_ack_0, ack => testConfigure_CP_0_elements(181)); -- 
    -- CP-element group 182:  transition  input  bypass 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	277 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	207 
    -- CP-element group 182:  members (3) 
      -- CP-element group 182: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_793_update_completed_
      -- CP-element group 182: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_793_Update/$exit
      -- CP-element group 182: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_793_Update/ca
      -- 
    ca_2064_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_793_inst_ack_1, ack => testConfigure_CP_0_elements(182)); -- 
    -- CP-element group 183:  transition  input  output  bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	180 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	184 
    -- CP-element group 183:  members (6) 
      -- CP-element group 183: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_807_sample_completed_
      -- CP-element group 183: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_807_update_start_
      -- CP-element group 183: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_807_Sample/$exit
      -- CP-element group 183: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_807_Sample/ra
      -- CP-element group 183: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_807_Update/$entry
      -- CP-element group 183: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_807_Update/cr
      -- 
    ra_2073_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_807_inst_ack_0, ack => testConfigure_CP_0_elements(183)); -- 
    cr_2077_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2077_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(183), ack => RPIPE_ConvTranspose_input_pipe_807_inst_req_1); -- 
    -- CP-element group 184:  fork  transition  input  output  bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	183 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	185 
    -- CP-element group 184: 	187 
    -- CP-element group 184:  members (9) 
      -- CP-element group 184: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_807_update_completed_
      -- CP-element group 184: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_807_Update/$exit
      -- CP-element group 184: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_807_Update/ca
      -- CP-element group 184: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_811_sample_start_
      -- CP-element group 184: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_811_Sample/$entry
      -- CP-element group 184: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_811_Sample/rr
      -- CP-element group 184: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_825_sample_start_
      -- CP-element group 184: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_825_Sample/$entry
      -- CP-element group 184: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_825_Sample/rr
      -- 
    ca_2078_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_807_inst_ack_1, ack => testConfigure_CP_0_elements(184)); -- 
    rr_2086_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2086_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(184), ack => type_cast_811_inst_req_0); -- 
    rr_2100_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2100_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(184), ack => RPIPE_ConvTranspose_input_pipe_825_inst_req_0); -- 
    -- CP-element group 185:  transition  input  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	184 
    -- CP-element group 185: successors 
    -- CP-element group 185:  members (3) 
      -- CP-element group 185: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_811_sample_completed_
      -- CP-element group 185: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_811_Sample/$exit
      -- CP-element group 185: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_811_Sample/ra
      -- 
    ra_2087_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_811_inst_ack_0, ack => testConfigure_CP_0_elements(185)); -- 
    -- CP-element group 186:  transition  input  bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	277 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	207 
    -- CP-element group 186:  members (3) 
      -- CP-element group 186: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_811_update_completed_
      -- CP-element group 186: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_811_Update/$exit
      -- CP-element group 186: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_811_Update/ca
      -- 
    ca_2092_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_811_inst_ack_1, ack => testConfigure_CP_0_elements(186)); -- 
    -- CP-element group 187:  transition  input  output  bypass 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	184 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	188 
    -- CP-element group 187:  members (6) 
      -- CP-element group 187: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_825_sample_completed_
      -- CP-element group 187: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_825_update_start_
      -- CP-element group 187: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_825_Sample/$exit
      -- CP-element group 187: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_825_Sample/ra
      -- CP-element group 187: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_825_Update/$entry
      -- CP-element group 187: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_825_Update/cr
      -- 
    ra_2101_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_825_inst_ack_0, ack => testConfigure_CP_0_elements(187)); -- 
    cr_2105_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2105_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(187), ack => RPIPE_ConvTranspose_input_pipe_825_inst_req_1); -- 
    -- CP-element group 188:  fork  transition  input  output  bypass 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	187 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	189 
    -- CP-element group 188: 	191 
    -- CP-element group 188:  members (9) 
      -- CP-element group 188: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_843_Sample/$entry
      -- CP-element group 188: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_843_Sample/rr
      -- CP-element group 188: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_843_sample_start_
      -- CP-element group 188: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_825_update_completed_
      -- CP-element group 188: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_825_Update/$exit
      -- CP-element group 188: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_825_Update/ca
      -- CP-element group 188: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_829_sample_start_
      -- CP-element group 188: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_829_Sample/$entry
      -- CP-element group 188: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_829_Sample/rr
      -- 
    ca_2106_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_825_inst_ack_1, ack => testConfigure_CP_0_elements(188)); -- 
    rr_2114_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2114_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(188), ack => type_cast_829_inst_req_0); -- 
    rr_2128_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2128_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(188), ack => RPIPE_ConvTranspose_input_pipe_843_inst_req_0); -- 
    -- CP-element group 189:  transition  input  bypass 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	188 
    -- CP-element group 189: successors 
    -- CP-element group 189:  members (3) 
      -- CP-element group 189: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_829_sample_completed_
      -- CP-element group 189: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_829_Sample/$exit
      -- CP-element group 189: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_829_Sample/ra
      -- 
    ra_2115_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_829_inst_ack_0, ack => testConfigure_CP_0_elements(189)); -- 
    -- CP-element group 190:  transition  input  bypass 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	277 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	207 
    -- CP-element group 190:  members (3) 
      -- CP-element group 190: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_829_Update/ca
      -- CP-element group 190: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_829_Update/$exit
      -- CP-element group 190: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_829_update_completed_
      -- 
    ca_2120_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_829_inst_ack_1, ack => testConfigure_CP_0_elements(190)); -- 
    -- CP-element group 191:  transition  input  output  bypass 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	188 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	192 
    -- CP-element group 191:  members (6) 
      -- CP-element group 191: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_843_sample_completed_
      -- CP-element group 191: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_843_Update/cr
      -- CP-element group 191: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_843_update_start_
      -- CP-element group 191: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_843_Sample/ra
      -- CP-element group 191: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_843_Sample/$exit
      -- CP-element group 191: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_843_Update/$entry
      -- 
    ra_2129_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_843_inst_ack_0, ack => testConfigure_CP_0_elements(191)); -- 
    cr_2133_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2133_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(191), ack => RPIPE_ConvTranspose_input_pipe_843_inst_req_1); -- 
    -- CP-element group 192:  fork  transition  input  output  bypass 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	191 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	193 
    -- CP-element group 192: 	195 
    -- CP-element group 192:  members (9) 
      -- CP-element group 192: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_843_Update/$exit
      -- CP-element group 192: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_861_Sample/rr
      -- CP-element group 192: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_861_Sample/$entry
      -- CP-element group 192: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_843_update_completed_
      -- CP-element group 192: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_843_Update/ca
      -- CP-element group 192: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_847_sample_start_
      -- CP-element group 192: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_847_Sample/$entry
      -- CP-element group 192: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_847_Sample/rr
      -- CP-element group 192: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_861_sample_start_
      -- 
    ca_2134_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_843_inst_ack_1, ack => testConfigure_CP_0_elements(192)); -- 
    rr_2142_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2142_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(192), ack => type_cast_847_inst_req_0); -- 
    rr_2156_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2156_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(192), ack => RPIPE_ConvTranspose_input_pipe_861_inst_req_0); -- 
    -- CP-element group 193:  transition  input  bypass 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	192 
    -- CP-element group 193: successors 
    -- CP-element group 193:  members (3) 
      -- CP-element group 193: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_847_sample_completed_
      -- CP-element group 193: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_847_Sample/$exit
      -- CP-element group 193: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_847_Sample/ra
      -- 
    ra_2143_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_847_inst_ack_0, ack => testConfigure_CP_0_elements(193)); -- 
    -- CP-element group 194:  transition  input  bypass 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	277 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	207 
    -- CP-element group 194:  members (3) 
      -- CP-element group 194: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_847_update_completed_
      -- CP-element group 194: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_847_Update/ca
      -- CP-element group 194: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_847_Update/$exit
      -- 
    ca_2148_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_847_inst_ack_1, ack => testConfigure_CP_0_elements(194)); -- 
    -- CP-element group 195:  transition  input  output  bypass 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	192 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	196 
    -- CP-element group 195:  members (6) 
      -- CP-element group 195: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_861_Update/$entry
      -- CP-element group 195: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_861_Update/cr
      -- CP-element group 195: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_861_Sample/$exit
      -- CP-element group 195: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_861_Sample/ra
      -- CP-element group 195: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_861_update_start_
      -- CP-element group 195: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_861_sample_completed_
      -- 
    ra_2157_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_861_inst_ack_0, ack => testConfigure_CP_0_elements(195)); -- 
    cr_2161_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2161_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(195), ack => RPIPE_ConvTranspose_input_pipe_861_inst_req_1); -- 
    -- CP-element group 196:  fork  transition  input  output  bypass 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	195 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	197 
    -- CP-element group 196: 	199 
    -- CP-element group 196:  members (9) 
      -- CP-element group 196: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_861_Update/$exit
      -- CP-element group 196: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_861_Update/ca
      -- CP-element group 196: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_865_sample_start_
      -- CP-element group 196: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_861_update_completed_
      -- CP-element group 196: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_879_Sample/rr
      -- CP-element group 196: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_879_Sample/$entry
      -- CP-element group 196: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_879_sample_start_
      -- CP-element group 196: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_865_Sample/rr
      -- CP-element group 196: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_865_Sample/$entry
      -- 
    ca_2162_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_861_inst_ack_1, ack => testConfigure_CP_0_elements(196)); -- 
    rr_2170_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2170_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(196), ack => type_cast_865_inst_req_0); -- 
    rr_2184_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2184_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(196), ack => RPIPE_ConvTranspose_input_pipe_879_inst_req_0); -- 
    -- CP-element group 197:  transition  input  bypass 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	196 
    -- CP-element group 197: successors 
    -- CP-element group 197:  members (3) 
      -- CP-element group 197: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_865_sample_completed_
      -- CP-element group 197: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_865_Sample/ra
      -- CP-element group 197: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_865_Sample/$exit
      -- 
    ra_2171_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_865_inst_ack_0, ack => testConfigure_CP_0_elements(197)); -- 
    -- CP-element group 198:  transition  input  bypass 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	277 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	207 
    -- CP-element group 198:  members (3) 
      -- CP-element group 198: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_865_Update/ca
      -- CP-element group 198: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_865_Update/$exit
      -- CP-element group 198: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_865_update_completed_
      -- 
    ca_2176_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_865_inst_ack_1, ack => testConfigure_CP_0_elements(198)); -- 
    -- CP-element group 199:  transition  input  output  bypass 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	196 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	200 
    -- CP-element group 199:  members (6) 
      -- CP-element group 199: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_879_Update/cr
      -- CP-element group 199: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_879_Update/$entry
      -- CP-element group 199: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_879_Sample/ra
      -- CP-element group 199: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_879_Sample/$exit
      -- CP-element group 199: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_879_update_start_
      -- CP-element group 199: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_879_sample_completed_
      -- 
    ra_2185_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_879_inst_ack_0, ack => testConfigure_CP_0_elements(199)); -- 
    cr_2189_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2189_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(199), ack => RPIPE_ConvTranspose_input_pipe_879_inst_req_1); -- 
    -- CP-element group 200:  fork  transition  input  output  bypass 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	199 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	201 
    -- CP-element group 200: 	203 
    -- CP-element group 200:  members (9) 
      -- CP-element group 200: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_897_sample_start_
      -- CP-element group 200: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_883_Sample/$entry
      -- CP-element group 200: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_883_Sample/rr
      -- CP-element group 200: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_897_Sample/$entry
      -- CP-element group 200: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_897_Sample/rr
      -- CP-element group 200: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_883_sample_start_
      -- CP-element group 200: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_879_Update/ca
      -- CP-element group 200: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_879_Update/$exit
      -- CP-element group 200: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_879_update_completed_
      -- 
    ca_2190_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 200_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_879_inst_ack_1, ack => testConfigure_CP_0_elements(200)); -- 
    rr_2198_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2198_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(200), ack => type_cast_883_inst_req_0); -- 
    rr_2212_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2212_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(200), ack => RPIPE_ConvTranspose_input_pipe_897_inst_req_0); -- 
    -- CP-element group 201:  transition  input  bypass 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	200 
    -- CP-element group 201: successors 
    -- CP-element group 201:  members (3) 
      -- CP-element group 201: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_883_Sample/ra
      -- CP-element group 201: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_883_Sample/$exit
      -- CP-element group 201: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_883_sample_completed_
      -- 
    ra_2199_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_883_inst_ack_0, ack => testConfigure_CP_0_elements(201)); -- 
    -- CP-element group 202:  transition  input  bypass 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	277 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	207 
    -- CP-element group 202:  members (3) 
      -- CP-element group 202: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_883_Update/ca
      -- CP-element group 202: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_883_Update/$exit
      -- CP-element group 202: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_883_update_completed_
      -- 
    ca_2204_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_883_inst_ack_1, ack => testConfigure_CP_0_elements(202)); -- 
    -- CP-element group 203:  transition  input  output  bypass 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	200 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	204 
    -- CP-element group 203:  members (6) 
      -- CP-element group 203: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_897_sample_completed_
      -- CP-element group 203: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_897_update_start_
      -- CP-element group 203: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_897_Sample/$exit
      -- CP-element group 203: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_897_Sample/ra
      -- CP-element group 203: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_897_Update/$entry
      -- CP-element group 203: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_897_Update/cr
      -- 
    ra_2213_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 203_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_897_inst_ack_0, ack => testConfigure_CP_0_elements(203)); -- 
    cr_2217_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2217_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(203), ack => RPIPE_ConvTranspose_input_pipe_897_inst_req_1); -- 
    -- CP-element group 204:  transition  input  output  bypass 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	203 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	205 
    -- CP-element group 204:  members (6) 
      -- CP-element group 204: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_897_update_completed_
      -- CP-element group 204: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_897_Update/$exit
      -- CP-element group 204: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_897_Update/ca
      -- CP-element group 204: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_901_sample_start_
      -- CP-element group 204: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_901_Sample/rr
      -- CP-element group 204: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_901_Sample/$entry
      -- 
    ca_2218_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 204_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_897_inst_ack_1, ack => testConfigure_CP_0_elements(204)); -- 
    rr_2226_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2226_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(204), ack => type_cast_901_inst_req_0); -- 
    -- CP-element group 205:  transition  input  bypass 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	204 
    -- CP-element group 205: successors 
    -- CP-element group 205:  members (3) 
      -- CP-element group 205: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_901_sample_completed_
      -- CP-element group 205: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_901_Sample/ra
      -- CP-element group 205: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_901_Sample/$exit
      -- 
    ra_2227_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_901_inst_ack_0, ack => testConfigure_CP_0_elements(205)); -- 
    -- CP-element group 206:  transition  input  bypass 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	277 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	207 
    -- CP-element group 206:  members (3) 
      -- CP-element group 206: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_901_Update/$exit
      -- CP-element group 206: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_901_Update/ca
      -- CP-element group 206: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_901_update_completed_
      -- 
    ca_2232_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 206_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_901_inst_ack_1, ack => testConfigure_CP_0_elements(206)); -- 
    -- CP-element group 207:  join  transition  output  bypass 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	174 
    -- CP-element group 207: 	178 
    -- CP-element group 207: 	182 
    -- CP-element group 207: 	186 
    -- CP-element group 207: 	190 
    -- CP-element group 207: 	194 
    -- CP-element group 207: 	198 
    -- CP-element group 207: 	202 
    -- CP-element group 207: 	206 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	208 
    -- CP-element group 207:  members (9) 
      -- CP-element group 207: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/ptr_deref_909_sample_start_
      -- CP-element group 207: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/ptr_deref_909_Sample/word_access_start/word_0/rr
      -- CP-element group 207: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/ptr_deref_909_Sample/word_access_start/word_0/$entry
      -- CP-element group 207: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/ptr_deref_909_Sample/word_access_start/$entry
      -- CP-element group 207: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/ptr_deref_909_Sample/ptr_deref_909_Split/split_ack
      -- CP-element group 207: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/ptr_deref_909_Sample/ptr_deref_909_Split/split_req
      -- CP-element group 207: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/ptr_deref_909_Sample/ptr_deref_909_Split/$exit
      -- CP-element group 207: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/ptr_deref_909_Sample/ptr_deref_909_Split/$entry
      -- CP-element group 207: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/ptr_deref_909_Sample/$entry
      -- 
    rr_2270_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2270_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(207), ack => ptr_deref_909_store_0_req_0); -- 
    testConfigure_cp_element_group_207: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_207"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(174) & testConfigure_CP_0_elements(178) & testConfigure_CP_0_elements(182) & testConfigure_CP_0_elements(186) & testConfigure_CP_0_elements(190) & testConfigure_CP_0_elements(194) & testConfigure_CP_0_elements(198) & testConfigure_CP_0_elements(202) & testConfigure_CP_0_elements(206);
      gj_testConfigure_cp_element_group_207 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(207), clk => clk, reset => reset); --
    end block;
    -- CP-element group 208:  transition  input  bypass 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	207 
    -- CP-element group 208: successors 
    -- CP-element group 208:  members (5) 
      -- CP-element group 208: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/ptr_deref_909_sample_completed_
      -- CP-element group 208: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/ptr_deref_909_Sample/word_access_start/word_0/ra
      -- CP-element group 208: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/ptr_deref_909_Sample/word_access_start/word_0/$exit
      -- CP-element group 208: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/ptr_deref_909_Sample/word_access_start/$exit
      -- CP-element group 208: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/ptr_deref_909_Sample/$exit
      -- 
    ra_2271_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 208_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_909_store_0_ack_0, ack => testConfigure_CP_0_elements(208)); -- 
    -- CP-element group 209:  transition  input  bypass 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	277 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	210 
    -- CP-element group 209:  members (5) 
      -- CP-element group 209: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/ptr_deref_909_update_completed_
      -- CP-element group 209: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/ptr_deref_909_Update/word_access_complete/word_0/ca
      -- CP-element group 209: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/ptr_deref_909_Update/word_access_complete/word_0/$exit
      -- CP-element group 209: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/ptr_deref_909_Update/word_access_complete/$exit
      -- CP-element group 209: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/ptr_deref_909_Update/$exit
      -- 
    ca_2282_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_909_store_0_ack_1, ack => testConfigure_CP_0_elements(209)); -- 
    -- CP-element group 210:  branch  join  transition  place  output  bypass 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	171 
    -- CP-element group 210: 	209 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	211 
    -- CP-element group 210: 	212 
    -- CP-element group 210:  members (10) 
      -- CP-element group 210: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922__exit__
      -- CP-element group 210: 	 branch_block_stmt_34/if_stmt_923__entry__
      -- CP-element group 210: 	 branch_block_stmt_34/if_stmt_923_else_link/$entry
      -- CP-element group 210: 	 branch_block_stmt_34/if_stmt_923_if_link/$entry
      -- CP-element group 210: 	 branch_block_stmt_34/if_stmt_923_eval_test/branch_req
      -- CP-element group 210: 	 branch_block_stmt_34/if_stmt_923_eval_test/$exit
      -- CP-element group 210: 	 branch_block_stmt_34/if_stmt_923_eval_test/$entry
      -- CP-element group 210: 	 branch_block_stmt_34/if_stmt_923_dead_link/$entry
      -- CP-element group 210: 	 branch_block_stmt_34/R_exitcond_924_place
      -- CP-element group 210: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/$exit
      -- 
    branch_req_2290_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2290_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(210), ack => if_stmt_923_branch_req_0); -- 
    testConfigure_cp_element_group_210: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_210"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(171) & testConfigure_CP_0_elements(209);
      gj_testConfigure_cp_element_group_210 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(210), clk => clk, reset => reset); --
    end block;
    -- CP-element group 211:  merge  transition  place  input  bypass 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	210 
    -- CP-element group 211: successors 
    -- CP-element group 211: 	278 
    -- CP-element group 211:  members (13) 
      -- CP-element group 211: 	 branch_block_stmt_34/merge_stmt_929__exit__
      -- CP-element group 211: 	 branch_block_stmt_34/forx_xend204x_xloopexit_forx_xend204
      -- CP-element group 211: 	 branch_block_stmt_34/forx_xbody150_forx_xend204x_xloopexit
      -- CP-element group 211: 	 branch_block_stmt_34/if_stmt_923_if_link/if_choice_transition
      -- CP-element group 211: 	 branch_block_stmt_34/if_stmt_923_if_link/$exit
      -- CP-element group 211: 	 branch_block_stmt_34/forx_xbody150_forx_xend204x_xloopexit_PhiReq/$entry
      -- CP-element group 211: 	 branch_block_stmt_34/forx_xbody150_forx_xend204x_xloopexit_PhiReq/$exit
      -- CP-element group 211: 	 branch_block_stmt_34/merge_stmt_929_PhiReqMerge
      -- CP-element group 211: 	 branch_block_stmt_34/merge_stmt_929_PhiAck/$entry
      -- CP-element group 211: 	 branch_block_stmt_34/merge_stmt_929_PhiAck/$exit
      -- CP-element group 211: 	 branch_block_stmt_34/merge_stmt_929_PhiAck/dummy
      -- CP-element group 211: 	 branch_block_stmt_34/forx_xend204x_xloopexit_forx_xend204_PhiReq/$entry
      -- CP-element group 211: 	 branch_block_stmt_34/forx_xend204x_xloopexit_forx_xend204_PhiReq/$exit
      -- 
    if_choice_transition_2295_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 211_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_923_branch_ack_1, ack => testConfigure_CP_0_elements(211)); -- 
    -- CP-element group 212:  fork  transition  place  input  output  bypass 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	210 
    -- CP-element group 212: successors 
    -- CP-element group 212: 	273 
    -- CP-element group 212: 	274 
    -- CP-element group 212:  members (12) 
      -- CP-element group 212: 	 branch_block_stmt_34/forx_xbody150_forx_xbody150
      -- CP-element group 212: 	 branch_block_stmt_34/if_stmt_923_else_link/else_choice_transition
      -- CP-element group 212: 	 branch_block_stmt_34/if_stmt_923_else_link/$exit
      -- CP-element group 212: 	 branch_block_stmt_34/forx_xbody150_forx_xbody150_PhiReq/$entry
      -- CP-element group 212: 	 branch_block_stmt_34/forx_xbody150_forx_xbody150_PhiReq/phi_stmt_760/$entry
      -- CP-element group 212: 	 branch_block_stmt_34/forx_xbody150_forx_xbody150_PhiReq/phi_stmt_760/phi_stmt_760_sources/$entry
      -- CP-element group 212: 	 branch_block_stmt_34/forx_xbody150_forx_xbody150_PhiReq/phi_stmt_760/phi_stmt_760_sources/type_cast_766/$entry
      -- CP-element group 212: 	 branch_block_stmt_34/forx_xbody150_forx_xbody150_PhiReq/phi_stmt_760/phi_stmt_760_sources/type_cast_766/SplitProtocol/$entry
      -- CP-element group 212: 	 branch_block_stmt_34/forx_xbody150_forx_xbody150_PhiReq/phi_stmt_760/phi_stmt_760_sources/type_cast_766/SplitProtocol/Sample/$entry
      -- CP-element group 212: 	 branch_block_stmt_34/forx_xbody150_forx_xbody150_PhiReq/phi_stmt_760/phi_stmt_760_sources/type_cast_766/SplitProtocol/Sample/rr
      -- CP-element group 212: 	 branch_block_stmt_34/forx_xbody150_forx_xbody150_PhiReq/phi_stmt_760/phi_stmt_760_sources/type_cast_766/SplitProtocol/Update/$entry
      -- CP-element group 212: 	 branch_block_stmt_34/forx_xbody150_forx_xbody150_PhiReq/phi_stmt_760/phi_stmt_760_sources/type_cast_766/SplitProtocol/Update/cr
      -- 
    else_choice_transition_2299_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 212_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_923_branch_ack_0, ack => testConfigure_CP_0_elements(212)); -- 
    rr_2962_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2962_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(212), ack => type_cast_766_inst_req_0); -- 
    cr_2967_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2967_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(212), ack => type_cast_766_inst_req_1); -- 
    -- CP-element group 213:  transition  input  bypass 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	279 
    -- CP-element group 213: successors 
    -- CP-element group 213:  members (5) 
      -- CP-element group 213: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_942_Sample/$exit
      -- CP-element group 213: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_942_Sample/word_access_start/$exit
      -- CP-element group 213: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_942_Sample/word_access_start/word_0/$exit
      -- CP-element group 213: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_942_Sample/word_access_start/word_0/ra
      -- CP-element group 213: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_942_sample_completed_
      -- 
    ra_2338_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_942_load_0_ack_0, ack => testConfigure_CP_0_elements(213)); -- 
    -- CP-element group 214:  transition  input  bypass 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	279 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	219 
    -- CP-element group 214:  members (9) 
      -- CP-element group 214: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_942_Update/$exit
      -- CP-element group 214: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_942_Update/word_access_complete/$exit
      -- CP-element group 214: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_942_Update/word_access_complete/word_0/$exit
      -- CP-element group 214: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_942_Update/word_access_complete/word_0/ca
      -- CP-element group 214: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_942_Update/ptr_deref_942_Merge/$entry
      -- CP-element group 214: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_942_Update/ptr_deref_942_Merge/$exit
      -- CP-element group 214: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_942_Update/ptr_deref_942_Merge/merge_req
      -- CP-element group 214: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_942_Update/ptr_deref_942_Merge/merge_ack
      -- CP-element group 214: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_942_update_completed_
      -- 
    ca_2349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 214_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_942_load_0_ack_1, ack => testConfigure_CP_0_elements(214)); -- 
    -- CP-element group 215:  transition  input  bypass 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	279 
    -- CP-element group 215: successors 
    -- CP-element group 215:  members (5) 
      -- CP-element group 215: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_954_Sample/word_access_start/word_0/ra
      -- CP-element group 215: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_954_Sample/word_access_start/word_0/$exit
      -- CP-element group 215: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_954_Sample/word_access_start/$exit
      -- CP-element group 215: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_954_sample_completed_
      -- CP-element group 215: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_954_Sample/$exit
      -- 
    ra_2388_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 215_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_954_load_0_ack_0, ack => testConfigure_CP_0_elements(215)); -- 
    -- CP-element group 216:  transition  input  bypass 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	279 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	219 
    -- CP-element group 216:  members (9) 
      -- CP-element group 216: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_954_Update/$exit
      -- CP-element group 216: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_954_update_completed_
      -- CP-element group 216: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_954_Update/ptr_deref_954_Merge/merge_ack
      -- CP-element group 216: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_954_Update/ptr_deref_954_Merge/merge_req
      -- CP-element group 216: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_954_Update/ptr_deref_954_Merge/$exit
      -- CP-element group 216: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_954_Update/ptr_deref_954_Merge/$entry
      -- CP-element group 216: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_954_Update/word_access_complete/word_0/ca
      -- CP-element group 216: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_954_Update/word_access_complete/word_0/$exit
      -- CP-element group 216: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_954_Update/word_access_complete/$exit
      -- 
    ca_2399_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_954_load_0_ack_1, ack => testConfigure_CP_0_elements(216)); -- 
    -- CP-element group 217:  transition  input  bypass 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	279 
    -- CP-element group 217: successors 
    -- CP-element group 217:  members (5) 
      -- CP-element group 217: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_966_Sample/$exit
      -- CP-element group 217: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_966_Sample/word_access_start/$exit
      -- CP-element group 217: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_966_Sample/word_access_start/word_0/$exit
      -- CP-element group 217: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_966_sample_completed_
      -- CP-element group 217: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_966_Sample/word_access_start/word_0/ra
      -- 
    ra_2438_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 217_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_966_load_0_ack_0, ack => testConfigure_CP_0_elements(217)); -- 
    -- CP-element group 218:  transition  input  bypass 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	279 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	219 
    -- CP-element group 218:  members (9) 
      -- CP-element group 218: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_966_Update/ptr_deref_966_Merge/merge_ack
      -- CP-element group 218: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_966_Update/ptr_deref_966_Merge/merge_req
      -- CP-element group 218: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_966_update_completed_
      -- CP-element group 218: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_966_Update/ptr_deref_966_Merge/$exit
      -- CP-element group 218: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_966_Update/ptr_deref_966_Merge/$entry
      -- CP-element group 218: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_966_Update/word_access_complete/word_0/ca
      -- CP-element group 218: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_966_Update/word_access_complete/word_0/$exit
      -- CP-element group 218: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_966_Update/word_access_complete/$exit
      -- CP-element group 218: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_966_Update/$exit
      -- 
    ca_2449_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 218_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_966_load_0_ack_1, ack => testConfigure_CP_0_elements(218)); -- 
    -- CP-element group 219:  branch  join  transition  place  output  bypass 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	214 
    -- CP-element group 219: 	216 
    -- CP-element group 219: 	218 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	220 
    -- CP-element group 219: 	221 
    -- CP-element group 219:  members (10) 
      -- CP-element group 219: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983__exit__
      -- CP-element group 219: 	 branch_block_stmt_34/if_stmt_984__entry__
      -- CP-element group 219: 	 branch_block_stmt_34/if_stmt_984_eval_test/$entry
      -- CP-element group 219: 	 branch_block_stmt_34/if_stmt_984_dead_link/$entry
      -- CP-element group 219: 	 branch_block_stmt_34/if_stmt_984_eval_test/$exit
      -- CP-element group 219: 	 branch_block_stmt_34/if_stmt_984_if_link/$entry
      -- CP-element group 219: 	 branch_block_stmt_34/if_stmt_984_eval_test/branch_req
      -- CP-element group 219: 	 branch_block_stmt_34/R_cmp215226_985_place
      -- CP-element group 219: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/$exit
      -- CP-element group 219: 	 branch_block_stmt_34/if_stmt_984_else_link/$entry
      -- 
    branch_req_2462_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2462_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(219), ack => if_stmt_984_branch_req_0); -- 
    testConfigure_cp_element_group_219: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_219"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(214) & testConfigure_CP_0_elements(216) & testConfigure_CP_0_elements(218);
      gj_testConfigure_cp_element_group_219 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(219), clk => clk, reset => reset); --
    end block;
    -- CP-element group 220:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	219 
    -- CP-element group 220: successors 
    -- CP-element group 220: 	222 
    -- CP-element group 220: 	223 
    -- CP-element group 220:  members (18) 
      -- CP-element group 220: 	 branch_block_stmt_34/assign_stmt_996_to_assign_stmt_1025/$entry
      -- CP-element group 220: 	 branch_block_stmt_34/assign_stmt_996_to_assign_stmt_1025/type_cast_1011_Sample/rr
      -- CP-element group 220: 	 branch_block_stmt_34/merge_stmt_990__exit__
      -- CP-element group 220: 	 branch_block_stmt_34/assign_stmt_996_to_assign_stmt_1025__entry__
      -- CP-element group 220: 	 branch_block_stmt_34/assign_stmt_996_to_assign_stmt_1025/type_cast_1011_sample_start_
      -- CP-element group 220: 	 branch_block_stmt_34/if_stmt_984_if_link/if_choice_transition
      -- CP-element group 220: 	 branch_block_stmt_34/if_stmt_984_if_link/$exit
      -- CP-element group 220: 	 branch_block_stmt_34/assign_stmt_996_to_assign_stmt_1025/type_cast_1011_update_start_
      -- CP-element group 220: 	 branch_block_stmt_34/assign_stmt_996_to_assign_stmt_1025/type_cast_1011_Update/$entry
      -- CP-element group 220: 	 branch_block_stmt_34/assign_stmt_996_to_assign_stmt_1025/type_cast_1011_Sample/$entry
      -- CP-element group 220: 	 branch_block_stmt_34/forx_xend204_bbx_xnph
      -- CP-element group 220: 	 branch_block_stmt_34/assign_stmt_996_to_assign_stmt_1025/type_cast_1011_Update/cr
      -- CP-element group 220: 	 branch_block_stmt_34/forx_xend204_bbx_xnph_PhiReq/$entry
      -- CP-element group 220: 	 branch_block_stmt_34/forx_xend204_bbx_xnph_PhiReq/$exit
      -- CP-element group 220: 	 branch_block_stmt_34/merge_stmt_990_PhiReqMerge
      -- CP-element group 220: 	 branch_block_stmt_34/merge_stmt_990_PhiAck/$entry
      -- CP-element group 220: 	 branch_block_stmt_34/merge_stmt_990_PhiAck/$exit
      -- CP-element group 220: 	 branch_block_stmt_34/merge_stmt_990_PhiAck/dummy
      -- 
    if_choice_transition_2467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_984_branch_ack_1, ack => testConfigure_CP_0_elements(220)); -- 
    rr_2484_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2484_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(220), ack => type_cast_1011_inst_req_0); -- 
    cr_2489_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2489_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(220), ack => type_cast_1011_inst_req_1); -- 
    -- CP-element group 221:  transition  place  input  bypass 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	219 
    -- CP-element group 221: successors 
    -- CP-element group 221: 	286 
    -- CP-element group 221:  members (5) 
      -- CP-element group 221: 	 branch_block_stmt_34/forx_xend204_forx_xend224
      -- CP-element group 221: 	 branch_block_stmt_34/if_stmt_984_else_link/else_choice_transition
      -- CP-element group 221: 	 branch_block_stmt_34/if_stmt_984_else_link/$exit
      -- CP-element group 221: 	 branch_block_stmt_34/forx_xend204_forx_xend224_PhiReq/$entry
      -- CP-element group 221: 	 branch_block_stmt_34/forx_xend204_forx_xend224_PhiReq/$exit
      -- 
    else_choice_transition_2471_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_984_branch_ack_0, ack => testConfigure_CP_0_elements(221)); -- 
    -- CP-element group 222:  transition  input  bypass 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	220 
    -- CP-element group 222: successors 
    -- CP-element group 222:  members (3) 
      -- CP-element group 222: 	 branch_block_stmt_34/assign_stmt_996_to_assign_stmt_1025/type_cast_1011_Sample/$exit
      -- CP-element group 222: 	 branch_block_stmt_34/assign_stmt_996_to_assign_stmt_1025/type_cast_1011_Sample/ra
      -- CP-element group 222: 	 branch_block_stmt_34/assign_stmt_996_to_assign_stmt_1025/type_cast_1011_sample_completed_
      -- 
    ra_2485_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 222_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1011_inst_ack_0, ack => testConfigure_CP_0_elements(222)); -- 
    -- CP-element group 223:  transition  place  input  bypass 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	220 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	280 
    -- CP-element group 223:  members (9) 
      -- CP-element group 223: 	 branch_block_stmt_34/assign_stmt_996_to_assign_stmt_1025__exit__
      -- CP-element group 223: 	 branch_block_stmt_34/bbx_xnph_forx_xbody217
      -- CP-element group 223: 	 branch_block_stmt_34/assign_stmt_996_to_assign_stmt_1025/$exit
      -- CP-element group 223: 	 branch_block_stmt_34/assign_stmt_996_to_assign_stmt_1025/type_cast_1011_update_completed_
      -- CP-element group 223: 	 branch_block_stmt_34/assign_stmt_996_to_assign_stmt_1025/type_cast_1011_Update/ca
      -- CP-element group 223: 	 branch_block_stmt_34/assign_stmt_996_to_assign_stmt_1025/type_cast_1011_Update/$exit
      -- CP-element group 223: 	 branch_block_stmt_34/bbx_xnph_forx_xbody217_PhiReq/$entry
      -- CP-element group 223: 	 branch_block_stmt_34/bbx_xnph_forx_xbody217_PhiReq/phi_stmt_1028/$entry
      -- CP-element group 223: 	 branch_block_stmt_34/bbx_xnph_forx_xbody217_PhiReq/phi_stmt_1028/phi_stmt_1028_sources/$entry
      -- 
    ca_2490_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 223_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1011_inst_ack_1, ack => testConfigure_CP_0_elements(223)); -- 
    -- CP-element group 224:  transition  input  bypass 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	285 
    -- CP-element group 224: successors 
    -- CP-element group 224: 	230 
    -- CP-element group 224:  members (3) 
      -- CP-element group 224: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/array_obj_ref_1040_final_index_sum_regn_Sample/ack
      -- CP-element group 224: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/array_obj_ref_1040_final_index_sum_regn_Sample/$exit
      -- CP-element group 224: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/array_obj_ref_1040_final_index_sum_regn_sample_complete
      -- 
    ack_2519_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1040_index_offset_ack_0, ack => testConfigure_CP_0_elements(224)); -- 
    -- CP-element group 225:  transition  input  output  bypass 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	285 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	226 
    -- CP-element group 225:  members (11) 
      -- CP-element group 225: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/array_obj_ref_1040_final_index_sum_regn_Update/$exit
      -- CP-element group 225: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/array_obj_ref_1040_offset_calculated
      -- CP-element group 225: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/addr_of_1041_request/req
      -- CP-element group 225: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/array_obj_ref_1040_final_index_sum_regn_Update/ack
      -- CP-element group 225: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/array_obj_ref_1040_root_address_calculated
      -- CP-element group 225: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/addr_of_1041_request/$entry
      -- CP-element group 225: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/addr_of_1041_sample_start_
      -- CP-element group 225: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/array_obj_ref_1040_base_plus_offset/sum_rename_ack
      -- CP-element group 225: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/array_obj_ref_1040_base_plus_offset/sum_rename_req
      -- CP-element group 225: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/array_obj_ref_1040_base_plus_offset/$exit
      -- CP-element group 225: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/array_obj_ref_1040_base_plus_offset/$entry
      -- 
    ack_2524_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 225_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1040_index_offset_ack_1, ack => testConfigure_CP_0_elements(225)); -- 
    req_2533_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2533_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(225), ack => addr_of_1041_final_reg_req_0); -- 
    -- CP-element group 226:  transition  input  bypass 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	225 
    -- CP-element group 226: successors 
    -- CP-element group 226:  members (3) 
      -- CP-element group 226: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/addr_of_1041_request/ack
      -- CP-element group 226: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/addr_of_1041_request/$exit
      -- CP-element group 226: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/addr_of_1041_sample_completed_
      -- 
    ack_2534_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 226_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1041_final_reg_ack_0, ack => testConfigure_CP_0_elements(226)); -- 
    -- CP-element group 227:  join  fork  transition  input  output  bypass 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	285 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	228 
    -- CP-element group 227:  members (28) 
      -- CP-element group 227: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/ptr_deref_1044_word_addrgen/root_register_req
      -- CP-element group 227: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/ptr_deref_1044_base_plus_offset/sum_rename_req
      -- CP-element group 227: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/ptr_deref_1044_Sample/ptr_deref_1044_Split/split_ack
      -- CP-element group 227: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/ptr_deref_1044_root_address_calculated
      -- CP-element group 227: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/ptr_deref_1044_word_address_calculated
      -- CP-element group 227: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/ptr_deref_1044_base_plus_offset/$exit
      -- CP-element group 227: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/addr_of_1041_complete/$exit
      -- CP-element group 227: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/ptr_deref_1044_base_plus_offset/$entry
      -- CP-element group 227: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/addr_of_1041_update_completed_
      -- CP-element group 227: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/ptr_deref_1044_Sample/ptr_deref_1044_Split/split_req
      -- CP-element group 227: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/ptr_deref_1044_base_address_calculated
      -- CP-element group 227: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/ptr_deref_1044_Sample/ptr_deref_1044_Split/$exit
      -- CP-element group 227: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/ptr_deref_1044_word_addrgen/$entry
      -- CP-element group 227: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/ptr_deref_1044_word_addrgen/$exit
      -- CP-element group 227: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/addr_of_1041_complete/ack
      -- CP-element group 227: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/ptr_deref_1044_Sample/ptr_deref_1044_Split/$entry
      -- CP-element group 227: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/ptr_deref_1044_base_addr_resize/base_resize_ack
      -- CP-element group 227: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/ptr_deref_1044_Sample/$entry
      -- CP-element group 227: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/ptr_deref_1044_base_addr_resize/base_resize_req
      -- CP-element group 227: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/ptr_deref_1044_sample_start_
      -- CP-element group 227: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/ptr_deref_1044_base_addr_resize/$exit
      -- CP-element group 227: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/ptr_deref_1044_base_plus_offset/sum_rename_ack
      -- CP-element group 227: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/ptr_deref_1044_base_addr_resize/$entry
      -- CP-element group 227: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/ptr_deref_1044_word_addrgen/root_register_ack
      -- CP-element group 227: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/ptr_deref_1044_base_address_resized
      -- CP-element group 227: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/ptr_deref_1044_Sample/word_access_start/$entry
      -- CP-element group 227: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/ptr_deref_1044_Sample/word_access_start/word_0/$entry
      -- CP-element group 227: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/ptr_deref_1044_Sample/word_access_start/word_0/rr
      -- 
    ack_2539_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 227_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1041_final_reg_ack_1, ack => testConfigure_CP_0_elements(227)); -- 
    rr_2577_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2577_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(227), ack => ptr_deref_1044_store_0_req_0); -- 
    -- CP-element group 228:  transition  input  bypass 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	227 
    -- CP-element group 228: successors 
    -- CP-element group 228:  members (5) 
      -- CP-element group 228: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/ptr_deref_1044_Sample/$exit
      -- CP-element group 228: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/ptr_deref_1044_sample_completed_
      -- CP-element group 228: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/ptr_deref_1044_Sample/word_access_start/$exit
      -- CP-element group 228: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/ptr_deref_1044_Sample/word_access_start/word_0/$exit
      -- CP-element group 228: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/ptr_deref_1044_Sample/word_access_start/word_0/ra
      -- 
    ra_2578_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 228_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1044_store_0_ack_0, ack => testConfigure_CP_0_elements(228)); -- 
    -- CP-element group 229:  transition  input  bypass 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	285 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	230 
    -- CP-element group 229:  members (5) 
      -- CP-element group 229: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/ptr_deref_1044_update_completed_
      -- CP-element group 229: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/ptr_deref_1044_Update/$exit
      -- CP-element group 229: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/ptr_deref_1044_Update/word_access_complete/$exit
      -- CP-element group 229: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/ptr_deref_1044_Update/word_access_complete/word_0/$exit
      -- CP-element group 229: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/ptr_deref_1044_Update/word_access_complete/word_0/ca
      -- 
    ca_2589_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 229_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1044_store_0_ack_1, ack => testConfigure_CP_0_elements(229)); -- 
    -- CP-element group 230:  branch  join  transition  place  output  bypass 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	224 
    -- CP-element group 230: 	229 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	231 
    -- CP-element group 230: 	232 
    -- CP-element group 230:  members (10) 
      -- CP-element group 230: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058__exit__
      -- CP-element group 230: 	 branch_block_stmt_34/if_stmt_1059__entry__
      -- CP-element group 230: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/$exit
      -- CP-element group 230: 	 branch_block_stmt_34/if_stmt_1059_dead_link/$entry
      -- CP-element group 230: 	 branch_block_stmt_34/if_stmt_1059_eval_test/$entry
      -- CP-element group 230: 	 branch_block_stmt_34/if_stmt_1059_eval_test/$exit
      -- CP-element group 230: 	 branch_block_stmt_34/if_stmt_1059_eval_test/branch_req
      -- CP-element group 230: 	 branch_block_stmt_34/R_exitcond1_1060_place
      -- CP-element group 230: 	 branch_block_stmt_34/if_stmt_1059_if_link/$entry
      -- CP-element group 230: 	 branch_block_stmt_34/if_stmt_1059_else_link/$entry
      -- 
    branch_req_2597_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2597_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(230), ack => if_stmt_1059_branch_req_0); -- 
    testConfigure_cp_element_group_230: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_230"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(224) & testConfigure_CP_0_elements(229);
      gj_testConfigure_cp_element_group_230 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(230), clk => clk, reset => reset); --
    end block;
    -- CP-element group 231:  merge  transition  place  input  bypass 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	230 
    -- CP-element group 231: successors 
    -- CP-element group 231: 	286 
    -- CP-element group 231:  members (13) 
      -- CP-element group 231: 	 branch_block_stmt_34/merge_stmt_1065__exit__
      -- CP-element group 231: 	 branch_block_stmt_34/forx_xend224x_xloopexit_forx_xend224
      -- CP-element group 231: 	 branch_block_stmt_34/if_stmt_1059_if_link/$exit
      -- CP-element group 231: 	 branch_block_stmt_34/if_stmt_1059_if_link/if_choice_transition
      -- CP-element group 231: 	 branch_block_stmt_34/forx_xbody217_forx_xend224x_xloopexit
      -- CP-element group 231: 	 branch_block_stmt_34/forx_xbody217_forx_xend224x_xloopexit_PhiReq/$entry
      -- CP-element group 231: 	 branch_block_stmt_34/forx_xbody217_forx_xend224x_xloopexit_PhiReq/$exit
      -- CP-element group 231: 	 branch_block_stmt_34/merge_stmt_1065_PhiReqMerge
      -- CP-element group 231: 	 branch_block_stmt_34/merge_stmt_1065_PhiAck/$entry
      -- CP-element group 231: 	 branch_block_stmt_34/merge_stmt_1065_PhiAck/$exit
      -- CP-element group 231: 	 branch_block_stmt_34/merge_stmt_1065_PhiAck/dummy
      -- CP-element group 231: 	 branch_block_stmt_34/forx_xend224x_xloopexit_forx_xend224_PhiReq/$entry
      -- CP-element group 231: 	 branch_block_stmt_34/forx_xend224x_xloopexit_forx_xend224_PhiReq/$exit
      -- 
    if_choice_transition_2602_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 231_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1059_branch_ack_1, ack => testConfigure_CP_0_elements(231)); -- 
    -- CP-element group 232:  fork  transition  place  input  output  bypass 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	230 
    -- CP-element group 232: successors 
    -- CP-element group 232: 	281 
    -- CP-element group 232: 	282 
    -- CP-element group 232:  members (12) 
      -- CP-element group 232: 	 branch_block_stmt_34/if_stmt_1059_else_link/$exit
      -- CP-element group 232: 	 branch_block_stmt_34/if_stmt_1059_else_link/else_choice_transition
      -- CP-element group 232: 	 branch_block_stmt_34/forx_xbody217_forx_xbody217
      -- CP-element group 232: 	 branch_block_stmt_34/forx_xbody217_forx_xbody217_PhiReq/$entry
      -- CP-element group 232: 	 branch_block_stmt_34/forx_xbody217_forx_xbody217_PhiReq/phi_stmt_1028/$entry
      -- CP-element group 232: 	 branch_block_stmt_34/forx_xbody217_forx_xbody217_PhiReq/phi_stmt_1028/phi_stmt_1028_sources/$entry
      -- CP-element group 232: 	 branch_block_stmt_34/forx_xbody217_forx_xbody217_PhiReq/phi_stmt_1028/phi_stmt_1028_sources/type_cast_1034/$entry
      -- CP-element group 232: 	 branch_block_stmt_34/forx_xbody217_forx_xbody217_PhiReq/phi_stmt_1028/phi_stmt_1028_sources/type_cast_1034/SplitProtocol/$entry
      -- CP-element group 232: 	 branch_block_stmt_34/forx_xbody217_forx_xbody217_PhiReq/phi_stmt_1028/phi_stmt_1028_sources/type_cast_1034/SplitProtocol/Sample/$entry
      -- CP-element group 232: 	 branch_block_stmt_34/forx_xbody217_forx_xbody217_PhiReq/phi_stmt_1028/phi_stmt_1028_sources/type_cast_1034/SplitProtocol/Sample/rr
      -- CP-element group 232: 	 branch_block_stmt_34/forx_xbody217_forx_xbody217_PhiReq/phi_stmt_1028/phi_stmt_1028_sources/type_cast_1034/SplitProtocol/Update/$entry
      -- CP-element group 232: 	 branch_block_stmt_34/forx_xbody217_forx_xbody217_PhiReq/phi_stmt_1028/phi_stmt_1028_sources/type_cast_1034/SplitProtocol/Update/cr
      -- 
    else_choice_transition_2606_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 232_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1059_branch_ack_0, ack => testConfigure_CP_0_elements(232)); -- 
    rr_3039_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3039_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(232), ack => type_cast_1034_inst_req_0); -- 
    cr_3044_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3044_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(232), ack => type_cast_1034_inst_req_1); -- 
    -- CP-element group 233:  transition  output  delay-element  bypass 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	0 
    -- CP-element group 233: successors 
    -- CP-element group 233: 	237 
    -- CP-element group 233:  members (5) 
      -- CP-element group 233: 	 branch_block_stmt_34/bbx_xnph246_forx_xbody_PhiReq/$exit
      -- CP-element group 233: 	 branch_block_stmt_34/bbx_xnph246_forx_xbody_PhiReq/phi_stmt_37/$exit
      -- CP-element group 233: 	 branch_block_stmt_34/bbx_xnph246_forx_xbody_PhiReq/phi_stmt_37/phi_stmt_37_sources/$exit
      -- CP-element group 233: 	 branch_block_stmt_34/bbx_xnph246_forx_xbody_PhiReq/phi_stmt_37/phi_stmt_37_sources/type_cast_41_konst_delay_trans
      -- CP-element group 233: 	 branch_block_stmt_34/bbx_xnph246_forx_xbody_PhiReq/phi_stmt_37/phi_stmt_37_req
      -- 
    phi_stmt_37_req_2622_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_37_req_2622_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(233), ack => phi_stmt_37_req_0); -- 
    -- Element group testConfigure_CP_0_elements(233) is a control-delay.
    cp_element_233_delay: control_delay_element  generic map(name => " 233_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(0), ack => testConfigure_CP_0_elements(233), clk => clk, reset =>reset);
    -- CP-element group 234:  transition  input  bypass 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	22 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	236 
    -- CP-element group 234:  members (2) 
      -- CP-element group 234: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_37/phi_stmt_37_sources/type_cast_43/SplitProtocol/Sample/$exit
      -- CP-element group 234: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_37/phi_stmt_37_sources/type_cast_43/SplitProtocol/Sample/ra
      -- 
    ra_2642_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 234_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_43_inst_ack_0, ack => testConfigure_CP_0_elements(234)); -- 
    -- CP-element group 235:  transition  input  bypass 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	22 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	236 
    -- CP-element group 235:  members (2) 
      -- CP-element group 235: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_37/phi_stmt_37_sources/type_cast_43/SplitProtocol/Update/$exit
      -- CP-element group 235: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_37/phi_stmt_37_sources/type_cast_43/SplitProtocol/Update/ca
      -- 
    ca_2647_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 235_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_43_inst_ack_1, ack => testConfigure_CP_0_elements(235)); -- 
    -- CP-element group 236:  join  transition  output  bypass 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	234 
    -- CP-element group 236: 	235 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	237 
    -- CP-element group 236:  members (6) 
      -- CP-element group 236: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 236: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_37/$exit
      -- CP-element group 236: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_37/phi_stmt_37_sources/$exit
      -- CP-element group 236: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_37/phi_stmt_37_sources/type_cast_43/$exit
      -- CP-element group 236: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_37/phi_stmt_37_sources/type_cast_43/SplitProtocol/$exit
      -- CP-element group 236: 	 branch_block_stmt_34/forx_xbody_forx_xbody_PhiReq/phi_stmt_37/phi_stmt_37_req
      -- 
    phi_stmt_37_req_2648_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_37_req_2648_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(236), ack => phi_stmt_37_req_1); -- 
    testConfigure_cp_element_group_236: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_236"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(234) & testConfigure_CP_0_elements(235);
      gj_testConfigure_cp_element_group_236 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(236), clk => clk, reset => reset); --
    end block;
    -- CP-element group 237:  merge  transition  place  bypass 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	233 
    -- CP-element group 237: 	236 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	238 
    -- CP-element group 237:  members (2) 
      -- CP-element group 237: 	 branch_block_stmt_34/merge_stmt_36_PhiReqMerge
      -- CP-element group 237: 	 branch_block_stmt_34/merge_stmt_36_PhiAck/$entry
      -- 
    testConfigure_CP_0_elements(237) <= OrReduce(testConfigure_CP_0_elements(233) & testConfigure_CP_0_elements(236));
    -- CP-element group 238:  fork  transition  place  input  output  bypass 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	237 
    -- CP-element group 238: successors 
    -- CP-element group 238: 	11 
    -- CP-element group 238: 	15 
    -- CP-element group 238: 	18 
    -- CP-element group 238: 	1 
    -- CP-element group 238: 	2 
    -- CP-element group 238: 	4 
    -- CP-element group 238: 	5 
    -- CP-element group 238: 	8 
    -- CP-element group 238:  members (43) 
      -- CP-element group 238: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/array_obj_ref_49_final_index_sum_regn_Update/$entry
      -- CP-element group 238: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/array_obj_ref_49_final_index_sum_regn_Update/req
      -- CP-element group 238: 	 branch_block_stmt_34/merge_stmt_36__exit__
      -- CP-element group 238: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97__entry__
      -- CP-element group 238: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/$entry
      -- CP-element group 238: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/addr_of_50_update_start_
      -- CP-element group 238: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/array_obj_ref_49_index_resized_1
      -- CP-element group 238: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/array_obj_ref_49_index_scaled_1
      -- CP-element group 238: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/array_obj_ref_49_index_computed_1
      -- CP-element group 238: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/array_obj_ref_49_index_resize_1/$entry
      -- CP-element group 238: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/array_obj_ref_49_index_resize_1/$exit
      -- CP-element group 238: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/array_obj_ref_49_index_resize_1/index_resize_req
      -- CP-element group 238: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/array_obj_ref_49_index_resize_1/index_resize_ack
      -- CP-element group 238: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/array_obj_ref_49_index_scale_1/$entry
      -- CP-element group 238: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/array_obj_ref_49_index_scale_1/$exit
      -- CP-element group 238: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/array_obj_ref_49_index_scale_1/scale_rename_req
      -- CP-element group 238: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/array_obj_ref_49_index_scale_1/scale_rename_ack
      -- CP-element group 238: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/array_obj_ref_49_final_index_sum_regn_update_start
      -- CP-element group 238: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/array_obj_ref_49_final_index_sum_regn_Sample/$entry
      -- CP-element group 238: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/array_obj_ref_49_final_index_sum_regn_Sample/req
      -- CP-element group 238: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/addr_of_50_complete/$entry
      -- CP-element group 238: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/addr_of_50_complete/req
      -- CP-element group 238: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/RPIPE_ConvTranspose_input_pipe_53_sample_start_
      -- CP-element group 238: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/RPIPE_ConvTranspose_input_pipe_53_Sample/$entry
      -- CP-element group 238: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/RPIPE_ConvTranspose_input_pipe_53_Sample/rr
      -- CP-element group 238: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/type_cast_57_update_start_
      -- CP-element group 238: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/type_cast_57_Update/$entry
      -- CP-element group 238: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/type_cast_57_Update/cr
      -- CP-element group 238: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_60_update_start_
      -- CP-element group 238: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_60_Update/$entry
      -- CP-element group 238: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_60_Update/word_access_complete/$entry
      -- CP-element group 238: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_60_Update/word_access_complete/word_0/$entry
      -- CP-element group 238: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_60_Update/word_access_complete/word_0/cr
      -- CP-element group 238: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/type_cast_74_update_start_
      -- CP-element group 238: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/type_cast_74_Update/$entry
      -- CP-element group 238: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/type_cast_74_Update/cr
      -- CP-element group 238: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_82_update_start_
      -- CP-element group 238: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_82_Update/$entry
      -- CP-element group 238: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_82_Update/word_access_complete/$entry
      -- CP-element group 238: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_82_Update/word_access_complete/word_0/$entry
      -- CP-element group 238: 	 branch_block_stmt_34/assign_stmt_51_to_assign_stmt_97/ptr_deref_82_Update/word_access_complete/word_0/cr
      -- CP-element group 238: 	 branch_block_stmt_34/merge_stmt_36_PhiAck/$exit
      -- CP-element group 238: 	 branch_block_stmt_34/merge_stmt_36_PhiAck/phi_stmt_37_ack
      -- 
    phi_stmt_37_ack_2653_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 238_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_37_ack_0, ack => testConfigure_CP_0_elements(238)); -- 
    req_124_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_124_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(238), ack => array_obj_ref_49_index_offset_req_1); -- 
    req_119_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_119_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(238), ack => array_obj_ref_49_index_offset_req_0); -- 
    req_139_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_139_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(238), ack => addr_of_50_final_reg_req_1); -- 
    rr_148_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_148_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(238), ack => RPIPE_ConvTranspose_input_pipe_53_inst_req_0); -- 
    cr_167_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_167_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(238), ack => type_cast_57_inst_req_1); -- 
    cr_217_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_217_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(238), ack => ptr_deref_60_store_0_req_1); -- 
    cr_245_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_245_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(238), ack => type_cast_74_inst_req_1); -- 
    cr_295_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_295_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(238), ack => ptr_deref_82_store_0_req_1); -- 
    -- CP-element group 239:  transition  input  bypass 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	44 
    -- CP-element group 239: successors 
    -- CP-element group 239: 	241 
    -- CP-element group 239:  members (2) 
      -- CP-element group 239: 	 branch_block_stmt_34/forx_xbody16_forx_xbody16_PhiReq/phi_stmt_107/phi_stmt_107_sources/type_cast_110/SplitProtocol/Sample/$exit
      -- CP-element group 239: 	 branch_block_stmt_34/forx_xbody16_forx_xbody16_PhiReq/phi_stmt_107/phi_stmt_107_sources/type_cast_110/SplitProtocol/Sample/ra
      -- 
    ra_2685_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 239_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_110_inst_ack_0, ack => testConfigure_CP_0_elements(239)); -- 
    -- CP-element group 240:  transition  input  bypass 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	44 
    -- CP-element group 240: successors 
    -- CP-element group 240: 	241 
    -- CP-element group 240:  members (2) 
      -- CP-element group 240: 	 branch_block_stmt_34/forx_xbody16_forx_xbody16_PhiReq/phi_stmt_107/phi_stmt_107_sources/type_cast_110/SplitProtocol/Update/$exit
      -- CP-element group 240: 	 branch_block_stmt_34/forx_xbody16_forx_xbody16_PhiReq/phi_stmt_107/phi_stmt_107_sources/type_cast_110/SplitProtocol/Update/ca
      -- 
    ca_2690_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 240_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_110_inst_ack_1, ack => testConfigure_CP_0_elements(240)); -- 
    -- CP-element group 241:  join  transition  output  bypass 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	239 
    -- CP-element group 241: 	240 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	243 
    -- CP-element group 241:  members (6) 
      -- CP-element group 241: 	 branch_block_stmt_34/forx_xbody16_forx_xbody16_PhiReq/$exit
      -- CP-element group 241: 	 branch_block_stmt_34/forx_xbody16_forx_xbody16_PhiReq/phi_stmt_107/$exit
      -- CP-element group 241: 	 branch_block_stmt_34/forx_xbody16_forx_xbody16_PhiReq/phi_stmt_107/phi_stmt_107_sources/$exit
      -- CP-element group 241: 	 branch_block_stmt_34/forx_xbody16_forx_xbody16_PhiReq/phi_stmt_107/phi_stmt_107_sources/type_cast_110/$exit
      -- CP-element group 241: 	 branch_block_stmt_34/forx_xbody16_forx_xbody16_PhiReq/phi_stmt_107/phi_stmt_107_sources/type_cast_110/SplitProtocol/$exit
      -- CP-element group 241: 	 branch_block_stmt_34/forx_xbody16_forx_xbody16_PhiReq/phi_stmt_107/phi_stmt_107_req
      -- 
    phi_stmt_107_req_2691_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_107_req_2691_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(241), ack => phi_stmt_107_req_0); -- 
    testConfigure_cp_element_group_241: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_241"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(239) & testConfigure_CP_0_elements(240);
      gj_testConfigure_cp_element_group_241 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(241), clk => clk, reset => reset); --
    end block;
    -- CP-element group 242:  transition  output  delay-element  bypass 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	21 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	243 
    -- CP-element group 242:  members (5) 
      -- CP-element group 242: 	 branch_block_stmt_34/forx_xbody16x_xpreheader_forx_xbody16_PhiReq/$exit
      -- CP-element group 242: 	 branch_block_stmt_34/forx_xbody16x_xpreheader_forx_xbody16_PhiReq/phi_stmt_107/$exit
      -- CP-element group 242: 	 branch_block_stmt_34/forx_xbody16x_xpreheader_forx_xbody16_PhiReq/phi_stmt_107/phi_stmt_107_sources/$exit
      -- CP-element group 242: 	 branch_block_stmt_34/forx_xbody16x_xpreheader_forx_xbody16_PhiReq/phi_stmt_107/phi_stmt_107_sources/type_cast_113_konst_delay_trans
      -- CP-element group 242: 	 branch_block_stmt_34/forx_xbody16x_xpreheader_forx_xbody16_PhiReq/phi_stmt_107/phi_stmt_107_req
      -- 
    phi_stmt_107_req_2702_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_107_req_2702_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(242), ack => phi_stmt_107_req_1); -- 
    -- Element group testConfigure_CP_0_elements(242) is a control-delay.
    cp_element_242_delay: control_delay_element  generic map(name => " 242_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(21), ack => testConfigure_CP_0_elements(242), clk => clk, reset =>reset);
    -- CP-element group 243:  merge  transition  place  bypass 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	241 
    -- CP-element group 243: 	242 
    -- CP-element group 243: successors 
    -- CP-element group 243: 	244 
    -- CP-element group 243:  members (2) 
      -- CP-element group 243: 	 branch_block_stmt_34/merge_stmt_106_PhiReqMerge
      -- CP-element group 243: 	 branch_block_stmt_34/merge_stmt_106_PhiAck/$entry
      -- 
    testConfigure_CP_0_elements(243) <= OrReduce(testConfigure_CP_0_elements(241) & testConfigure_CP_0_elements(242));
    -- CP-element group 244:  fork  transition  place  input  output  bypass 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	243 
    -- CP-element group 244: successors 
    -- CP-element group 244: 	30 
    -- CP-element group 244: 	27 
    -- CP-element group 244: 	33 
    -- CP-element group 244: 	37 
    -- CP-element group 244: 	40 
    -- CP-element group 244: 	23 
    -- CP-element group 244: 	24 
    -- CP-element group 244: 	26 
    -- CP-element group 244:  members (43) 
      -- CP-element group 244: 	 branch_block_stmt_34/merge_stmt_106__exit__
      -- CP-element group 244: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166__entry__
      -- CP-element group 244: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/array_obj_ref_119_index_scale_1/$entry
      -- CP-element group 244: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/array_obj_ref_119_index_scale_1/$exit
      -- CP-element group 244: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/array_obj_ref_119_index_scale_1/scale_rename_req
      -- CP-element group 244: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/array_obj_ref_119_index_scale_1/scale_rename_ack
      -- CP-element group 244: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/array_obj_ref_119_final_index_sum_regn_update_start
      -- CP-element group 244: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/array_obj_ref_119_final_index_sum_regn_Sample/$entry
      -- CP-element group 244: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/array_obj_ref_119_final_index_sum_regn_Sample/req
      -- CP-element group 244: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/array_obj_ref_119_final_index_sum_regn_Update/$entry
      -- CP-element group 244: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/array_obj_ref_119_final_index_sum_regn_Update/req
      -- CP-element group 244: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/$entry
      -- CP-element group 244: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/addr_of_120_update_start_
      -- CP-element group 244: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/array_obj_ref_119_index_resized_1
      -- CP-element group 244: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/array_obj_ref_119_index_scaled_1
      -- CP-element group 244: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/array_obj_ref_119_index_computed_1
      -- CP-element group 244: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/array_obj_ref_119_index_resize_1/$entry
      -- CP-element group 244: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/array_obj_ref_119_index_resize_1/$exit
      -- CP-element group 244: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/array_obj_ref_119_index_resize_1/index_resize_req
      -- CP-element group 244: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/array_obj_ref_119_index_resize_1/index_resize_ack
      -- CP-element group 244: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/addr_of_120_complete/$entry
      -- CP-element group 244: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/addr_of_120_complete/req
      -- CP-element group 244: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/RPIPE_ConvTranspose_input_pipe_123_sample_start_
      -- CP-element group 244: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/RPIPE_ConvTranspose_input_pipe_123_Sample/$entry
      -- CP-element group 244: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/RPIPE_ConvTranspose_input_pipe_123_Sample/rr
      -- CP-element group 244: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/type_cast_127_update_start_
      -- CP-element group 244: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/type_cast_127_Update/$entry
      -- CP-element group 244: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/type_cast_127_Update/cr
      -- CP-element group 244: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_130_update_start_
      -- CP-element group 244: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_130_Update/$entry
      -- CP-element group 244: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_130_Update/word_access_complete/$entry
      -- CP-element group 244: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_130_Update/word_access_complete/word_0/$entry
      -- CP-element group 244: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_130_Update/word_access_complete/word_0/cr
      -- CP-element group 244: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/type_cast_144_update_start_
      -- CP-element group 244: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/type_cast_144_Update/$entry
      -- CP-element group 244: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/type_cast_144_Update/cr
      -- CP-element group 244: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_152_update_start_
      -- CP-element group 244: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_152_Update/$entry
      -- CP-element group 244: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_152_Update/word_access_complete/$entry
      -- CP-element group 244: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_152_Update/word_access_complete/word_0/$entry
      -- CP-element group 244: 	 branch_block_stmt_34/assign_stmt_121_to_assign_stmt_166/ptr_deref_152_Update/word_access_complete/word_0/cr
      -- CP-element group 244: 	 branch_block_stmt_34/merge_stmt_106_PhiAck/$exit
      -- CP-element group 244: 	 branch_block_stmt_34/merge_stmt_106_PhiAck/phi_stmt_107_ack
      -- 
    phi_stmt_107_ack_2707_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 244_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_107_ack_0, ack => testConfigure_CP_0_elements(244)); -- 
    req_344_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_344_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(244), ack => array_obj_ref_119_index_offset_req_0); -- 
    req_349_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_349_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(244), ack => array_obj_ref_119_index_offset_req_1); -- 
    req_364_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_364_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(244), ack => addr_of_120_final_reg_req_1); -- 
    rr_373_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_373_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(244), ack => RPIPE_ConvTranspose_input_pipe_123_inst_req_0); -- 
    cr_392_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_392_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(244), ack => type_cast_127_inst_req_1); -- 
    cr_442_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_442_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(244), ack => ptr_deref_130_store_0_req_1); -- 
    cr_470_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_470_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(244), ack => type_cast_144_inst_req_1); -- 
    cr_520_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_520_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(244), ack => ptr_deref_152_store_0_req_1); -- 
    -- CP-element group 245:  transition  output  delay-element  bypass 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	46 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	249 
    -- CP-element group 245:  members (4) 
      -- CP-element group 245: 	 branch_block_stmt_34/bbx_xnph240_forx_xbody41_PhiReq/phi_stmt_179/$exit
      -- CP-element group 245: 	 branch_block_stmt_34/bbx_xnph240_forx_xbody41_PhiReq/phi_stmt_179/phi_stmt_179_sources/$exit
      -- CP-element group 245: 	 branch_block_stmt_34/bbx_xnph240_forx_xbody41_PhiReq/phi_stmt_179/phi_stmt_179_sources/type_cast_183_konst_delay_trans
      -- CP-element group 245: 	 branch_block_stmt_34/bbx_xnph240_forx_xbody41_PhiReq/phi_stmt_179/phi_stmt_179_req
      -- 
    phi_stmt_179_req_2730_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_179_req_2730_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(245), ack => phi_stmt_179_req_0); -- 
    -- Element group testConfigure_CP_0_elements(245) is a control-delay.
    cp_element_245_delay: control_delay_element  generic map(name => " 245_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(46), ack => testConfigure_CP_0_elements(245), clk => clk, reset =>reset);
    -- CP-element group 246:  transition  input  bypass 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	46 
    -- CP-element group 246: successors 
    -- CP-element group 246: 	248 
    -- CP-element group 246:  members (2) 
      -- CP-element group 246: 	 branch_block_stmt_34/bbx_xnph240_forx_xbody41_PhiReq/phi_stmt_186/phi_stmt_186_sources/type_cast_189/SplitProtocol/Sample/$exit
      -- CP-element group 246: 	 branch_block_stmt_34/bbx_xnph240_forx_xbody41_PhiReq/phi_stmt_186/phi_stmt_186_sources/type_cast_189/SplitProtocol/Sample/ra
      -- 
    ra_2747_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 246_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_189_inst_ack_0, ack => testConfigure_CP_0_elements(246)); -- 
    -- CP-element group 247:  transition  input  bypass 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	46 
    -- CP-element group 247: successors 
    -- CP-element group 247: 	248 
    -- CP-element group 247:  members (2) 
      -- CP-element group 247: 	 branch_block_stmt_34/bbx_xnph240_forx_xbody41_PhiReq/phi_stmt_186/phi_stmt_186_sources/type_cast_189/SplitProtocol/Update/$exit
      -- CP-element group 247: 	 branch_block_stmt_34/bbx_xnph240_forx_xbody41_PhiReq/phi_stmt_186/phi_stmt_186_sources/type_cast_189/SplitProtocol/Update/ca
      -- 
    ca_2752_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 247_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_189_inst_ack_1, ack => testConfigure_CP_0_elements(247)); -- 
    -- CP-element group 248:  join  transition  output  bypass 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	246 
    -- CP-element group 248: 	247 
    -- CP-element group 248: successors 
    -- CP-element group 248: 	249 
    -- CP-element group 248:  members (5) 
      -- CP-element group 248: 	 branch_block_stmt_34/bbx_xnph240_forx_xbody41_PhiReq/phi_stmt_186/$exit
      -- CP-element group 248: 	 branch_block_stmt_34/bbx_xnph240_forx_xbody41_PhiReq/phi_stmt_186/phi_stmt_186_sources/$exit
      -- CP-element group 248: 	 branch_block_stmt_34/bbx_xnph240_forx_xbody41_PhiReq/phi_stmt_186/phi_stmt_186_sources/type_cast_189/$exit
      -- CP-element group 248: 	 branch_block_stmt_34/bbx_xnph240_forx_xbody41_PhiReq/phi_stmt_186/phi_stmt_186_sources/type_cast_189/SplitProtocol/$exit
      -- CP-element group 248: 	 branch_block_stmt_34/bbx_xnph240_forx_xbody41_PhiReq/phi_stmt_186/phi_stmt_186_req
      -- 
    phi_stmt_186_req_2753_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_186_req_2753_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(248), ack => phi_stmt_186_req_0); -- 
    testConfigure_cp_element_group_248: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_248"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(246) & testConfigure_CP_0_elements(247);
      gj_testConfigure_cp_element_group_248 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(248), clk => clk, reset => reset); --
    end block;
    -- CP-element group 249:  join  transition  bypass 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	245 
    -- CP-element group 249: 	248 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	257 
    -- CP-element group 249:  members (1) 
      -- CP-element group 249: 	 branch_block_stmt_34/bbx_xnph240_forx_xbody41_PhiReq/$exit
      -- 
    testConfigure_cp_element_group_249: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_249"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(245) & testConfigure_CP_0_elements(248);
      gj_testConfigure_cp_element_group_249 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(249), clk => clk, reset => reset); --
    end block;
    -- CP-element group 250:  transition  input  bypass 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	55 
    -- CP-element group 250: successors 
    -- CP-element group 250: 	252 
    -- CP-element group 250:  members (2) 
      -- CP-element group 250: 	 branch_block_stmt_34/forx_xbody41_forx_xbody41_PhiReq/phi_stmt_179/phi_stmt_179_sources/type_cast_185/SplitProtocol/Sample/$exit
      -- CP-element group 250: 	 branch_block_stmt_34/forx_xbody41_forx_xbody41_PhiReq/phi_stmt_179/phi_stmt_179_sources/type_cast_185/SplitProtocol/Sample/ra
      -- 
    ra_2773_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 250_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_185_inst_ack_0, ack => testConfigure_CP_0_elements(250)); -- 
    -- CP-element group 251:  transition  input  bypass 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	55 
    -- CP-element group 251: successors 
    -- CP-element group 251: 	252 
    -- CP-element group 251:  members (2) 
      -- CP-element group 251: 	 branch_block_stmt_34/forx_xbody41_forx_xbody41_PhiReq/phi_stmt_179/phi_stmt_179_sources/type_cast_185/SplitProtocol/Update/$exit
      -- CP-element group 251: 	 branch_block_stmt_34/forx_xbody41_forx_xbody41_PhiReq/phi_stmt_179/phi_stmt_179_sources/type_cast_185/SplitProtocol/Update/ca
      -- 
    ca_2778_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 251_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_185_inst_ack_1, ack => testConfigure_CP_0_elements(251)); -- 
    -- CP-element group 252:  join  transition  output  bypass 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	250 
    -- CP-element group 252: 	251 
    -- CP-element group 252: successors 
    -- CP-element group 252: 	256 
    -- CP-element group 252:  members (5) 
      -- CP-element group 252: 	 branch_block_stmt_34/forx_xbody41_forx_xbody41_PhiReq/phi_stmt_179/$exit
      -- CP-element group 252: 	 branch_block_stmt_34/forx_xbody41_forx_xbody41_PhiReq/phi_stmt_179/phi_stmt_179_sources/$exit
      -- CP-element group 252: 	 branch_block_stmt_34/forx_xbody41_forx_xbody41_PhiReq/phi_stmt_179/phi_stmt_179_sources/type_cast_185/$exit
      -- CP-element group 252: 	 branch_block_stmt_34/forx_xbody41_forx_xbody41_PhiReq/phi_stmt_179/phi_stmt_179_sources/type_cast_185/SplitProtocol/$exit
      -- CP-element group 252: 	 branch_block_stmt_34/forx_xbody41_forx_xbody41_PhiReq/phi_stmt_179/phi_stmt_179_req
      -- 
    phi_stmt_179_req_2779_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_179_req_2779_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(252), ack => phi_stmt_179_req_1); -- 
    testConfigure_cp_element_group_252: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_252"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(250) & testConfigure_CP_0_elements(251);
      gj_testConfigure_cp_element_group_252 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(252), clk => clk, reset => reset); --
    end block;
    -- CP-element group 253:  transition  input  bypass 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	55 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	255 
    -- CP-element group 253:  members (2) 
      -- CP-element group 253: 	 branch_block_stmt_34/forx_xbody41_forx_xbody41_PhiReq/phi_stmt_186/phi_stmt_186_sources/type_cast_191/SplitProtocol/Sample/$exit
      -- CP-element group 253: 	 branch_block_stmt_34/forx_xbody41_forx_xbody41_PhiReq/phi_stmt_186/phi_stmt_186_sources/type_cast_191/SplitProtocol/Sample/ra
      -- 
    ra_2796_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 253_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_191_inst_ack_0, ack => testConfigure_CP_0_elements(253)); -- 
    -- CP-element group 254:  transition  input  bypass 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	55 
    -- CP-element group 254: successors 
    -- CP-element group 254: 	255 
    -- CP-element group 254:  members (2) 
      -- CP-element group 254: 	 branch_block_stmt_34/forx_xbody41_forx_xbody41_PhiReq/phi_stmt_186/phi_stmt_186_sources/type_cast_191/SplitProtocol/Update/$exit
      -- CP-element group 254: 	 branch_block_stmt_34/forx_xbody41_forx_xbody41_PhiReq/phi_stmt_186/phi_stmt_186_sources/type_cast_191/SplitProtocol/Update/ca
      -- 
    ca_2801_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 254_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_191_inst_ack_1, ack => testConfigure_CP_0_elements(254)); -- 
    -- CP-element group 255:  join  transition  output  bypass 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	253 
    -- CP-element group 255: 	254 
    -- CP-element group 255: successors 
    -- CP-element group 255: 	256 
    -- CP-element group 255:  members (5) 
      -- CP-element group 255: 	 branch_block_stmt_34/forx_xbody41_forx_xbody41_PhiReq/phi_stmt_186/$exit
      -- CP-element group 255: 	 branch_block_stmt_34/forx_xbody41_forx_xbody41_PhiReq/phi_stmt_186/phi_stmt_186_sources/$exit
      -- CP-element group 255: 	 branch_block_stmt_34/forx_xbody41_forx_xbody41_PhiReq/phi_stmt_186/phi_stmt_186_sources/type_cast_191/$exit
      -- CP-element group 255: 	 branch_block_stmt_34/forx_xbody41_forx_xbody41_PhiReq/phi_stmt_186/phi_stmt_186_sources/type_cast_191/SplitProtocol/$exit
      -- CP-element group 255: 	 branch_block_stmt_34/forx_xbody41_forx_xbody41_PhiReq/phi_stmt_186/phi_stmt_186_req
      -- 
    phi_stmt_186_req_2802_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_186_req_2802_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(255), ack => phi_stmt_186_req_1); -- 
    testConfigure_cp_element_group_255: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_255"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(253) & testConfigure_CP_0_elements(254);
      gj_testConfigure_cp_element_group_255 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(255), clk => clk, reset => reset); --
    end block;
    -- CP-element group 256:  join  transition  bypass 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	252 
    -- CP-element group 256: 	255 
    -- CP-element group 256: successors 
    -- CP-element group 256: 	257 
    -- CP-element group 256:  members (1) 
      -- CP-element group 256: 	 branch_block_stmt_34/forx_xbody41_forx_xbody41_PhiReq/$exit
      -- 
    testConfigure_cp_element_group_256: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_256"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(252) & testConfigure_CP_0_elements(255);
      gj_testConfigure_cp_element_group_256 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(256), clk => clk, reset => reset); --
    end block;
    -- CP-element group 257:  merge  fork  transition  place  bypass 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	249 
    -- CP-element group 257: 	256 
    -- CP-element group 257: successors 
    -- CP-element group 257: 	258 
    -- CP-element group 257: 	259 
    -- CP-element group 257:  members (2) 
      -- CP-element group 257: 	 branch_block_stmt_34/merge_stmt_178_PhiReqMerge
      -- CP-element group 257: 	 branch_block_stmt_34/merge_stmt_178_PhiAck/$entry
      -- 
    testConfigure_CP_0_elements(257) <= OrReduce(testConfigure_CP_0_elements(249) & testConfigure_CP_0_elements(256));
    -- CP-element group 258:  transition  input  bypass 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	257 
    -- CP-element group 258: successors 
    -- CP-element group 258: 	260 
    -- CP-element group 258:  members (1) 
      -- CP-element group 258: 	 branch_block_stmt_34/merge_stmt_178_PhiAck/phi_stmt_179_ack
      -- 
    phi_stmt_179_ack_2807_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 258_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_179_ack_0, ack => testConfigure_CP_0_elements(258)); -- 
    -- CP-element group 259:  transition  input  bypass 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	257 
    -- CP-element group 259: successors 
    -- CP-element group 259: 	260 
    -- CP-element group 259:  members (1) 
      -- CP-element group 259: 	 branch_block_stmt_34/merge_stmt_178_PhiAck/phi_stmt_186_ack
      -- 
    phi_stmt_186_ack_2808_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 259_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_186_ack_0, ack => testConfigure_CP_0_elements(259)); -- 
    -- CP-element group 260:  join  fork  transition  place  output  bypass 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	258 
    -- CP-element group 260: 	259 
    -- CP-element group 260: successors 
    -- CP-element group 260: 	51 
    -- CP-element group 260: 	50 
    -- CP-element group 260: 	47 
    -- CP-element group 260: 	48 
    -- CP-element group 260:  members (39) 
      -- CP-element group 260: 	 branch_block_stmt_34/merge_stmt_178__exit__
      -- CP-element group 260: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216__entry__
      -- CP-element group 260: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/$entry
      -- CP-element group 260: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/addr_of_196_sample_start_
      -- CP-element group 260: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/addr_of_196_update_start_
      -- CP-element group 260: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/array_obj_ref_195_root_address_calculated
      -- CP-element group 260: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/array_obj_ref_195_offset_calculated
      -- CP-element group 260: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/array_obj_ref_195_index_resized_0
      -- CP-element group 260: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/array_obj_ref_195_index_scaled_0
      -- CP-element group 260: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/array_obj_ref_195_index_computed_0
      -- CP-element group 260: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/array_obj_ref_195_index_resize_0/$entry
      -- CP-element group 260: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/array_obj_ref_195_index_resize_0/$exit
      -- CP-element group 260: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/array_obj_ref_195_index_resize_0/index_resize_req
      -- CP-element group 260: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/array_obj_ref_195_index_resize_0/index_resize_ack
      -- CP-element group 260: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/array_obj_ref_195_index_scale_0/$entry
      -- CP-element group 260: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/array_obj_ref_195_index_scale_0/$exit
      -- CP-element group 260: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/array_obj_ref_195_index_scale_0/scale_rename_req
      -- CP-element group 260: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/array_obj_ref_195_index_scale_0/scale_rename_ack
      -- CP-element group 260: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/array_obj_ref_195_final_index_sum_regn/$entry
      -- CP-element group 260: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/array_obj_ref_195_final_index_sum_regn/$exit
      -- CP-element group 260: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/array_obj_ref_195_final_index_sum_regn/req
      -- CP-element group 260: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/array_obj_ref_195_final_index_sum_regn/ack
      -- CP-element group 260: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/array_obj_ref_195_base_plus_offset/$entry
      -- CP-element group 260: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/array_obj_ref_195_base_plus_offset/$exit
      -- CP-element group 260: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/array_obj_ref_195_base_plus_offset/sum_rename_req
      -- CP-element group 260: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/array_obj_ref_195_base_plus_offset/sum_rename_ack
      -- CP-element group 260: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/addr_of_196_request/$entry
      -- CP-element group 260: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/addr_of_196_request/req
      -- CP-element group 260: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/addr_of_196_complete/$entry
      -- CP-element group 260: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/addr_of_196_complete/req
      -- CP-element group 260: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/ptr_deref_199_update_start_
      -- CP-element group 260: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/ptr_deref_199_Update/$entry
      -- CP-element group 260: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/ptr_deref_199_Update/word_access_complete/$entry
      -- CP-element group 260: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/ptr_deref_199_Update/word_access_complete/word_0/$entry
      -- CP-element group 260: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/ptr_deref_199_Update/word_access_complete/word_0/cr
      -- CP-element group 260: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/RPIPE_ConvTranspose_input_pipe_203_sample_start_
      -- CP-element group 260: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/RPIPE_ConvTranspose_input_pipe_203_Sample/$entry
      -- CP-element group 260: 	 branch_block_stmt_34/assign_stmt_197_to_assign_stmt_216/RPIPE_ConvTranspose_input_pipe_203_Sample/rr
      -- CP-element group 260: 	 branch_block_stmt_34/merge_stmt_178_PhiAck/$exit
      -- 
    req_594_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_594_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(260), ack => addr_of_196_final_reg_req_0); -- 
    req_599_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_599_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(260), ack => addr_of_196_final_reg_req_1); -- 
    cr_649_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_649_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(260), ack => ptr_deref_199_store_0_req_1); -- 
    rr_658_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_658_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(260), ack => RPIPE_ConvTranspose_input_pipe_203_inst_req_0); -- 
    testConfigure_cp_element_group_260: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_260"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(258) & testConfigure_CP_0_elements(259);
      gj_testConfigure_cp_element_group_260 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(260), clk => clk, reset => reset); --
    end block;
    -- CP-element group 261:  transition  input  bypass 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	54 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	263 
    -- CP-element group 261:  members (2) 
      -- CP-element group 261: 	 branch_block_stmt_34/forx_xbody41_forx_xend49_PhiReq/phi_stmt_224/phi_stmt_224_sources/type_cast_227/SplitProtocol/Sample/$exit
      -- CP-element group 261: 	 branch_block_stmt_34/forx_xbody41_forx_xend49_PhiReq/phi_stmt_224/phi_stmt_224_sources/type_cast_227/SplitProtocol/Sample/ra
      -- 
    ra_2832_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 261_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_227_inst_ack_0, ack => testConfigure_CP_0_elements(261)); -- 
    -- CP-element group 262:  transition  input  bypass 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	54 
    -- CP-element group 262: successors 
    -- CP-element group 262: 	263 
    -- CP-element group 262:  members (2) 
      -- CP-element group 262: 	 branch_block_stmt_34/forx_xbody41_forx_xend49_PhiReq/phi_stmt_224/phi_stmt_224_sources/type_cast_227/SplitProtocol/Update/$exit
      -- CP-element group 262: 	 branch_block_stmt_34/forx_xbody41_forx_xend49_PhiReq/phi_stmt_224/phi_stmt_224_sources/type_cast_227/SplitProtocol/Update/ca
      -- 
    ca_2837_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 262_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_227_inst_ack_1, ack => testConfigure_CP_0_elements(262)); -- 
    -- CP-element group 263:  join  transition  place  output  bypass 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	261 
    -- CP-element group 263: 	262 
    -- CP-element group 263: successors 
    -- CP-element group 263: 	264 
    -- CP-element group 263:  members (8) 
      -- CP-element group 263: 	 branch_block_stmt_34/forx_xbody41_forx_xend49_PhiReq/$exit
      -- CP-element group 263: 	 branch_block_stmt_34/forx_xbody41_forx_xend49_PhiReq/phi_stmt_224/$exit
      -- CP-element group 263: 	 branch_block_stmt_34/forx_xbody41_forx_xend49_PhiReq/phi_stmt_224/phi_stmt_224_sources/$exit
      -- CP-element group 263: 	 branch_block_stmt_34/forx_xbody41_forx_xend49_PhiReq/phi_stmt_224/phi_stmt_224_sources/type_cast_227/$exit
      -- CP-element group 263: 	 branch_block_stmt_34/forx_xbody41_forx_xend49_PhiReq/phi_stmt_224/phi_stmt_224_sources/type_cast_227/SplitProtocol/$exit
      -- CP-element group 263: 	 branch_block_stmt_34/forx_xbody41_forx_xend49_PhiReq/phi_stmt_224/phi_stmt_224_req
      -- CP-element group 263: 	 branch_block_stmt_34/merge_stmt_223_PhiReqMerge
      -- CP-element group 263: 	 branch_block_stmt_34/merge_stmt_223_PhiAck/$entry
      -- 
    phi_stmt_224_req_2838_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_224_req_2838_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(263), ack => phi_stmt_224_req_0); -- 
    testConfigure_cp_element_group_263: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_263"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(261) & testConfigure_CP_0_elements(262);
      gj_testConfigure_cp_element_group_263 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(263), clk => clk, reset => reset); --
    end block;
    -- CP-element group 264:  merge  transition  place  input  bypass 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	263 
    -- CP-element group 264: successors 
    -- CP-element group 264: 	56 
    -- CP-element group 264:  members (4) 
      -- CP-element group 264: 	 branch_block_stmt_34/merge_stmt_223__exit__
      -- CP-element group 264: 	 branch_block_stmt_34/assign_stmt_231_to_assign_stmt_493__entry__
      -- CP-element group 264: 	 branch_block_stmt_34/merge_stmt_223_PhiAck/$exit
      -- CP-element group 264: 	 branch_block_stmt_34/merge_stmt_223_PhiAck/phi_stmt_224_ack
      -- 
    phi_stmt_224_ack_2843_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 264_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_224_ack_0, ack => testConfigure_CP_0_elements(264)); -- 
    -- CP-element group 265:  merge  branch  transition  place  output  bypass 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	122 
    -- CP-element group 265: 	167 
    -- CP-element group 265: successors 
    -- CP-element group 265: 	123 
    -- CP-element group 265: 	124 
    -- CP-element group 265:  members (17) 
      -- CP-element group 265: 	 branch_block_stmt_34/merge_stmt_502__exit__
      -- CP-element group 265: 	 branch_block_stmt_34/assign_stmt_508__entry__
      -- CP-element group 265: 	 branch_block_stmt_34/assign_stmt_508__exit__
      -- CP-element group 265: 	 branch_block_stmt_34/if_stmt_509__entry__
      -- CP-element group 265: 	 branch_block_stmt_34/assign_stmt_508/$entry
      -- CP-element group 265: 	 branch_block_stmt_34/assign_stmt_508/$exit
      -- CP-element group 265: 	 branch_block_stmt_34/if_stmt_509_dead_link/$entry
      -- CP-element group 265: 	 branch_block_stmt_34/if_stmt_509_eval_test/$entry
      -- CP-element group 265: 	 branch_block_stmt_34/if_stmt_509_eval_test/$exit
      -- CP-element group 265: 	 branch_block_stmt_34/if_stmt_509_eval_test/branch_req
      -- CP-element group 265: 	 branch_block_stmt_34/R_cmp148229_510_place
      -- CP-element group 265: 	 branch_block_stmt_34/if_stmt_509_if_link/$entry
      -- CP-element group 265: 	 branch_block_stmt_34/if_stmt_509_else_link/$entry
      -- CP-element group 265: 	 branch_block_stmt_34/merge_stmt_502_PhiReqMerge
      -- CP-element group 265: 	 branch_block_stmt_34/merge_stmt_502_PhiAck/$entry
      -- CP-element group 265: 	 branch_block_stmt_34/merge_stmt_502_PhiAck/$exit
      -- CP-element group 265: 	 branch_block_stmt_34/merge_stmt_502_PhiAck/dummy
      -- 
    branch_req_1572_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1572_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(265), ack => if_stmt_509_branch_req_0); -- 
    testConfigure_CP_0_elements(265) <= OrReduce(testConfigure_CP_0_elements(122) & testConfigure_CP_0_elements(167));
    -- CP-element group 266:  transition  output  delay-element  bypass 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	126 
    -- CP-element group 266: successors 
    -- CP-element group 266: 	270 
    -- CP-element group 266:  members (5) 
      -- CP-element group 266: 	 branch_block_stmt_34/bbx_xnph235_forx_xbody90_PhiReq/$exit
      -- CP-element group 266: 	 branch_block_stmt_34/bbx_xnph235_forx_xbody90_PhiReq/phi_stmt_553/$exit
      -- CP-element group 266: 	 branch_block_stmt_34/bbx_xnph235_forx_xbody90_PhiReq/phi_stmt_553/phi_stmt_553_sources/$exit
      -- CP-element group 266: 	 branch_block_stmt_34/bbx_xnph235_forx_xbody90_PhiReq/phi_stmt_553/phi_stmt_553_sources/type_cast_557_konst_delay_trans
      -- CP-element group 266: 	 branch_block_stmt_34/bbx_xnph235_forx_xbody90_PhiReq/phi_stmt_553/phi_stmt_553_req
      -- 
    phi_stmt_553_req_2889_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_553_req_2889_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(266), ack => phi_stmt_553_req_0); -- 
    -- Element group testConfigure_CP_0_elements(266) is a control-delay.
    cp_element_266_delay: control_delay_element  generic map(name => " 266_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(126), ack => testConfigure_CP_0_elements(266), clk => clk, reset =>reset);
    -- CP-element group 267:  transition  input  bypass 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	168 
    -- CP-element group 267: successors 
    -- CP-element group 267: 	269 
    -- CP-element group 267:  members (2) 
      -- CP-element group 267: 	 branch_block_stmt_34/forx_xbody90_forx_xbody90_PhiReq/phi_stmt_553/phi_stmt_553_sources/type_cast_559/SplitProtocol/Sample/$exit
      -- CP-element group 267: 	 branch_block_stmt_34/forx_xbody90_forx_xbody90_PhiReq/phi_stmt_553/phi_stmt_553_sources/type_cast_559/SplitProtocol/Sample/ra
      -- 
    ra_2909_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 267_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_559_inst_ack_0, ack => testConfigure_CP_0_elements(267)); -- 
    -- CP-element group 268:  transition  input  bypass 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	168 
    -- CP-element group 268: successors 
    -- CP-element group 268: 	269 
    -- CP-element group 268:  members (2) 
      -- CP-element group 268: 	 branch_block_stmt_34/forx_xbody90_forx_xbody90_PhiReq/phi_stmt_553/phi_stmt_553_sources/type_cast_559/SplitProtocol/Update/$exit
      -- CP-element group 268: 	 branch_block_stmt_34/forx_xbody90_forx_xbody90_PhiReq/phi_stmt_553/phi_stmt_553_sources/type_cast_559/SplitProtocol/Update/ca
      -- 
    ca_2914_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 268_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_559_inst_ack_1, ack => testConfigure_CP_0_elements(268)); -- 
    -- CP-element group 269:  join  transition  output  bypass 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: 	267 
    -- CP-element group 269: 	268 
    -- CP-element group 269: successors 
    -- CP-element group 269: 	270 
    -- CP-element group 269:  members (6) 
      -- CP-element group 269: 	 branch_block_stmt_34/forx_xbody90_forx_xbody90_PhiReq/$exit
      -- CP-element group 269: 	 branch_block_stmt_34/forx_xbody90_forx_xbody90_PhiReq/phi_stmt_553/$exit
      -- CP-element group 269: 	 branch_block_stmt_34/forx_xbody90_forx_xbody90_PhiReq/phi_stmt_553/phi_stmt_553_sources/$exit
      -- CP-element group 269: 	 branch_block_stmt_34/forx_xbody90_forx_xbody90_PhiReq/phi_stmt_553/phi_stmt_553_sources/type_cast_559/$exit
      -- CP-element group 269: 	 branch_block_stmt_34/forx_xbody90_forx_xbody90_PhiReq/phi_stmt_553/phi_stmt_553_sources/type_cast_559/SplitProtocol/$exit
      -- CP-element group 269: 	 branch_block_stmt_34/forx_xbody90_forx_xbody90_PhiReq/phi_stmt_553/phi_stmt_553_req
      -- 
    phi_stmt_553_req_2915_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_553_req_2915_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(269), ack => phi_stmt_553_req_1); -- 
    testConfigure_cp_element_group_269: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_269"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(267) & testConfigure_CP_0_elements(268);
      gj_testConfigure_cp_element_group_269 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(269), clk => clk, reset => reset); --
    end block;
    -- CP-element group 270:  merge  transition  place  bypass 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	266 
    -- CP-element group 270: 	269 
    -- CP-element group 270: successors 
    -- CP-element group 270: 	271 
    -- CP-element group 270:  members (2) 
      -- CP-element group 270: 	 branch_block_stmt_34/merge_stmt_552_PhiReqMerge
      -- CP-element group 270: 	 branch_block_stmt_34/merge_stmt_552_PhiAck/$entry
      -- 
    testConfigure_CP_0_elements(270) <= OrReduce(testConfigure_CP_0_elements(266) & testConfigure_CP_0_elements(269));
    -- CP-element group 271:  fork  transition  place  input  output  bypass 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	270 
    -- CP-element group 271: successors 
    -- CP-element group 271: 	127 
    -- CP-element group 271: 	128 
    -- CP-element group 271: 	130 
    -- CP-element group 271: 	131 
    -- CP-element group 271: 	134 
    -- CP-element group 271: 	138 
    -- CP-element group 271: 	142 
    -- CP-element group 271: 	146 
    -- CP-element group 271: 	150 
    -- CP-element group 271: 	154 
    -- CP-element group 271: 	158 
    -- CP-element group 271: 	162 
    -- CP-element group 271: 	165 
    -- CP-element group 271:  members (56) 
      -- CP-element group 271: 	 branch_block_stmt_34/merge_stmt_552__exit__
      -- CP-element group 271: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715__entry__
      -- CP-element group 271: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/$entry
      -- CP-element group 271: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/addr_of_566_update_start_
      -- CP-element group 271: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/array_obj_ref_565_index_resized_1
      -- CP-element group 271: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/array_obj_ref_565_index_scaled_1
      -- CP-element group 271: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/array_obj_ref_565_index_computed_1
      -- CP-element group 271: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/array_obj_ref_565_index_resize_1/$entry
      -- CP-element group 271: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/array_obj_ref_565_index_resize_1/$exit
      -- CP-element group 271: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/array_obj_ref_565_index_resize_1/index_resize_req
      -- CP-element group 271: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/array_obj_ref_565_index_resize_1/index_resize_ack
      -- CP-element group 271: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/array_obj_ref_565_index_scale_1/$entry
      -- CP-element group 271: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/array_obj_ref_565_index_scale_1/$exit
      -- CP-element group 271: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/array_obj_ref_565_index_scale_1/scale_rename_req
      -- CP-element group 271: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/array_obj_ref_565_index_scale_1/scale_rename_ack
      -- CP-element group 271: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/array_obj_ref_565_final_index_sum_regn_update_start
      -- CP-element group 271: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/array_obj_ref_565_final_index_sum_regn_Sample/$entry
      -- CP-element group 271: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/array_obj_ref_565_final_index_sum_regn_Sample/req
      -- CP-element group 271: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/array_obj_ref_565_final_index_sum_regn_Update/$entry
      -- CP-element group 271: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/array_obj_ref_565_final_index_sum_regn_Update/req
      -- CP-element group 271: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/addr_of_566_complete/$entry
      -- CP-element group 271: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/addr_of_566_complete/req
      -- CP-element group 271: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_569_sample_start_
      -- CP-element group 271: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_569_Sample/$entry
      -- CP-element group 271: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/RPIPE_ConvTranspose_input_pipe_569_Sample/rr
      -- CP-element group 271: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_573_update_start_
      -- CP-element group 271: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_573_Update/$entry
      -- CP-element group 271: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_573_Update/cr
      -- CP-element group 271: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_586_update_start_
      -- CP-element group 271: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_586_Update/$entry
      -- CP-element group 271: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_586_Update/cr
      -- CP-element group 271: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_604_update_start_
      -- CP-element group 271: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_604_Update/$entry
      -- CP-element group 271: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_604_Update/cr
      -- CP-element group 271: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_622_update_start_
      -- CP-element group 271: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_622_Update/$entry
      -- CP-element group 271: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_622_Update/cr
      -- CP-element group 271: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_640_update_start_
      -- CP-element group 271: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_640_Update/$entry
      -- CP-element group 271: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_640_Update/cr
      -- CP-element group 271: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_658_update_start_
      -- CP-element group 271: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_658_Update/$entry
      -- CP-element group 271: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_658_Update/cr
      -- CP-element group 271: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_676_update_start_
      -- CP-element group 271: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_676_Update/$entry
      -- CP-element group 271: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_676_Update/cr
      -- CP-element group 271: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_694_update_start_
      -- CP-element group 271: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_694_Update/$entry
      -- CP-element group 271: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/type_cast_694_Update/cr
      -- CP-element group 271: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/ptr_deref_702_update_start_
      -- CP-element group 271: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/ptr_deref_702_Update/$entry
      -- CP-element group 271: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/ptr_deref_702_Update/word_access_complete/$entry
      -- CP-element group 271: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/ptr_deref_702_Update/word_access_complete/word_0/$entry
      -- CP-element group 271: 	 branch_block_stmt_34/assign_stmt_567_to_assign_stmt_715/ptr_deref_702_Update/word_access_complete/word_0/cr
      -- CP-element group 271: 	 branch_block_stmt_34/merge_stmt_552_PhiAck/$exit
      -- CP-element group 271: 	 branch_block_stmt_34/merge_stmt_552_PhiAck/phi_stmt_553_ack
      -- 
    phi_stmt_553_ack_2920_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 271_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_553_ack_0, ack => testConfigure_CP_0_elements(271)); -- 
    req_1628_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1628_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(271), ack => array_obj_ref_565_index_offset_req_0); -- 
    req_1633_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1633_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(271), ack => array_obj_ref_565_index_offset_req_1); -- 
    req_1648_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1648_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(271), ack => addr_of_566_final_reg_req_1); -- 
    rr_1657_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1657_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(271), ack => RPIPE_ConvTranspose_input_pipe_569_inst_req_0); -- 
    cr_1676_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1676_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(271), ack => type_cast_573_inst_req_1); -- 
    cr_1704_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1704_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(271), ack => type_cast_586_inst_req_1); -- 
    cr_1732_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1732_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(271), ack => type_cast_604_inst_req_1); -- 
    cr_1760_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1760_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(271), ack => type_cast_622_inst_req_1); -- 
    cr_1788_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1788_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(271), ack => type_cast_640_inst_req_1); -- 
    cr_1816_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1816_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(271), ack => type_cast_658_inst_req_1); -- 
    cr_1844_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1844_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(271), ack => type_cast_676_inst_req_1); -- 
    cr_1872_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1872_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(271), ack => type_cast_694_inst_req_1); -- 
    cr_1922_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1922_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(271), ack => ptr_deref_702_store_0_req_1); -- 
    -- CP-element group 272:  transition  output  delay-element  bypass 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	170 
    -- CP-element group 272: successors 
    -- CP-element group 272: 	276 
    -- CP-element group 272:  members (5) 
      -- CP-element group 272: 	 branch_block_stmt_34/bbx_xnph231_forx_xbody150_PhiReq/$exit
      -- CP-element group 272: 	 branch_block_stmt_34/bbx_xnph231_forx_xbody150_PhiReq/phi_stmt_760/$exit
      -- CP-element group 272: 	 branch_block_stmt_34/bbx_xnph231_forx_xbody150_PhiReq/phi_stmt_760/phi_stmt_760_sources/$exit
      -- CP-element group 272: 	 branch_block_stmt_34/bbx_xnph231_forx_xbody150_PhiReq/phi_stmt_760/phi_stmt_760_sources/type_cast_764_konst_delay_trans
      -- CP-element group 272: 	 branch_block_stmt_34/bbx_xnph231_forx_xbody150_PhiReq/phi_stmt_760/phi_stmt_760_req
      -- 
    phi_stmt_760_req_2943_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_760_req_2943_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(272), ack => phi_stmt_760_req_0); -- 
    -- Element group testConfigure_CP_0_elements(272) is a control-delay.
    cp_element_272_delay: control_delay_element  generic map(name => " 272_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(170), ack => testConfigure_CP_0_elements(272), clk => clk, reset =>reset);
    -- CP-element group 273:  transition  input  bypass 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: 	212 
    -- CP-element group 273: successors 
    -- CP-element group 273: 	275 
    -- CP-element group 273:  members (2) 
      -- CP-element group 273: 	 branch_block_stmt_34/forx_xbody150_forx_xbody150_PhiReq/phi_stmt_760/phi_stmt_760_sources/type_cast_766/SplitProtocol/Sample/$exit
      -- CP-element group 273: 	 branch_block_stmt_34/forx_xbody150_forx_xbody150_PhiReq/phi_stmt_760/phi_stmt_760_sources/type_cast_766/SplitProtocol/Sample/ra
      -- 
    ra_2963_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 273_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_766_inst_ack_0, ack => testConfigure_CP_0_elements(273)); -- 
    -- CP-element group 274:  transition  input  bypass 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	212 
    -- CP-element group 274: successors 
    -- CP-element group 274: 	275 
    -- CP-element group 274:  members (2) 
      -- CP-element group 274: 	 branch_block_stmt_34/forx_xbody150_forx_xbody150_PhiReq/phi_stmt_760/phi_stmt_760_sources/type_cast_766/SplitProtocol/Update/$exit
      -- CP-element group 274: 	 branch_block_stmt_34/forx_xbody150_forx_xbody150_PhiReq/phi_stmt_760/phi_stmt_760_sources/type_cast_766/SplitProtocol/Update/ca
      -- 
    ca_2968_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 274_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_766_inst_ack_1, ack => testConfigure_CP_0_elements(274)); -- 
    -- CP-element group 275:  join  transition  output  bypass 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	273 
    -- CP-element group 275: 	274 
    -- CP-element group 275: successors 
    -- CP-element group 275: 	276 
    -- CP-element group 275:  members (6) 
      -- CP-element group 275: 	 branch_block_stmt_34/forx_xbody150_forx_xbody150_PhiReq/$exit
      -- CP-element group 275: 	 branch_block_stmt_34/forx_xbody150_forx_xbody150_PhiReq/phi_stmt_760/$exit
      -- CP-element group 275: 	 branch_block_stmt_34/forx_xbody150_forx_xbody150_PhiReq/phi_stmt_760/phi_stmt_760_sources/$exit
      -- CP-element group 275: 	 branch_block_stmt_34/forx_xbody150_forx_xbody150_PhiReq/phi_stmt_760/phi_stmt_760_sources/type_cast_766/$exit
      -- CP-element group 275: 	 branch_block_stmt_34/forx_xbody150_forx_xbody150_PhiReq/phi_stmt_760/phi_stmt_760_sources/type_cast_766/SplitProtocol/$exit
      -- CP-element group 275: 	 branch_block_stmt_34/forx_xbody150_forx_xbody150_PhiReq/phi_stmt_760/phi_stmt_760_req
      -- 
    phi_stmt_760_req_2969_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_760_req_2969_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(275), ack => phi_stmt_760_req_1); -- 
    testConfigure_cp_element_group_275: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_275"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(273) & testConfigure_CP_0_elements(274);
      gj_testConfigure_cp_element_group_275 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(275), clk => clk, reset => reset); --
    end block;
    -- CP-element group 276:  merge  transition  place  bypass 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	272 
    -- CP-element group 276: 	275 
    -- CP-element group 276: successors 
    -- CP-element group 276: 	277 
    -- CP-element group 276:  members (2) 
      -- CP-element group 276: 	 branch_block_stmt_34/merge_stmt_759_PhiReqMerge
      -- CP-element group 276: 	 branch_block_stmt_34/merge_stmt_759_PhiAck/$entry
      -- 
    testConfigure_CP_0_elements(276) <= OrReduce(testConfigure_CP_0_elements(272) & testConfigure_CP_0_elements(275));
    -- CP-element group 277:  fork  transition  place  input  output  bypass 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	276 
    -- CP-element group 277: successors 
    -- CP-element group 277: 	171 
    -- CP-element group 277: 	172 
    -- CP-element group 277: 	174 
    -- CP-element group 277: 	175 
    -- CP-element group 277: 	178 
    -- CP-element group 277: 	182 
    -- CP-element group 277: 	186 
    -- CP-element group 277: 	190 
    -- CP-element group 277: 	194 
    -- CP-element group 277: 	198 
    -- CP-element group 277: 	202 
    -- CP-element group 277: 	206 
    -- CP-element group 277: 	209 
    -- CP-element group 277:  members (56) 
      -- CP-element group 277: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_901_Update/cr
      -- CP-element group 277: 	 branch_block_stmt_34/merge_stmt_759__exit__
      -- CP-element group 277: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922__entry__
      -- CP-element group 277: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_901_Update/$entry
      -- CP-element group 277: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_847_update_start_
      -- CP-element group 277: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_883_Update/$entry
      -- CP-element group 277: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_883_Update/cr
      -- CP-element group 277: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/ptr_deref_909_update_start_
      -- CP-element group 277: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_901_update_start_
      -- CP-element group 277: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_883_update_start_
      -- CP-element group 277: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_847_Update/cr
      -- CP-element group 277: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_847_Update/$entry
      -- CP-element group 277: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/ptr_deref_909_Update/word_access_complete/word_0/cr
      -- CP-element group 277: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/ptr_deref_909_Update/word_access_complete/word_0/$entry
      -- CP-element group 277: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/ptr_deref_909_Update/word_access_complete/$entry
      -- CP-element group 277: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/ptr_deref_909_Update/$entry
      -- CP-element group 277: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_865_Update/cr
      -- CP-element group 277: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_865_Update/$entry
      -- CP-element group 277: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_829_Update/cr
      -- CP-element group 277: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_865_update_start_
      -- CP-element group 277: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_829_Update/$entry
      -- CP-element group 277: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/$entry
      -- CP-element group 277: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/addr_of_773_update_start_
      -- CP-element group 277: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/array_obj_ref_772_index_resized_1
      -- CP-element group 277: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/array_obj_ref_772_index_scaled_1
      -- CP-element group 277: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/array_obj_ref_772_index_computed_1
      -- CP-element group 277: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/array_obj_ref_772_index_resize_1/$entry
      -- CP-element group 277: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/array_obj_ref_772_index_resize_1/$exit
      -- CP-element group 277: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/array_obj_ref_772_index_resize_1/index_resize_req
      -- CP-element group 277: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/array_obj_ref_772_index_resize_1/index_resize_ack
      -- CP-element group 277: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/array_obj_ref_772_index_scale_1/$entry
      -- CP-element group 277: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/array_obj_ref_772_index_scale_1/$exit
      -- CP-element group 277: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/array_obj_ref_772_index_scale_1/scale_rename_req
      -- CP-element group 277: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/array_obj_ref_772_index_scale_1/scale_rename_ack
      -- CP-element group 277: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/array_obj_ref_772_final_index_sum_regn_update_start
      -- CP-element group 277: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/array_obj_ref_772_final_index_sum_regn_Sample/$entry
      -- CP-element group 277: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/array_obj_ref_772_final_index_sum_regn_Sample/req
      -- CP-element group 277: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/array_obj_ref_772_final_index_sum_regn_Update/$entry
      -- CP-element group 277: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/array_obj_ref_772_final_index_sum_regn_Update/req
      -- CP-element group 277: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/addr_of_773_complete/$entry
      -- CP-element group 277: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/addr_of_773_complete/req
      -- CP-element group 277: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_776_sample_start_
      -- CP-element group 277: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_776_Sample/$entry
      -- CP-element group 277: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/RPIPE_ConvTranspose_input_pipe_776_Sample/rr
      -- CP-element group 277: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_780_update_start_
      -- CP-element group 277: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_780_Update/$entry
      -- CP-element group 277: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_780_Update/cr
      -- CP-element group 277: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_793_update_start_
      -- CP-element group 277: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_793_Update/$entry
      -- CP-element group 277: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_793_Update/cr
      -- CP-element group 277: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_811_update_start_
      -- CP-element group 277: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_811_Update/$entry
      -- CP-element group 277: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_811_Update/cr
      -- CP-element group 277: 	 branch_block_stmt_34/assign_stmt_774_to_assign_stmt_922/type_cast_829_update_start_
      -- CP-element group 277: 	 branch_block_stmt_34/merge_stmt_759_PhiAck/$exit
      -- CP-element group 277: 	 branch_block_stmt_34/merge_stmt_759_PhiAck/phi_stmt_760_ack
      -- 
    phi_stmt_760_ack_2974_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 277_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_760_ack_0, ack => testConfigure_CP_0_elements(277)); -- 
    cr_2231_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2231_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(277), ack => type_cast_901_inst_req_1); -- 
    cr_2203_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2203_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(277), ack => type_cast_883_inst_req_1); -- 
    cr_2147_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2147_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(277), ack => type_cast_847_inst_req_1); -- 
    cr_2281_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2281_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(277), ack => ptr_deref_909_store_0_req_1); -- 
    cr_2175_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2175_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(277), ack => type_cast_865_inst_req_1); -- 
    cr_2119_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2119_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(277), ack => type_cast_829_inst_req_1); -- 
    req_1987_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1987_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(277), ack => array_obj_ref_772_index_offset_req_0); -- 
    req_1992_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1992_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(277), ack => array_obj_ref_772_index_offset_req_1); -- 
    req_2007_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2007_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(277), ack => addr_of_773_final_reg_req_1); -- 
    rr_2016_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2016_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(277), ack => RPIPE_ConvTranspose_input_pipe_776_inst_req_0); -- 
    cr_2035_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2035_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(277), ack => type_cast_780_inst_req_1); -- 
    cr_2063_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2063_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(277), ack => type_cast_793_inst_req_1); -- 
    cr_2091_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2091_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(277), ack => type_cast_811_inst_req_1); -- 
    -- CP-element group 278:  merge  place  bypass 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	124 
    -- CP-element group 278: 	211 
    -- CP-element group 278: successors 
    -- CP-element group 278: 	279 
    -- CP-element group 278:  members (1) 
      -- CP-element group 278: 	 branch_block_stmt_34/merge_stmt_931_PhiReqMerge
      -- 
    testConfigure_CP_0_elements(278) <= OrReduce(testConfigure_CP_0_elements(124) & testConfigure_CP_0_elements(211));
    -- CP-element group 279:  join  fork  transition  place  output  bypass 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	278 
    -- CP-element group 279: successors 
    -- CP-element group 279: 	213 
    -- CP-element group 279: 	214 
    -- CP-element group 279: 	215 
    -- CP-element group 279: 	216 
    -- CP-element group 279: 	217 
    -- CP-element group 279: 	218 
    -- CP-element group 279:  members (84) 
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_942_base_addr_resize/$entry
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_942_base_address_calculated
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_942_word_address_calculated
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_942_root_address_calculated
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_942_base_plus_offset/sum_rename_req
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_954_Sample/word_access_start/word_0/$entry
      -- CP-element group 279: 	 branch_block_stmt_34/merge_stmt_931__exit__
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983__entry__
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_942_Sample/word_access_start/$entry
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_942_base_plus_offset/sum_rename_ack
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_942_word_addrgen/root_register_ack
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_966_word_addrgen/root_register_req
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_942_Sample/$entry
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_966_word_addrgen/root_register_ack
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_942_base_addr_resize/$exit
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_942_Sample/word_access_start/word_0/$entry
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_942_word_addrgen/$entry
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_942_base_address_resized
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_942_Sample/word_access_start/word_0/rr
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_942_Update/$entry
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_942_base_addr_resize/base_resize_ack
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_954_base_addr_resize/$exit
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_942_base_plus_offset/$exit
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_954_Update/$entry
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_966_Sample/$entry
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_942_base_addr_resize/base_resize_req
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_942_word_addrgen/root_register_req
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_954_Sample/word_access_start/word_0/rr
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_966_word_addrgen/$entry
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_966_word_addrgen/$exit
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_942_base_plus_offset/$entry
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_942_Update/word_access_complete/$entry
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_942_Update/word_access_complete/word_0/$entry
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_942_word_addrgen/$exit
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_942_Update/word_access_complete/word_0/cr
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_966_Sample/word_access_start/$entry
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_966_Sample/word_access_start/word_0/$entry
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_954_sample_start_
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_954_update_start_
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_966_Sample/word_access_start/word_0/rr
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_954_base_address_calculated
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_954_word_address_calculated
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_954_root_address_calculated
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_954_base_address_resized
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_954_Update/word_access_complete/$entry
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_954_base_addr_resize/$entry
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_942_update_start_
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_954_Sample/word_access_start/$entry
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_954_Sample/$entry
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_954_word_addrgen/root_register_ack
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_966_base_plus_offset/sum_rename_ack
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_966_base_plus_offset/sum_rename_req
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_954_word_addrgen/root_register_req
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_954_word_addrgen/$exit
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_954_word_addrgen/$entry
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_966_base_plus_offset/$exit
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_942_sample_start_
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_954_base_plus_offset/sum_rename_ack
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/$entry
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_954_base_plus_offset/sum_rename_req
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_966_base_plus_offset/$entry
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_966_base_addr_resize/base_resize_ack
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_966_base_addr_resize/base_resize_req
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_966_base_addr_resize/$exit
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_966_base_addr_resize/$entry
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_966_base_address_resized
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_966_root_address_calculated
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_966_word_address_calculated
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_966_base_address_calculated
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_966_update_start_
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_966_sample_start_
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_966_Update/word_access_complete/word_0/cr
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_966_Update/word_access_complete/word_0/$entry
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_966_Update/word_access_complete/$entry
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_966_Update/$entry
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_954_Update/word_access_complete/word_0/cr
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_954_base_plus_offset/$exit
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_954_base_plus_offset/$entry
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_954_Update/word_access_complete/word_0/$entry
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_954_base_addr_resize/base_resize_ack
      -- CP-element group 279: 	 branch_block_stmt_34/assign_stmt_939_to_assign_stmt_983/ptr_deref_954_base_addr_resize/base_resize_req
      -- CP-element group 279: 	 branch_block_stmt_34/merge_stmt_931_PhiAck/$entry
      -- CP-element group 279: 	 branch_block_stmt_34/merge_stmt_931_PhiAck/$exit
      -- CP-element group 279: 	 branch_block_stmt_34/merge_stmt_931_PhiAck/dummy
      -- 
    rr_2337_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2337_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(279), ack => ptr_deref_942_load_0_req_0); -- 
    rr_2387_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2387_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(279), ack => ptr_deref_954_load_0_req_0); -- 
    cr_2348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(279), ack => ptr_deref_942_load_0_req_1); -- 
    rr_2437_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2437_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(279), ack => ptr_deref_966_load_0_req_0); -- 
    cr_2448_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2448_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(279), ack => ptr_deref_966_load_0_req_1); -- 
    cr_2398_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2398_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(279), ack => ptr_deref_954_load_0_req_1); -- 
    testConfigure_CP_0_elements(279) <= testConfigure_CP_0_elements(278);
    -- CP-element group 280:  transition  output  delay-element  bypass 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	223 
    -- CP-element group 280: successors 
    -- CP-element group 280: 	284 
    -- CP-element group 280:  members (5) 
      -- CP-element group 280: 	 branch_block_stmt_34/bbx_xnph_forx_xbody217_PhiReq/$exit
      -- CP-element group 280: 	 branch_block_stmt_34/bbx_xnph_forx_xbody217_PhiReq/phi_stmt_1028/$exit
      -- CP-element group 280: 	 branch_block_stmt_34/bbx_xnph_forx_xbody217_PhiReq/phi_stmt_1028/phi_stmt_1028_sources/$exit
      -- CP-element group 280: 	 branch_block_stmt_34/bbx_xnph_forx_xbody217_PhiReq/phi_stmt_1028/phi_stmt_1028_sources/type_cast_1032_konst_delay_trans
      -- CP-element group 280: 	 branch_block_stmt_34/bbx_xnph_forx_xbody217_PhiReq/phi_stmt_1028/phi_stmt_1028_req
      -- 
    phi_stmt_1028_req_3020_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1028_req_3020_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(280), ack => phi_stmt_1028_req_0); -- 
    -- Element group testConfigure_CP_0_elements(280) is a control-delay.
    cp_element_280_delay: control_delay_element  generic map(name => " 280_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(223), ack => testConfigure_CP_0_elements(280), clk => clk, reset =>reset);
    -- CP-element group 281:  transition  input  bypass 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	232 
    -- CP-element group 281: successors 
    -- CP-element group 281: 	283 
    -- CP-element group 281:  members (2) 
      -- CP-element group 281: 	 branch_block_stmt_34/forx_xbody217_forx_xbody217_PhiReq/phi_stmt_1028/phi_stmt_1028_sources/type_cast_1034/SplitProtocol/Sample/$exit
      -- CP-element group 281: 	 branch_block_stmt_34/forx_xbody217_forx_xbody217_PhiReq/phi_stmt_1028/phi_stmt_1028_sources/type_cast_1034/SplitProtocol/Sample/ra
      -- 
    ra_3040_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 281_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1034_inst_ack_0, ack => testConfigure_CP_0_elements(281)); -- 
    -- CP-element group 282:  transition  input  bypass 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	232 
    -- CP-element group 282: successors 
    -- CP-element group 282: 	283 
    -- CP-element group 282:  members (2) 
      -- CP-element group 282: 	 branch_block_stmt_34/forx_xbody217_forx_xbody217_PhiReq/phi_stmt_1028/phi_stmt_1028_sources/type_cast_1034/SplitProtocol/Update/$exit
      -- CP-element group 282: 	 branch_block_stmt_34/forx_xbody217_forx_xbody217_PhiReq/phi_stmt_1028/phi_stmt_1028_sources/type_cast_1034/SplitProtocol/Update/ca
      -- 
    ca_3045_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 282_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1034_inst_ack_1, ack => testConfigure_CP_0_elements(282)); -- 
    -- CP-element group 283:  join  transition  output  bypass 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: 	281 
    -- CP-element group 283: 	282 
    -- CP-element group 283: successors 
    -- CP-element group 283: 	284 
    -- CP-element group 283:  members (6) 
      -- CP-element group 283: 	 branch_block_stmt_34/forx_xbody217_forx_xbody217_PhiReq/$exit
      -- CP-element group 283: 	 branch_block_stmt_34/forx_xbody217_forx_xbody217_PhiReq/phi_stmt_1028/$exit
      -- CP-element group 283: 	 branch_block_stmt_34/forx_xbody217_forx_xbody217_PhiReq/phi_stmt_1028/phi_stmt_1028_sources/$exit
      -- CP-element group 283: 	 branch_block_stmt_34/forx_xbody217_forx_xbody217_PhiReq/phi_stmt_1028/phi_stmt_1028_sources/type_cast_1034/$exit
      -- CP-element group 283: 	 branch_block_stmt_34/forx_xbody217_forx_xbody217_PhiReq/phi_stmt_1028/phi_stmt_1028_sources/type_cast_1034/SplitProtocol/$exit
      -- CP-element group 283: 	 branch_block_stmt_34/forx_xbody217_forx_xbody217_PhiReq/phi_stmt_1028/phi_stmt_1028_req
      -- 
    phi_stmt_1028_req_3046_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1028_req_3046_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(283), ack => phi_stmt_1028_req_1); -- 
    testConfigure_cp_element_group_283: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_283"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(281) & testConfigure_CP_0_elements(282);
      gj_testConfigure_cp_element_group_283 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(283), clk => clk, reset => reset); --
    end block;
    -- CP-element group 284:  merge  transition  place  bypass 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	280 
    -- CP-element group 284: 	283 
    -- CP-element group 284: successors 
    -- CP-element group 284: 	285 
    -- CP-element group 284:  members (2) 
      -- CP-element group 284: 	 branch_block_stmt_34/merge_stmt_1027_PhiReqMerge
      -- CP-element group 284: 	 branch_block_stmt_34/merge_stmt_1027_PhiAck/$entry
      -- 
    testConfigure_CP_0_elements(284) <= OrReduce(testConfigure_CP_0_elements(280) & testConfigure_CP_0_elements(283));
    -- CP-element group 285:  fork  transition  place  input  output  bypass 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: 	284 
    -- CP-element group 285: successors 
    -- CP-element group 285: 	224 
    -- CP-element group 285: 	225 
    -- CP-element group 285: 	227 
    -- CP-element group 285: 	229 
    -- CP-element group 285:  members (29) 
      -- CP-element group 285: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/array_obj_ref_1040_index_resized_1
      -- CP-element group 285: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/array_obj_ref_1040_final_index_sum_regn_Update/req
      -- CP-element group 285: 	 branch_block_stmt_34/merge_stmt_1027__exit__
      -- CP-element group 285: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058__entry__
      -- CP-element group 285: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/addr_of_1041_complete/$entry
      -- CP-element group 285: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/array_obj_ref_1040_index_scaled_1
      -- CP-element group 285: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/array_obj_ref_1040_index_computed_1
      -- CP-element group 285: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/array_obj_ref_1040_index_resize_1/$entry
      -- CP-element group 285: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/addr_of_1041_complete/req
      -- CP-element group 285: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/array_obj_ref_1040_final_index_sum_regn_Update/$entry
      -- CP-element group 285: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/array_obj_ref_1040_final_index_sum_regn_Sample/req
      -- CP-element group 285: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/addr_of_1041_update_start_
      -- CP-element group 285: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/array_obj_ref_1040_final_index_sum_regn_Sample/$entry
      -- CP-element group 285: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/array_obj_ref_1040_final_index_sum_regn_update_start
      -- CP-element group 285: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/ptr_deref_1044_update_start_
      -- CP-element group 285: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/$entry
      -- CP-element group 285: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/array_obj_ref_1040_index_scale_1/scale_rename_ack
      -- CP-element group 285: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/array_obj_ref_1040_index_scale_1/scale_rename_req
      -- CP-element group 285: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/array_obj_ref_1040_index_scale_1/$exit
      -- CP-element group 285: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/array_obj_ref_1040_index_scale_1/$entry
      -- CP-element group 285: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/array_obj_ref_1040_index_resize_1/index_resize_ack
      -- CP-element group 285: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/array_obj_ref_1040_index_resize_1/index_resize_req
      -- CP-element group 285: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/array_obj_ref_1040_index_resize_1/$exit
      -- CP-element group 285: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/ptr_deref_1044_Update/$entry
      -- CP-element group 285: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/ptr_deref_1044_Update/word_access_complete/$entry
      -- CP-element group 285: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/ptr_deref_1044_Update/word_access_complete/word_0/$entry
      -- CP-element group 285: 	 branch_block_stmt_34/assign_stmt_1042_to_assign_stmt_1058/ptr_deref_1044_Update/word_access_complete/word_0/cr
      -- CP-element group 285: 	 branch_block_stmt_34/merge_stmt_1027_PhiAck/$exit
      -- CP-element group 285: 	 branch_block_stmt_34/merge_stmt_1027_PhiAck/phi_stmt_1028_ack
      -- 
    phi_stmt_1028_ack_3051_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 285_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1028_ack_0, ack => testConfigure_CP_0_elements(285)); -- 
    req_2523_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2523_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(285), ack => array_obj_ref_1040_index_offset_req_1); -- 
    req_2538_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2538_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(285), ack => addr_of_1041_final_reg_req_1); -- 
    req_2518_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2518_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(285), ack => array_obj_ref_1040_index_offset_req_0); -- 
    cr_2588_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2588_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(285), ack => ptr_deref_1044_store_0_req_1); -- 
    -- CP-element group 286:  merge  transition  place  bypass 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	221 
    -- CP-element group 286: 	231 
    -- CP-element group 286: successors 
    -- CP-element group 286:  members (20) 
      -- CP-element group 286: 	 $exit
      -- CP-element group 286: 	 branch_block_stmt_34/$exit
      -- CP-element group 286: 	 branch_block_stmt_34/branch_block_stmt_34__exit__
      -- CP-element group 286: 	 branch_block_stmt_34/merge_stmt_1067__exit__
      -- CP-element group 286: 	 branch_block_stmt_34/assign_stmt_1071__entry__
      -- CP-element group 286: 	 branch_block_stmt_34/assign_stmt_1071__exit__
      -- CP-element group 286: 	 branch_block_stmt_34/return__
      -- CP-element group 286: 	 branch_block_stmt_34/merge_stmt_1073__exit__
      -- CP-element group 286: 	 branch_block_stmt_34/assign_stmt_1071/$entry
      -- CP-element group 286: 	 branch_block_stmt_34/assign_stmt_1071/$exit
      -- CP-element group 286: 	 branch_block_stmt_34/merge_stmt_1067_PhiReqMerge
      -- CP-element group 286: 	 branch_block_stmt_34/merge_stmt_1067_PhiAck/$entry
      -- CP-element group 286: 	 branch_block_stmt_34/merge_stmt_1067_PhiAck/$exit
      -- CP-element group 286: 	 branch_block_stmt_34/merge_stmt_1067_PhiAck/dummy
      -- CP-element group 286: 	 branch_block_stmt_34/return___PhiReq/$entry
      -- CP-element group 286: 	 branch_block_stmt_34/return___PhiReq/$exit
      -- CP-element group 286: 	 branch_block_stmt_34/merge_stmt_1073_PhiReqMerge
      -- CP-element group 286: 	 branch_block_stmt_34/merge_stmt_1073_PhiAck/$entry
      -- CP-element group 286: 	 branch_block_stmt_34/merge_stmt_1073_PhiAck/$exit
      -- CP-element group 286: 	 branch_block_stmt_34/merge_stmt_1073_PhiAck/dummy
      -- 
    testConfigure_CP_0_elements(286) <= OrReduce(testConfigure_CP_0_elements(221) & testConfigure_CP_0_elements(231));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_indvar253_771_resized : std_logic_vector(10 downto 0);
    signal R_indvar253_771_scaled : std_logic_vector(10 downto 0);
    signal R_indvar265_564_resized : std_logic_vector(13 downto 0);
    signal R_indvar265_564_scaled : std_logic_vector(13 downto 0);
    signal R_indvar277_194_resized : std_logic_vector(0 downto 0);
    signal R_indvar277_194_scaled : std_logic_vector(0 downto 0);
    signal R_indvar280_118_resized : std_logic_vector(6 downto 0);
    signal R_indvar280_118_scaled : std_logic_vector(6 downto 0);
    signal R_indvar283_48_resized : std_logic_vector(6 downto 0);
    signal R_indvar283_48_scaled : std_logic_vector(6 downto 0);
    signal R_indvar_1039_resized : std_logic_vector(13 downto 0);
    signal R_indvar_1039_scaled : std_logic_vector(13 downto 0);
    signal STORE_padding_229_data_0 : std_logic_vector(7 downto 0);
    signal STORE_padding_229_word_address_0 : std_logic_vector(0 downto 0);
    signal add105_610 : std_logic_vector(63 downto 0);
    signal add111_628 : std_logic_vector(63 downto 0);
    signal add117_646 : std_logic_vector(63 downto 0);
    signal add123_664 : std_logic_vector(63 downto 0);
    signal add129_682 : std_logic_vector(63 downto 0);
    signal add135_700 : std_logic_vector(63 downto 0);
    signal add160_799 : std_logic_vector(63 downto 0);
    signal add166_817 : std_logic_vector(63 downto 0);
    signal add172_835 : std_logic_vector(63 downto 0);
    signal add178_853 : std_logic_vector(63 downto 0);
    signal add184_871 : std_logic_vector(63 downto 0);
    signal add190_889 : std_logic_vector(63 downto 0);
    signal add196_907 : std_logic_vector(63 downto 0);
    signal add29_150 : std_logic_vector(31 downto 0);
    signal add57_268 : std_logic_vector(31 downto 0);
    signal add64_317 : std_logic_vector(31 downto 0);
    signal add71_366 : std_logic_vector(31 downto 0);
    signal add99_592 : std_logic_vector(63 downto 0);
    signal add_80 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1040_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1040_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1040_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1040_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1040_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1040_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_119_constant_part_of_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_119_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_119_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_119_offset_scale_factor_1 : std_logic_vector(6 downto 0);
    signal array_obj_ref_119_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_119_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_195_final_offset : std_logic_vector(0 downto 0);
    signal array_obj_ref_195_offset_scale_factor_0 : std_logic_vector(0 downto 0);
    signal array_obj_ref_195_resized_base_address : std_logic_vector(0 downto 0);
    signal array_obj_ref_195_root_address : std_logic_vector(0 downto 0);
    signal array_obj_ref_49_constant_part_of_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_49_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_49_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_49_offset_scale_factor_1 : std_logic_vector(6 downto 0);
    signal array_obj_ref_49_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_49_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_565_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_565_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_565_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_565_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_565_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_565_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_772_constant_part_of_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_772_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_772_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_772_offset_scale_factor_1 : std_logic_vector(10 downto 0);
    signal array_obj_ref_772_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_772_root_address : std_logic_vector(10 downto 0);
    signal arrayidx10_51 : std_logic_vector(31 downto 0);
    signal arrayidx139_567 : std_logic_vector(31 downto 0);
    signal arrayidx200_774 : std_logic_vector(31 downto 0);
    signal arrayidx220_1042 : std_logic_vector(31 downto 0);
    signal arrayidx32_121 : std_logic_vector(31 downto 0);
    signal arrayidx45_197 : std_logic_vector(31 downto 0);
    signal call102_601 : std_logic_vector(7 downto 0);
    signal call108_619 : std_logic_vector(7 downto 0);
    signal call114_637 : std_logic_vector(7 downto 0);
    signal call120_655 : std_logic_vector(7 downto 0);
    signal call126_673 : std_logic_vector(7 downto 0);
    signal call132_691 : std_logic_vector(7 downto 0);
    signal call153_777 : std_logic_vector(7 downto 0);
    signal call157_790 : std_logic_vector(7 downto 0);
    signal call163_808 : std_logic_vector(7 downto 0);
    signal call169_826 : std_logic_vector(7 downto 0);
    signal call175_844 : std_logic_vector(7 downto 0);
    signal call17_124 : std_logic_vector(7 downto 0);
    signal call181_862 : std_logic_vector(7 downto 0);
    signal call187_880 : std_logic_vector(7 downto 0);
    signal call193_898 : std_logic_vector(7 downto 0);
    signal call27_141 : std_logic_vector(7 downto 0);
    signal call42237_176 : std_logic_vector(7 downto 0);
    signal call42239_186 : std_logic_vector(7 downto 0);
    signal call42_204 : std_logic_vector(7 downto 0);
    signal call42x_xlcssa_224 : std_logic_vector(7 downto 0);
    signal call51_234 : std_logic_vector(7 downto 0);
    signal call55_259 : std_logic_vector(7 downto 0);
    signal call58_283 : std_logic_vector(7 downto 0);
    signal call62_308 : std_logic_vector(7 downto 0);
    signal call65_332 : std_logic_vector(7 downto 0);
    signal call69_357 : std_logic_vector(7 downto 0);
    signal call6_71 : std_logic_vector(7 downto 0);
    signal call92_570 : std_logic_vector(7 downto 0);
    signal call96_583 : std_logic_vector(7 downto 0);
    signal call_54 : std_logic_vector(7 downto 0);
    signal cmp148229_508 : std_logic_vector(0 downto 0);
    signal cmp215226_983 : std_logic_vector(0 downto 0);
    signal cmp88233_493 : std_logic_vector(0 downto 0);
    signal conv104_605 : std_logic_vector(63 downto 0);
    signal conv110_623 : std_logic_vector(63 downto 0);
    signal conv116_641 : std_logic_vector(63 downto 0);
    signal conv122_659 : std_logic_vector(63 downto 0);
    signal conv128_677 : std_logic_vector(63 downto 0);
    signal conv134_695 : std_logic_vector(63 downto 0);
    signal conv154_781 : std_logic_vector(63 downto 0);
    signal conv159_794 : std_logic_vector(63 downto 0);
    signal conv165_812 : std_logic_vector(63 downto 0);
    signal conv171_830 : std_logic_vector(63 downto 0);
    signal conv177_848 : std_logic_vector(63 downto 0);
    signal conv183_866 : std_logic_vector(63 downto 0);
    signal conv189_884 : std_logic_vector(63 downto 0);
    signal conv18_128 : std_logic_vector(31 downto 0);
    signal conv195_902 : std_logic_vector(63 downto 0);
    signal conv28_145 : std_logic_vector(31 downto 0);
    signal conv52_238 : std_logic_vector(31 downto 0);
    signal conv56_263 : std_logic_vector(31 downto 0);
    signal conv59_287 : std_logic_vector(31 downto 0);
    signal conv63_312 : std_logic_vector(31 downto 0);
    signal conv66_336 : std_logic_vector(31 downto 0);
    signal conv70_361 : std_logic_vector(31 downto 0);
    signal conv7_75 : std_logic_vector(31 downto 0);
    signal conv93_574 : std_logic_vector(63 downto 0);
    signal conv98_587 : std_logic_vector(63 downto 0);
    signal conv_58 : std_logic_vector(31 downto 0);
    signal exitcond1_1058 : std_logic_vector(0 downto 0);
    signal exitcond2_715 : std_logic_vector(0 downto 0);
    signal exitcond3_216 : std_logic_vector(0 downto 0);
    signal exitcond4_166 : std_logic_vector(0 downto 0);
    signal exitcond5_97 : std_logic_vector(0 downto 0);
    signal exitcond_922 : std_logic_vector(0 downto 0);
    signal iNsTr_19_246 : std_logic_vector(31 downto 0);
    signal iNsTr_22_276 : std_logic_vector(31 downto 0);
    signal iNsTr_25_295 : std_logic_vector(31 downto 0);
    signal iNsTr_28_325 : std_logic_vector(31 downto 0);
    signal iNsTr_31_344 : std_logic_vector(31 downto 0);
    signal iNsTr_34_374 : std_logic_vector(31 downto 0);
    signal iNsTr_36_386 : std_logic_vector(31 downto 0);
    signal iNsTr_37_398 : std_logic_vector(31 downto 0);
    signal iNsTr_38_410 : std_logic_vector(31 downto 0);
    signal iNsTr_39_432 : std_logic_vector(31 downto 0);
    signal iNsTr_40_444 : std_logic_vector(31 downto 0);
    signal iNsTr_41_456 : std_logic_vector(31 downto 0);
    signal iNsTr_42_468 : std_logic_vector(31 downto 0);
    signal iNsTr_44_537 : std_logic_vector(63 downto 0);
    signal iNsTr_57_744 : std_logic_vector(63 downto 0);
    signal iNsTr_59_939 : std_logic_vector(31 downto 0);
    signal iNsTr_60_951 : std_logic_vector(31 downto 0);
    signal iNsTr_61_963 : std_logic_vector(31 downto 0);
    signal iNsTr_74_1012 : std_logic_vector(63 downto 0);
    signal indvar253_760 : std_logic_vector(63 downto 0);
    signal indvar265_553 : std_logic_vector(63 downto 0);
    signal indvar277_179 : std_logic_vector(63 downto 0);
    signal indvar280_107 : std_logic_vector(63 downto 0);
    signal indvar283_37 : std_logic_vector(63 downto 0);
    signal indvar_1028 : std_logic_vector(63 downto 0);
    signal indvarx_xnext254_917 : std_logic_vector(63 downto 0);
    signal indvarx_xnext266_710 : std_logic_vector(63 downto 0);
    signal indvarx_xnext278_210 : std_logic_vector(63 downto 0);
    signal indvarx_xnext281_160 : std_logic_vector(63 downto 0);
    signal indvarx_xnext284_90 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_1053 : std_logic_vector(63 downto 0);
    signal mul208_972 : std_logic_vector(31 downto 0);
    signal mul210_977 : std_logic_vector(31 downto 0);
    signal mul76_424 : std_logic_vector(31 downto 0);
    signal mul80_477 : std_logic_vector(31 downto 0);
    signal mul82_482 : std_logic_vector(31 downto 0);
    signal mul84_487 : std_logic_vector(31 downto 0);
    signal mul_419 : std_logic_vector(31 downto 0);
    signal ptr_deref_1044_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1044_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1044_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1044_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1044_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1044_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_130_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_130_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_130_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_130_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_130_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_130_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_152_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_152_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_152_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_152_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_152_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_152_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_199_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_199_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_199_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_199_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_199_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_199_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_248_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_248_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_248_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_248_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_248_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_248_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_278_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_278_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_278_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_278_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_278_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_278_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_297_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_297_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_297_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_297_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_297_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_297_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_327_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_327_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_327_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_327_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_327_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_327_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_346_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_346_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_346_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_346_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_346_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_346_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_376_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_376_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_376_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_376_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_376_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_376_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_389_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_389_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_389_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_389_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_389_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_401_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_401_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_401_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_401_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_401_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_413_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_413_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_413_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_413_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_413_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_435_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_435_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_435_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_435_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_435_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_447_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_447_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_447_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_447_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_447_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_459_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_459_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_459_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_459_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_459_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_471_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_471_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_471_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_471_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_471_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_60_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_60_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_60_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_60_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_60_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_60_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_702_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_702_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_702_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_702_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_702_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_702_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_82_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_82_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_82_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_82_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_82_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_82_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_909_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_909_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_909_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_909_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_909_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_909_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_942_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_942_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_942_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_942_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_942_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_954_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_954_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_954_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_954_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_954_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_966_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_966_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_966_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_966_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_966_word_offset_0 : std_logic_vector(6 downto 0);
    signal shl101_598 : std_logic_vector(63 downto 0);
    signal shl107_616 : std_logic_vector(63 downto 0);
    signal shl113_634 : std_logic_vector(63 downto 0);
    signal shl119_652 : std_logic_vector(63 downto 0);
    signal shl125_670 : std_logic_vector(63 downto 0);
    signal shl131_688 : std_logic_vector(63 downto 0);
    signal shl156_787 : std_logic_vector(63 downto 0);
    signal shl162_805 : std_logic_vector(63 downto 0);
    signal shl168_823 : std_logic_vector(63 downto 0);
    signal shl174_841 : std_logic_vector(63 downto 0);
    signal shl180_859 : std_logic_vector(63 downto 0);
    signal shl186_877 : std_logic_vector(63 downto 0);
    signal shl192_895 : std_logic_vector(63 downto 0);
    signal shl26_138 : std_logic_vector(31 downto 0);
    signal shl54_256 : std_logic_vector(31 downto 0);
    signal shl61_305 : std_logic_vector(31 downto 0);
    signal shl68_354 : std_logic_vector(31 downto 0);
    signal shl95_580 : std_logic_vector(63 downto 0);
    signal shl_68 : std_logic_vector(31 downto 0);
    signal tmp206_943 : std_logic_vector(31 downto 0);
    signal tmp207_955 : std_logic_vector(31 downto 0);
    signal tmp209_967 : std_logic_vector(31 downto 0);
    signal tmp248_996 : std_logic_vector(31 downto 0);
    signal tmp248x_xop_1008 : std_logic_vector(31 downto 0);
    signal tmp249_1002 : std_logic_vector(0 downto 0);
    signal tmp252_1025 : std_logic_vector(63 downto 0);
    signal tmp258_728 : std_logic_vector(31 downto 0);
    signal tmp258x_xop_740 : std_logic_vector(31 downto 0);
    signal tmp259_734 : std_logic_vector(0 downto 0);
    signal tmp263_757 : std_logic_vector(63 downto 0);
    signal tmp269_521 : std_logic_vector(31 downto 0);
    signal tmp269x_xop_533 : std_logic_vector(31 downto 0);
    signal tmp270_527 : std_logic_vector(0 downto 0);
    signal tmp274_550 : std_logic_vector(63 downto 0);
    signal tmp73_390 : std_logic_vector(31 downto 0);
    signal tmp74_402 : std_logic_vector(31 downto 0);
    signal tmp75_414 : std_logic_vector(31 downto 0);
    signal tmp78_436 : std_logic_vector(31 downto 0);
    signal tmp79_448 : std_logic_vector(31 downto 0);
    signal tmp81_460 : std_logic_vector(31 downto 0);
    signal tmp83_472 : std_logic_vector(31 downto 0);
    signal type_cast_1000_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1006_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1016_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1023_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1032_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1034_wire : std_logic_vector(63 downto 0);
    signal type_cast_1046_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1051_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_110_wire : std_logic_vector(63 downto 0);
    signal type_cast_113_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_136_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_158_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_164_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_183_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_185_wire : std_logic_vector(63 downto 0);
    signal type_cast_189_wire : std_logic_vector(7 downto 0);
    signal type_cast_191_wire : std_logic_vector(7 downto 0);
    signal type_cast_208_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_214_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_227_wire : std_logic_vector(7 downto 0);
    signal type_cast_254_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_303_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_352_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_41_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_43_wire : std_logic_vector(63 downto 0);
    signal type_cast_491_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_506_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_519_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_525_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_531_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_541_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_548_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_557_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_559_wire : std_logic_vector(63 downto 0);
    signal type_cast_578_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_596_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_614_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_632_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_650_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_668_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_66_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_686_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_708_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_726_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_732_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_738_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_748_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_755_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_764_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_766_wire : std_logic_vector(63 downto 0);
    signal type_cast_785_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_803_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_821_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_839_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_857_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_875_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_88_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_893_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_915_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_94_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_981_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_994_wire_constant : std_logic_vector(31 downto 0);
    signal xx_xop286_750 : std_logic_vector(63 downto 0);
    signal xx_xop287_543 : std_logic_vector(63 downto 0);
    signal xx_xop_1018 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    STORE_padding_229_word_address_0 <= "0";
    array_obj_ref_1040_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1040_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1040_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1040_resized_base_address <= "00000000000000";
    array_obj_ref_119_constant_part_of_offset <= "0000011";
    array_obj_ref_119_offset_scale_factor_0 <= "1000000";
    array_obj_ref_119_offset_scale_factor_1 <= "0000001";
    array_obj_ref_119_resized_base_address <= "0000000";
    array_obj_ref_195_offset_scale_factor_0 <= "1";
    array_obj_ref_195_resized_base_address <= "0";
    array_obj_ref_49_constant_part_of_offset <= "0000011";
    array_obj_ref_49_offset_scale_factor_0 <= "1000000";
    array_obj_ref_49_offset_scale_factor_1 <= "0000001";
    array_obj_ref_49_resized_base_address <= "0000000";
    array_obj_ref_565_constant_part_of_offset <= "00000000000000";
    array_obj_ref_565_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_565_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_565_resized_base_address <= "00000000000000";
    array_obj_ref_772_constant_part_of_offset <= "00000100010";
    array_obj_ref_772_offset_scale_factor_0 <= "10000000000";
    array_obj_ref_772_offset_scale_factor_1 <= "00000000001";
    array_obj_ref_772_resized_base_address <= "00000000000";
    iNsTr_19_246 <= "00000000000000000000000000000011";
    iNsTr_22_276 <= "00000000000000000000000000000011";
    iNsTr_25_295 <= "00000000000000000000000000000100";
    iNsTr_28_325 <= "00000000000000000000000000000100";
    iNsTr_31_344 <= "00000000000000000000000000000101";
    iNsTr_34_374 <= "00000000000000000000000000000101";
    iNsTr_36_386 <= "00000000000000000000000000000011";
    iNsTr_37_398 <= "00000000000000000000000000000100";
    iNsTr_38_410 <= "00000000000000000000000000000101";
    iNsTr_39_432 <= "00000000000000000000000000000011";
    iNsTr_40_444 <= "00000000000000000000000000000100";
    iNsTr_41_456 <= "00000000000000000000000000000101";
    iNsTr_42_468 <= "00000000000000000000000000000110";
    iNsTr_59_939 <= "00000000000000000000000000000011";
    iNsTr_60_951 <= "00000000000000000000000000000100";
    iNsTr_61_963 <= "00000000000000000000000000000101";
    ptr_deref_1044_word_offset_0 <= "00000000000000";
    ptr_deref_130_word_offset_0 <= "0000000";
    ptr_deref_152_word_offset_0 <= "0000000";
    ptr_deref_199_word_offset_0 <= "0";
    ptr_deref_248_word_offset_0 <= "0000000";
    ptr_deref_278_word_offset_0 <= "0000000";
    ptr_deref_297_word_offset_0 <= "0000000";
    ptr_deref_327_word_offset_0 <= "0000000";
    ptr_deref_346_word_offset_0 <= "0000000";
    ptr_deref_376_word_offset_0 <= "0000000";
    ptr_deref_389_word_offset_0 <= "0000000";
    ptr_deref_401_word_offset_0 <= "0000000";
    ptr_deref_413_word_offset_0 <= "0000000";
    ptr_deref_435_word_offset_0 <= "0000000";
    ptr_deref_447_word_offset_0 <= "0000000";
    ptr_deref_459_word_offset_0 <= "0000000";
    ptr_deref_471_word_offset_0 <= "0000000";
    ptr_deref_60_word_offset_0 <= "0000000";
    ptr_deref_702_word_offset_0 <= "00000000000000";
    ptr_deref_82_word_offset_0 <= "0000000";
    ptr_deref_909_word_offset_0 <= "00000000000";
    ptr_deref_942_word_offset_0 <= "0000000";
    ptr_deref_954_word_offset_0 <= "0000000";
    ptr_deref_966_word_offset_0 <= "0000000";
    type_cast_1000_wire_constant <= "00000000000000000000000000000001";
    type_cast_1006_wire_constant <= "11111111111111111111111111111111";
    type_cast_1016_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1023_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1032_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1046_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1051_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_113_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_136_wire_constant <= "00000000000000000000000000001000";
    type_cast_158_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_164_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000100";
    type_cast_183_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_208_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_214_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_254_wire_constant <= "00000000000000000000000000001000";
    type_cast_303_wire_constant <= "00000000000000000000000000001000";
    type_cast_352_wire_constant <= "00000000000000000000000000001000";
    type_cast_41_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_491_wire_constant <= "00000000000000000000000000000111";
    type_cast_506_wire_constant <= "00000000000000000000000000000111";
    type_cast_519_wire_constant <= "00000000000000000000000000000011";
    type_cast_525_wire_constant <= "00000000000000000000000000000001";
    type_cast_531_wire_constant <= "11111111111111111111111111111111";
    type_cast_541_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_548_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_557_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_578_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_596_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_614_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_632_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_650_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_668_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_66_wire_constant <= "00000000000000000000000000001000";
    type_cast_686_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_708_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_726_wire_constant <= "00000000000000000000000000000011";
    type_cast_732_wire_constant <= "00000000000000000000000000000001";
    type_cast_738_wire_constant <= "11111111111111111111111111111111";
    type_cast_748_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_755_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_764_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_785_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_803_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_821_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_839_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_857_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_875_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_88_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_893_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_915_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_94_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    type_cast_981_wire_constant <= "00000000000000000000000000000011";
    type_cast_994_wire_constant <= "00000000000000000000000000000010";
    phi_stmt_1028: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1032_wire_constant & type_cast_1034_wire;
      req <= phi_stmt_1028_req_0 & phi_stmt_1028_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1028",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1028_ack_0,
          idata => idata,
          odata => indvar_1028,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1028
    phi_stmt_107: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_110_wire & type_cast_113_wire_constant;
      req <= phi_stmt_107_req_0 & phi_stmt_107_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_107",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_107_ack_0,
          idata => idata,
          odata => indvar280_107,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_107
    phi_stmt_179: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_183_wire_constant & type_cast_185_wire;
      req <= phi_stmt_179_req_0 & phi_stmt_179_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_179",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_179_ack_0,
          idata => idata,
          odata => indvar277_179,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_179
    phi_stmt_186: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_189_wire & type_cast_191_wire;
      req <= phi_stmt_186_req_0 & phi_stmt_186_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_186",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_186_ack_0,
          idata => idata,
          odata => call42239_186,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_186
    phi_stmt_224: Block -- phi operator 
      signal idata: std_logic_vector(7 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_227_wire;
      req(0) <= phi_stmt_224_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_224",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_224_ack_0,
          idata => idata,
          odata => call42x_xlcssa_224,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_224
    phi_stmt_37: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_41_wire_constant & type_cast_43_wire;
      req <= phi_stmt_37_req_0 & phi_stmt_37_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_37",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_37_ack_0,
          idata => idata,
          odata => indvar283_37,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_37
    phi_stmt_553: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_557_wire_constant & type_cast_559_wire;
      req <= phi_stmt_553_req_0 & phi_stmt_553_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_553",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_553_ack_0,
          idata => idata,
          odata => indvar265_553,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_553
    phi_stmt_760: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_764_wire_constant & type_cast_766_wire;
      req <= phi_stmt_760_req_0 & phi_stmt_760_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_760",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_760_ack_0,
          idata => idata,
          odata => indvar253_760,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_760
    -- flow-through select operator MUX_1024_inst
    tmp252_1025 <= xx_xop_1018 when (tmp249_1002(0) /=  '0') else type_cast_1023_wire_constant;
    -- flow-through select operator MUX_549_inst
    tmp274_550 <= xx_xop287_543 when (tmp270_527(0) /=  '0') else type_cast_548_wire_constant;
    -- flow-through select operator MUX_756_inst
    tmp263_757 <= xx_xop286_750 when (tmp259_734(0) /=  '0') else type_cast_755_wire_constant;
    addr_of_1041_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1041_final_reg_req_0;
      addr_of_1041_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1041_final_reg_req_1;
      addr_of_1041_final_reg_ack_1<= rack(0);
      addr_of_1041_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1041_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1040_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx220_1042,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_120_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_120_final_reg_req_0;
      addr_of_120_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_120_final_reg_req_1;
      addr_of_120_final_reg_ack_1<= rack(0);
      addr_of_120_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_120_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 7,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_119_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx32_121,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_196_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_196_final_reg_req_0;
      addr_of_196_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_196_final_reg_req_1;
      addr_of_196_final_reg_ack_1<= rack(0);
      addr_of_196_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_196_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_195_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx45_197,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_50_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_50_final_reg_req_0;
      addr_of_50_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_50_final_reg_req_1;
      addr_of_50_final_reg_ack_1<= rack(0);
      addr_of_50_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_50_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 7,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_49_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx10_51,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_566_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_566_final_reg_req_0;
      addr_of_566_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_566_final_reg_req_1;
      addr_of_566_final_reg_ack_1<= rack(0);
      addr_of_566_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_566_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_565_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx139_567,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_773_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_773_final_reg_req_0;
      addr_of_773_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_773_final_reg_req_1;
      addr_of_773_final_reg_ack_1<= rack(0);
      addr_of_773_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_773_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 11,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_772_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx200_774,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1011_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1011_inst_req_0;
      type_cast_1011_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1011_inst_req_1;
      type_cast_1011_inst_ack_1<= rack(0);
      type_cast_1011_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1011_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp248x_xop_1008,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_74_1012,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1034_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1034_inst_req_0;
      type_cast_1034_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1034_inst_req_1;
      type_cast_1034_inst_ack_1<= rack(0);
      type_cast_1034_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1034_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1053,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1034_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_110_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_110_inst_req_0;
      type_cast_110_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_110_inst_req_1;
      type_cast_110_inst_ack_1<= rack(0);
      type_cast_110_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_110_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext281_160,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_110_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_127_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_127_inst_req_0;
      type_cast_127_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_127_inst_req_1;
      type_cast_127_inst_ack_1<= rack(0);
      type_cast_127_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_127_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call17_124,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv18_128,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_144_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_144_inst_req_0;
      type_cast_144_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_144_inst_req_1;
      type_cast_144_inst_ack_1<= rack(0);
      type_cast_144_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_144_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call27_141,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv28_145,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_185_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_185_inst_req_0;
      type_cast_185_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_185_inst_req_1;
      type_cast_185_inst_ack_1<= rack(0);
      type_cast_185_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_185_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext278_210,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_185_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_189_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_189_inst_req_0;
      type_cast_189_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_189_inst_req_1;
      type_cast_189_inst_ack_1<= rack(0);
      type_cast_189_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_189_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call42237_176,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_189_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_191_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_191_inst_req_0;
      type_cast_191_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_191_inst_req_1;
      type_cast_191_inst_ack_1<= rack(0);
      type_cast_191_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_191_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call42_204,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_191_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_227_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_227_inst_req_0;
      type_cast_227_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_227_inst_req_1;
      type_cast_227_inst_ack_1<= rack(0);
      type_cast_227_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_227_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call42_204,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_227_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_237_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_237_inst_req_0;
      type_cast_237_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_237_inst_req_1;
      type_cast_237_inst_ack_1<= rack(0);
      type_cast_237_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_237_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call51_234,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv52_238,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_262_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_262_inst_req_0;
      type_cast_262_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_262_inst_req_1;
      type_cast_262_inst_ack_1<= rack(0);
      type_cast_262_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_262_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call55_259,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv56_263,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_286_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_286_inst_req_0;
      type_cast_286_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_286_inst_req_1;
      type_cast_286_inst_ack_1<= rack(0);
      type_cast_286_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_286_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call58_283,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv59_287,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_311_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_311_inst_req_0;
      type_cast_311_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_311_inst_req_1;
      type_cast_311_inst_ack_1<= rack(0);
      type_cast_311_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_311_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call62_308,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv63_312,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_335_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_335_inst_req_0;
      type_cast_335_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_335_inst_req_1;
      type_cast_335_inst_ack_1<= rack(0);
      type_cast_335_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_335_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call65_332,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv66_336,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_360_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_360_inst_req_0;
      type_cast_360_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_360_inst_req_1;
      type_cast_360_inst_ack_1<= rack(0);
      type_cast_360_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_360_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call69_357,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv70_361,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_43_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_43_inst_req_0;
      type_cast_43_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_43_inst_req_1;
      type_cast_43_inst_ack_1<= rack(0);
      type_cast_43_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_43_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext284_90,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_43_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_536_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_536_inst_req_0;
      type_cast_536_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_536_inst_req_1;
      type_cast_536_inst_ack_1<= rack(0);
      type_cast_536_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_536_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp269x_xop_533,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_44_537,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_559_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_559_inst_req_0;
      type_cast_559_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_559_inst_req_1;
      type_cast_559_inst_ack_1<= rack(0);
      type_cast_559_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_559_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext266_710,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_559_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_573_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_573_inst_req_0;
      type_cast_573_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_573_inst_req_1;
      type_cast_573_inst_ack_1<= rack(0);
      type_cast_573_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_573_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call92_570,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv93_574,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_57_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_57_inst_req_0;
      type_cast_57_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_57_inst_req_1;
      type_cast_57_inst_ack_1<= rack(0);
      type_cast_57_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_57_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_54,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_58,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_586_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_586_inst_req_0;
      type_cast_586_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_586_inst_req_1;
      type_cast_586_inst_ack_1<= rack(0);
      type_cast_586_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_586_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call96_583,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv98_587,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_604_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_604_inst_req_0;
      type_cast_604_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_604_inst_req_1;
      type_cast_604_inst_ack_1<= rack(0);
      type_cast_604_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_604_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call102_601,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv104_605,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_622_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_622_inst_req_0;
      type_cast_622_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_622_inst_req_1;
      type_cast_622_inst_ack_1<= rack(0);
      type_cast_622_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_622_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call108_619,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv110_623,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_640_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_640_inst_req_0;
      type_cast_640_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_640_inst_req_1;
      type_cast_640_inst_ack_1<= rack(0);
      type_cast_640_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_640_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call114_637,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv116_641,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_658_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_658_inst_req_0;
      type_cast_658_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_658_inst_req_1;
      type_cast_658_inst_ack_1<= rack(0);
      type_cast_658_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_658_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call120_655,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv122_659,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_676_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_676_inst_req_0;
      type_cast_676_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_676_inst_req_1;
      type_cast_676_inst_ack_1<= rack(0);
      type_cast_676_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_676_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call126_673,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv128_677,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_694_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_694_inst_req_0;
      type_cast_694_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_694_inst_req_1;
      type_cast_694_inst_ack_1<= rack(0);
      type_cast_694_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_694_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call132_691,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv134_695,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_743_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_743_inst_req_0;
      type_cast_743_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_743_inst_req_1;
      type_cast_743_inst_ack_1<= rack(0);
      type_cast_743_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_743_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp258x_xop_740,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_57_744,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_74_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_74_inst_req_0;
      type_cast_74_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_74_inst_req_1;
      type_cast_74_inst_ack_1<= rack(0);
      type_cast_74_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_74_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call6_71,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv7_75,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_766_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_766_inst_req_0;
      type_cast_766_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_766_inst_req_1;
      type_cast_766_inst_ack_1<= rack(0);
      type_cast_766_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_766_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext254_917,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_766_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_780_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_780_inst_req_0;
      type_cast_780_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_780_inst_req_1;
      type_cast_780_inst_ack_1<= rack(0);
      type_cast_780_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_780_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call153_777,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv154_781,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_793_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_793_inst_req_0;
      type_cast_793_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_793_inst_req_1;
      type_cast_793_inst_ack_1<= rack(0);
      type_cast_793_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_793_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call157_790,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv159_794,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_811_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_811_inst_req_0;
      type_cast_811_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_811_inst_req_1;
      type_cast_811_inst_ack_1<= rack(0);
      type_cast_811_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_811_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call163_808,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv165_812,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_829_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_829_inst_req_0;
      type_cast_829_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_829_inst_req_1;
      type_cast_829_inst_ack_1<= rack(0);
      type_cast_829_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_829_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call169_826,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv171_830,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_847_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_847_inst_req_0;
      type_cast_847_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_847_inst_req_1;
      type_cast_847_inst_ack_1<= rack(0);
      type_cast_847_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_847_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call175_844,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv177_848,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_865_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_865_inst_req_0;
      type_cast_865_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_865_inst_req_1;
      type_cast_865_inst_ack_1<= rack(0);
      type_cast_865_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_865_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call181_862,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv183_866,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_883_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_883_inst_req_0;
      type_cast_883_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_883_inst_req_1;
      type_cast_883_inst_ack_1<= rack(0);
      type_cast_883_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_883_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call187_880,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv189_884,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_901_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_901_inst_req_0;
      type_cast_901_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_901_inst_req_1;
      type_cast_901_inst_ack_1<= rack(0);
      type_cast_901_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_901_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call193_898,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv195_902,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence STORE_padding_229_gather_scatter
    process(call42x_xlcssa_224) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := call42x_xlcssa_224;
      ov(7 downto 0) := iv;
      STORE_padding_229_data_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1040_index_1_rename
    process(R_indvar_1039_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_1039_resized;
      ov(13 downto 0) := iv;
      R_indvar_1039_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1040_index_1_resize
    process(indvar_1028) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_1028;
      ov := iv(13 downto 0);
      R_indvar_1039_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1040_root_address_inst
    process(array_obj_ref_1040_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1040_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1040_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_119_index_1_rename
    process(R_indvar280_118_resized) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar280_118_resized;
      ov(6 downto 0) := iv;
      R_indvar280_118_scaled <= ov(6 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_119_index_1_resize
    process(indvar280_107) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar280_107;
      ov := iv(6 downto 0);
      R_indvar280_118_resized <= ov(6 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_119_root_address_inst
    process(array_obj_ref_119_final_offset) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_119_final_offset;
      ov(6 downto 0) := iv;
      array_obj_ref_119_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_195_index_0_rename
    process(R_indvar277_194_resized) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar277_194_resized;
      ov(0 downto 0) := iv;
      R_indvar277_194_scaled <= ov(0 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_195_index_0_resize
    process(indvar277_179) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar277_179;
      ov := iv(0 downto 0);
      R_indvar277_194_resized <= ov(0 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_195_index_offset
    process(R_indvar277_194_scaled) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar277_194_scaled;
      ov(0 downto 0) := iv;
      array_obj_ref_195_final_offset <= ov(0 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_195_root_address_inst
    process(array_obj_ref_195_final_offset) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_195_final_offset;
      ov(0 downto 0) := iv;
      array_obj_ref_195_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_49_index_1_rename
    process(R_indvar283_48_resized) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar283_48_resized;
      ov(6 downto 0) := iv;
      R_indvar283_48_scaled <= ov(6 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_49_index_1_resize
    process(indvar283_37) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar283_37;
      ov := iv(6 downto 0);
      R_indvar283_48_resized <= ov(6 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_49_root_address_inst
    process(array_obj_ref_49_final_offset) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_49_final_offset;
      ov(6 downto 0) := iv;
      array_obj_ref_49_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_565_index_1_rename
    process(R_indvar265_564_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar265_564_resized;
      ov(13 downto 0) := iv;
      R_indvar265_564_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_565_index_1_resize
    process(indvar265_553) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar265_553;
      ov := iv(13 downto 0);
      R_indvar265_564_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_565_root_address_inst
    process(array_obj_ref_565_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_565_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_565_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_772_index_1_rename
    process(R_indvar253_771_resized) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar253_771_resized;
      ov(10 downto 0) := iv;
      R_indvar253_771_scaled <= ov(10 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_772_index_1_resize
    process(indvar253_760) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar253_760;
      ov := iv(10 downto 0);
      R_indvar253_771_resized <= ov(10 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_772_root_address_inst
    process(array_obj_ref_772_final_offset) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_772_final_offset;
      ov(10 downto 0) := iv;
      array_obj_ref_772_root_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1044_addr_0
    process(ptr_deref_1044_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1044_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1044_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1044_base_resize
    process(arrayidx220_1042) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx220_1042;
      ov := iv(13 downto 0);
      ptr_deref_1044_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1044_gather_scatter
    process(type_cast_1046_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_1046_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_1044_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1044_root_address_inst
    process(ptr_deref_1044_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1044_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1044_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_130_addr_0
    process(ptr_deref_130_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_130_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_130_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_130_base_resize
    process(arrayidx32_121) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx32_121;
      ov := iv(6 downto 0);
      ptr_deref_130_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_130_gather_scatter
    process(conv18_128) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv18_128;
      ov(31 downto 0) := iv;
      ptr_deref_130_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_130_root_address_inst
    process(ptr_deref_130_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_130_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_130_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_152_addr_0
    process(ptr_deref_152_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_152_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_152_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_152_base_resize
    process(arrayidx32_121) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx32_121;
      ov := iv(6 downto 0);
      ptr_deref_152_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_152_gather_scatter
    process(add29_150) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add29_150;
      ov(31 downto 0) := iv;
      ptr_deref_152_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_152_root_address_inst
    process(ptr_deref_152_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_152_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_152_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_199_addr_0
    process(ptr_deref_199_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_199_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_199_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_199_base_resize
    process(arrayidx45_197) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx45_197;
      ov := iv(0 downto 0);
      ptr_deref_199_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_199_gather_scatter
    process(call42239_186) --
      variable iv : std_logic_vector(7 downto 0);
      variable ov : std_logic_vector(7 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := call42239_186;
      ov(7 downto 0) := iv;
      ptr_deref_199_data_0 <= ov(7 downto 0);
      --
    end process;
    -- equivalence ptr_deref_199_root_address_inst
    process(ptr_deref_199_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_199_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_199_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_248_addr_0
    process(ptr_deref_248_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_248_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_248_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_248_base_resize
    process(iNsTr_19_246) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_19_246;
      ov := iv(6 downto 0);
      ptr_deref_248_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_248_gather_scatter
    process(conv52_238) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv52_238;
      ov(31 downto 0) := iv;
      ptr_deref_248_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_248_root_address_inst
    process(ptr_deref_248_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_248_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_248_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_278_addr_0
    process(ptr_deref_278_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_278_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_278_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_278_base_resize
    process(iNsTr_22_276) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_22_276;
      ov := iv(6 downto 0);
      ptr_deref_278_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_278_gather_scatter
    process(add57_268) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add57_268;
      ov(31 downto 0) := iv;
      ptr_deref_278_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_278_root_address_inst
    process(ptr_deref_278_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_278_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_278_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_297_addr_0
    process(ptr_deref_297_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_297_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_297_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_297_base_resize
    process(iNsTr_25_295) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_25_295;
      ov := iv(6 downto 0);
      ptr_deref_297_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_297_gather_scatter
    process(conv59_287) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv59_287;
      ov(31 downto 0) := iv;
      ptr_deref_297_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_297_root_address_inst
    process(ptr_deref_297_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_297_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_297_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_327_addr_0
    process(ptr_deref_327_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_327_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_327_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_327_base_resize
    process(iNsTr_28_325) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_28_325;
      ov := iv(6 downto 0);
      ptr_deref_327_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_327_gather_scatter
    process(add64_317) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add64_317;
      ov(31 downto 0) := iv;
      ptr_deref_327_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_327_root_address_inst
    process(ptr_deref_327_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_327_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_327_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_346_addr_0
    process(ptr_deref_346_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_346_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_346_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_346_base_resize
    process(iNsTr_31_344) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_31_344;
      ov := iv(6 downto 0);
      ptr_deref_346_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_346_gather_scatter
    process(conv66_336) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv66_336;
      ov(31 downto 0) := iv;
      ptr_deref_346_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_346_root_address_inst
    process(ptr_deref_346_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_346_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_346_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_376_addr_0
    process(ptr_deref_376_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_376_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_376_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_376_base_resize
    process(iNsTr_34_374) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_34_374;
      ov := iv(6 downto 0);
      ptr_deref_376_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_376_gather_scatter
    process(add71_366) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add71_366;
      ov(31 downto 0) := iv;
      ptr_deref_376_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_376_root_address_inst
    process(ptr_deref_376_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_376_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_376_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_389_addr_0
    process(ptr_deref_389_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_389_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_389_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_389_base_resize
    process(iNsTr_36_386) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_36_386;
      ov := iv(6 downto 0);
      ptr_deref_389_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_389_gather_scatter
    process(ptr_deref_389_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_389_data_0;
      ov(31 downto 0) := iv;
      tmp73_390 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_389_root_address_inst
    process(ptr_deref_389_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_389_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_389_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_401_addr_0
    process(ptr_deref_401_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_401_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_401_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_401_base_resize
    process(iNsTr_37_398) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_37_398;
      ov := iv(6 downto 0);
      ptr_deref_401_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_401_gather_scatter
    process(ptr_deref_401_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_401_data_0;
      ov(31 downto 0) := iv;
      tmp74_402 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_401_root_address_inst
    process(ptr_deref_401_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_401_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_401_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_413_addr_0
    process(ptr_deref_413_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_413_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_413_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_413_base_resize
    process(iNsTr_38_410) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_38_410;
      ov := iv(6 downto 0);
      ptr_deref_413_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_413_gather_scatter
    process(ptr_deref_413_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_413_data_0;
      ov(31 downto 0) := iv;
      tmp75_414 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_413_root_address_inst
    process(ptr_deref_413_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_413_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_413_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_435_addr_0
    process(ptr_deref_435_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_435_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_435_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_435_base_resize
    process(iNsTr_39_432) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_39_432;
      ov := iv(6 downto 0);
      ptr_deref_435_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_435_gather_scatter
    process(ptr_deref_435_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_435_data_0;
      ov(31 downto 0) := iv;
      tmp78_436 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_435_root_address_inst
    process(ptr_deref_435_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_435_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_435_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_447_addr_0
    process(ptr_deref_447_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_447_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_447_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_447_base_resize
    process(iNsTr_40_444) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_40_444;
      ov := iv(6 downto 0);
      ptr_deref_447_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_447_gather_scatter
    process(ptr_deref_447_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_447_data_0;
      ov(31 downto 0) := iv;
      tmp79_448 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_447_root_address_inst
    process(ptr_deref_447_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_447_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_447_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_459_addr_0
    process(ptr_deref_459_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_459_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_459_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_459_base_resize
    process(iNsTr_41_456) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_41_456;
      ov := iv(6 downto 0);
      ptr_deref_459_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_459_gather_scatter
    process(ptr_deref_459_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_459_data_0;
      ov(31 downto 0) := iv;
      tmp81_460 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_459_root_address_inst
    process(ptr_deref_459_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_459_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_459_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_471_addr_0
    process(ptr_deref_471_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_471_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_471_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_471_base_resize
    process(iNsTr_42_468) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_42_468;
      ov := iv(6 downto 0);
      ptr_deref_471_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_471_gather_scatter
    process(ptr_deref_471_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_471_data_0;
      ov(31 downto 0) := iv;
      tmp83_472 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_471_root_address_inst
    process(ptr_deref_471_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_471_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_471_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_60_addr_0
    process(ptr_deref_60_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_60_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_60_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_60_base_resize
    process(arrayidx10_51) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx10_51;
      ov := iv(6 downto 0);
      ptr_deref_60_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_60_gather_scatter
    process(conv_58) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv_58;
      ov(31 downto 0) := iv;
      ptr_deref_60_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_60_root_address_inst
    process(ptr_deref_60_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_60_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_60_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_702_addr_0
    process(ptr_deref_702_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_702_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_702_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_702_base_resize
    process(arrayidx139_567) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx139_567;
      ov := iv(13 downto 0);
      ptr_deref_702_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_702_gather_scatter
    process(add135_700) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add135_700;
      ov(63 downto 0) := iv;
      ptr_deref_702_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_702_root_address_inst
    process(ptr_deref_702_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_702_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_702_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_82_addr_0
    process(ptr_deref_82_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_82_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_82_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_82_base_resize
    process(arrayidx10_51) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx10_51;
      ov := iv(6 downto 0);
      ptr_deref_82_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_82_gather_scatter
    process(add_80) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add_80;
      ov(31 downto 0) := iv;
      ptr_deref_82_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_82_root_address_inst
    process(ptr_deref_82_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_82_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_82_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_909_addr_0
    process(ptr_deref_909_root_address) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_909_root_address;
      ov(10 downto 0) := iv;
      ptr_deref_909_word_address_0 <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_909_base_resize
    process(arrayidx200_774) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx200_774;
      ov := iv(10 downto 0);
      ptr_deref_909_resized_base_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_909_gather_scatter
    process(add196_907) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add196_907;
      ov(63 downto 0) := iv;
      ptr_deref_909_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_909_root_address_inst
    process(ptr_deref_909_resized_base_address) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_909_resized_base_address;
      ov(10 downto 0) := iv;
      ptr_deref_909_root_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_942_addr_0
    process(ptr_deref_942_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_942_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_942_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_942_base_resize
    process(iNsTr_59_939) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_59_939;
      ov := iv(6 downto 0);
      ptr_deref_942_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_942_gather_scatter
    process(ptr_deref_942_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_942_data_0;
      ov(31 downto 0) := iv;
      tmp206_943 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_942_root_address_inst
    process(ptr_deref_942_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_942_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_942_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_954_addr_0
    process(ptr_deref_954_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_954_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_954_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_954_base_resize
    process(iNsTr_60_951) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_60_951;
      ov := iv(6 downto 0);
      ptr_deref_954_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_954_gather_scatter
    process(ptr_deref_954_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_954_data_0;
      ov(31 downto 0) := iv;
      tmp207_955 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_954_root_address_inst
    process(ptr_deref_954_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_954_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_954_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_966_addr_0
    process(ptr_deref_966_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_966_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_966_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_966_base_resize
    process(iNsTr_61_963) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_61_963;
      ov := iv(6 downto 0);
      ptr_deref_966_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_966_gather_scatter
    process(ptr_deref_966_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_966_data_0;
      ov(31 downto 0) := iv;
      tmp209_967 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_966_root_address_inst
    process(ptr_deref_966_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_966_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_966_root_address <= ov(6 downto 0);
      --
    end process;
    if_stmt_1059_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond1_1058;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1059_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1059_branch_req_0,
          ack0 => if_stmt_1059_branch_ack_0,
          ack1 => if_stmt_1059_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_167_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond4_166;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_167_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_167_branch_req_0,
          ack0 => if_stmt_167_branch_ack_0,
          ack1 => if_stmt_167_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_217_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond3_216;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_217_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_217_branch_req_0,
          ack0 => if_stmt_217_branch_ack_0,
          ack1 => if_stmt_217_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_494_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp88233_493;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_494_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_494_branch_req_0,
          ack0 => if_stmt_494_branch_ack_0,
          ack1 => if_stmt_494_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_509_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp148229_508;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_509_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_509_branch_req_0,
          ack0 => if_stmt_509_branch_ack_0,
          ack1 => if_stmt_509_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_716_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond2_715;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_716_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_716_branch_req_0,
          ack0 => if_stmt_716_branch_ack_0,
          ack1 => if_stmt_716_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_923_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond_922;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_923_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_923_branch_req_0,
          ack0 => if_stmt_923_branch_ack_0,
          ack1 => if_stmt_923_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_984_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp215226_983;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_984_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_984_branch_req_0,
          ack0 => if_stmt_984_branch_ack_0,
          ack1 => if_stmt_984_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_98_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond5_97;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_98_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_98_branch_req_0,
          ack0 => if_stmt_98_branch_ack_0,
          ack1 => if_stmt_98_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u32_u32_1007_inst
    process(tmp248_996) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp248_996, type_cast_1006_wire_constant, tmp_var);
      tmp248x_xop_1008 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_532_inst
    process(tmp269_521) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp269_521, type_cast_531_wire_constant, tmp_var);
      tmp269x_xop_533 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_739_inst
    process(tmp258_728) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp258_728, type_cast_738_wire_constant, tmp_var);
      tmp258x_xop_740 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1017_inst
    process(iNsTr_74_1012) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_74_1012, type_cast_1016_wire_constant, tmp_var);
      xx_xop_1018 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1052_inst
    process(indvar_1028) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1028, type_cast_1051_wire_constant, tmp_var);
      indvarx_xnext_1053 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_159_inst
    process(indvar280_107) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar280_107, type_cast_158_wire_constant, tmp_var);
      indvarx_xnext281_160 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_209_inst
    process(indvar277_179) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar277_179, type_cast_208_wire_constant, tmp_var);
      indvarx_xnext278_210 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_542_inst
    process(iNsTr_44_537) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_44_537, type_cast_541_wire_constant, tmp_var);
      xx_xop287_543 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_709_inst
    process(indvar265_553) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar265_553, type_cast_708_wire_constant, tmp_var);
      indvarx_xnext266_710 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_749_inst
    process(iNsTr_57_744) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_57_744, type_cast_748_wire_constant, tmp_var);
      xx_xop286_750 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_89_inst
    process(indvar283_37) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar283_37, type_cast_88_wire_constant, tmp_var);
      indvarx_xnext284_90 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_916_inst
    process(indvar253_760) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar253_760, type_cast_915_wire_constant, tmp_var);
      indvarx_xnext254_917 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1057_inst
    process(indvarx_xnext_1053, tmp252_1025) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_1053, tmp252_1025, tmp_var);
      exitcond1_1058 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_165_inst
    process(indvarx_xnext281_160) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext281_160, type_cast_164_wire_constant, tmp_var);
      exitcond4_166 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_215_inst
    process(indvarx_xnext278_210) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext278_210, type_cast_214_wire_constant, tmp_var);
      exitcond3_216 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_714_inst
    process(indvarx_xnext266_710, tmp274_550) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext266_710, tmp274_550, tmp_var);
      exitcond2_715 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_921_inst
    process(indvarx_xnext254_917, tmp263_757) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext254_917, tmp263_757, tmp_var);
      exitcond_922 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_95_inst
    process(indvarx_xnext284_90) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext284_90, type_cast_94_wire_constant, tmp_var);
      exitcond5_97 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_520_inst
    process(mul76_424) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul76_424, type_cast_519_wire_constant, tmp_var);
      tmp269_521 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_727_inst
    process(mul84_487) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul84_487, type_cast_726_wire_constant, tmp_var);
      tmp258_728 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_995_inst
    process(mul210_977) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul210_977, type_cast_994_wire_constant, tmp_var);
      tmp248_996 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_418_inst
    process(tmp74_402, tmp73_390) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp74_402, tmp73_390, tmp_var);
      mul_419 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_423_inst
    process(mul_419, tmp75_414) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_419, tmp75_414, tmp_var);
      mul76_424 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_476_inst
    process(tmp79_448, tmp78_436) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp79_448, tmp78_436, tmp_var);
      mul80_477 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_481_inst
    process(mul80_477, tmp81_460) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul80_477, tmp81_460, tmp_var);
      mul82_482 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_486_inst
    process(mul82_482, tmp83_472) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul82_482, tmp83_472, tmp_var);
      mul84_487 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_971_inst
    process(tmp207_955, tmp206_943) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp207_955, tmp206_943, tmp_var);
      mul208_972 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_976_inst
    process(mul208_972, tmp209_967) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul208_972, tmp209_967, tmp_var);
      mul210_977 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_149_inst
    process(conv28_145, shl26_138) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv28_145, shl26_138, tmp_var);
      add29_150 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_267_inst
    process(shl54_256, conv56_263) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl54_256, conv56_263, tmp_var);
      add57_268 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_316_inst
    process(shl61_305, conv63_312) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl61_305, conv63_312, tmp_var);
      add64_317 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_365_inst
    process(shl68_354, conv70_361) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl68_354, conv70_361, tmp_var);
      add71_366 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_79_inst
    process(conv7_75, shl_68) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv7_75, shl_68, tmp_var);
      add_80 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_591_inst
    process(shl95_580, conv98_587) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl95_580, conv98_587, tmp_var);
      add99_592 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_609_inst
    process(shl101_598, conv104_605) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl101_598, conv104_605, tmp_var);
      add105_610 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_627_inst
    process(shl107_616, conv110_623) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl107_616, conv110_623, tmp_var);
      add111_628 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_645_inst
    process(shl113_634, conv116_641) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl113_634, conv116_641, tmp_var);
      add117_646 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_663_inst
    process(shl119_652, conv122_659) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl119_652, conv122_659, tmp_var);
      add123_664 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_681_inst
    process(shl125_670, conv128_677) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl125_670, conv128_677, tmp_var);
      add129_682 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_699_inst
    process(shl131_688, conv134_695) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl131_688, conv134_695, tmp_var);
      add135_700 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_798_inst
    process(shl156_787, conv159_794) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl156_787, conv159_794, tmp_var);
      add160_799 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_816_inst
    process(shl162_805, conv165_812) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl162_805, conv165_812, tmp_var);
      add166_817 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_834_inst
    process(shl168_823, conv171_830) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl168_823, conv171_830, tmp_var);
      add172_835 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_852_inst
    process(shl174_841, conv177_848) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl174_841, conv177_848, tmp_var);
      add178_853 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_870_inst
    process(shl180_859, conv183_866) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl180_859, conv183_866, tmp_var);
      add184_871 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_888_inst
    process(shl186_877, conv189_884) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl186_877, conv189_884, tmp_var);
      add190_889 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_906_inst
    process(shl192_895, conv195_902) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl192_895, conv195_902, tmp_var);
      add196_907 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_137_inst
    process(conv18_128) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv18_128, type_cast_136_wire_constant, tmp_var);
      shl26_138 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_255_inst
    process(conv52_238) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv52_238, type_cast_254_wire_constant, tmp_var);
      shl54_256 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_304_inst
    process(conv59_287) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv59_287, type_cast_303_wire_constant, tmp_var);
      shl61_305 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_353_inst
    process(conv66_336) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv66_336, type_cast_352_wire_constant, tmp_var);
      shl68_354 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_67_inst
    process(conv_58) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv_58, type_cast_66_wire_constant, tmp_var);
      shl_68 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_579_inst
    process(conv93_574) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv93_574, type_cast_578_wire_constant, tmp_var);
      shl95_580 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_597_inst
    process(add99_592) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add99_592, type_cast_596_wire_constant, tmp_var);
      shl101_598 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_615_inst
    process(add105_610) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add105_610, type_cast_614_wire_constant, tmp_var);
      shl107_616 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_633_inst
    process(add111_628) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add111_628, type_cast_632_wire_constant, tmp_var);
      shl113_634 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_651_inst
    process(add117_646) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add117_646, type_cast_650_wire_constant, tmp_var);
      shl119_652 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_669_inst
    process(add123_664) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add123_664, type_cast_668_wire_constant, tmp_var);
      shl125_670 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_687_inst
    process(add129_682) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add129_682, type_cast_686_wire_constant, tmp_var);
      shl131_688 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_786_inst
    process(conv154_781) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv154_781, type_cast_785_wire_constant, tmp_var);
      shl156_787 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_804_inst
    process(add160_799) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add160_799, type_cast_803_wire_constant, tmp_var);
      shl162_805 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_822_inst
    process(add166_817) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add166_817, type_cast_821_wire_constant, tmp_var);
      shl168_823 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_840_inst
    process(add172_835) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add172_835, type_cast_839_wire_constant, tmp_var);
      shl174_841 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_858_inst
    process(add178_853) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add178_853, type_cast_857_wire_constant, tmp_var);
      shl180_859 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_876_inst
    process(add184_871) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add184_871, type_cast_875_wire_constant, tmp_var);
      shl186_877 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_894_inst
    process(add190_889) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add190_889, type_cast_893_wire_constant, tmp_var);
      shl192_895 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1001_inst
    process(tmp248_996) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp248_996, type_cast_1000_wire_constant, tmp_var);
      tmp249_1002 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_492_inst
    process(mul76_424) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul76_424, type_cast_491_wire_constant, tmp_var);
      cmp88233_493 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_507_inst
    process(mul84_487) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul84_487, type_cast_506_wire_constant, tmp_var);
      cmp148229_508 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_526_inst
    process(tmp269_521) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp269_521, type_cast_525_wire_constant, tmp_var);
      tmp270_527 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_733_inst
    process(tmp258_728) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp258_728, type_cast_732_wire_constant, tmp_var);
      tmp259_734 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_982_inst
    process(mul210_977) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul210_977, type_cast_981_wire_constant, tmp_var);
      cmp215226_983 <= tmp_var; --
    end process;
    -- shared split operator group (72) : array_obj_ref_1040_index_offset 
    ApIntAdd_group_72: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_1039_scaled;
      array_obj_ref_1040_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1040_index_offset_req_0;
      array_obj_ref_1040_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1040_index_offset_req_1;
      array_obj_ref_1040_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_72_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_72_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_72",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 72
    -- shared split operator group (73) : array_obj_ref_119_index_offset 
    ApIntAdd_group_73: Block -- 
      signal data_in: std_logic_vector(6 downto 0);
      signal data_out: std_logic_vector(6 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar280_118_scaled;
      array_obj_ref_119_final_offset <= data_out(6 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_119_index_offset_req_0;
      array_obj_ref_119_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_119_index_offset_req_1;
      array_obj_ref_119_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_73_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_73_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_73",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 7,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 7,
          constant_operand => "0000011",
          constant_width => 7,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 73
    -- shared split operator group (74) : array_obj_ref_49_index_offset 
    ApIntAdd_group_74: Block -- 
      signal data_in: std_logic_vector(6 downto 0);
      signal data_out: std_logic_vector(6 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar283_48_scaled;
      array_obj_ref_49_final_offset <= data_out(6 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_49_index_offset_req_0;
      array_obj_ref_49_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_49_index_offset_req_1;
      array_obj_ref_49_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_74_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_74_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_74",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 7,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 7,
          constant_operand => "0000011",
          constant_width => 7,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 74
    -- shared split operator group (75) : array_obj_ref_565_index_offset 
    ApIntAdd_group_75: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar265_564_scaled;
      array_obj_ref_565_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_565_index_offset_req_0;
      array_obj_ref_565_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_565_index_offset_req_1;
      array_obj_ref_565_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_75_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_75_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_75",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 75
    -- shared split operator group (76) : array_obj_ref_772_index_offset 
    ApIntAdd_group_76: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar253_771_scaled;
      array_obj_ref_772_final_offset <= data_out(10 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_772_index_offset_req_0;
      array_obj_ref_772_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_772_index_offset_req_1;
      array_obj_ref_772_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_76_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_76_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_76",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000100010",
          constant_width => 11,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 76
    -- shared load operator group (0) : ptr_deref_401_load_0 ptr_deref_413_load_0 ptr_deref_389_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(20 downto 0);
      signal data_out: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_401_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_413_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_389_load_0_req_0;
      ptr_deref_401_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_413_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_389_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_401_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_413_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_389_load_0_req_1;
      ptr_deref_401_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_413_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_389_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_401_word_address_0 & ptr_deref_413_word_address_0 & ptr_deref_389_word_address_0;
      ptr_deref_401_data_0 <= data_out(95 downto 64);
      ptr_deref_413_data_0 <= data_out(63 downto 32);
      ptr_deref_389_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 7,
        num_reqs => 3,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(6 downto 0),
          mtag => memory_space_1_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 32,
        num_reqs => 3,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(31 downto 0),
          mtag => memory_space_1_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_471_load_0 ptr_deref_435_load_0 ptr_deref_459_load_0 ptr_deref_447_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(27 downto 0);
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 3 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 3 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 3 downto 0);
      signal guard_vector : std_logic_vector( 3 downto 0);
      constant inBUFs : IntegerArray(3 downto 0) := (3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(3 downto 0) := (3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(3 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false);
      constant guardBuffering: IntegerArray(3 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2);
      -- 
    begin -- 
      reqL_unguarded(3) <= ptr_deref_471_load_0_req_0;
      reqL_unguarded(2) <= ptr_deref_435_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_459_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_447_load_0_req_0;
      ptr_deref_471_load_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_435_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_459_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_447_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(3) <= ptr_deref_471_load_0_req_1;
      reqR_unguarded(2) <= ptr_deref_435_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_459_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_447_load_0_req_1;
      ptr_deref_471_load_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_435_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_459_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_447_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      LoadGroup1_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 4, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_471_word_address_0 & ptr_deref_435_word_address_0 & ptr_deref_459_word_address_0 & ptr_deref_447_word_address_0;
      ptr_deref_471_data_0 <= data_out(127 downto 96);
      ptr_deref_435_data_0 <= data_out(95 downto 64);
      ptr_deref_459_data_0 <= data_out(63 downto 32);
      ptr_deref_447_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 7,
        num_reqs => 4,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(6 downto 0),
          mtag => memory_space_2_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 32,
        num_reqs => 4,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(31 downto 0),
          mtag => memory_space_2_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : ptr_deref_954_load_0 ptr_deref_942_load_0 ptr_deref_966_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(20 downto 0);
      signal data_out: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_954_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_942_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_966_load_0_req_0;
      ptr_deref_954_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_942_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_966_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_954_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_942_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_966_load_0_req_1;
      ptr_deref_954_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_942_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_966_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      LoadGroup2_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup2_gI: SplitGuardInterface generic map(name => "LoadGroup2_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_954_word_address_0 & ptr_deref_942_word_address_0 & ptr_deref_966_word_address_0;
      ptr_deref_954_data_0 <= data_out(95 downto 64);
      ptr_deref_942_data_0 <= data_out(63 downto 32);
      ptr_deref_966_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup2", addr_width => 7,
        num_reqs => 3,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(6 downto 0),
          mtag => memory_space_3_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup2 load-complete ",
        data_width => 32,
        num_reqs => 3,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(31 downto 0),
          mtag => memory_space_3_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared store operator group (0) : STORE_padding_229_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= STORE_padding_229_store_0_req_0;
      STORE_padding_229_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= STORE_padding_229_store_0_req_1;
      STORE_padding_229_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_padding_229_word_address_0;
      data_in <= STORE_padding_229_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 1,
        data_width => 8,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_7_sr_req(0),
          mack => memory_space_7_sr_ack(0),
          maddr => memory_space_7_sr_addr(0 downto 0),
          mdata => memory_space_7_sr_data(7 downto 0),
          mtag => memory_space_7_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_7_sc_req(0),
          mack => memory_space_7_sc_ack(0),
          mtag => memory_space_7_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : ptr_deref_1044_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1044_store_0_req_0;
      ptr_deref_1044_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1044_store_0_req_1;
      ptr_deref_1044_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup1_gI: SplitGuardInterface generic map(name => "StoreGroup1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1044_word_address_0;
      data_in <= ptr_deref_1044_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup1 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_6_sr_req(0),
          mack => memory_space_6_sr_ack(0),
          maddr => memory_space_6_sr_addr(13 downto 0),
          mdata => memory_space_6_sr_data(63 downto 0),
          mtag => memory_space_6_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup1 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_6_sc_req(0),
          mack => memory_space_6_sc_ack(0),
          mtag => memory_space_6_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared store operator group (2) : ptr_deref_130_store_0 ptr_deref_152_store_0 
    StoreGroup2: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_130_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_152_store_0_req_0;
      ptr_deref_130_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_152_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_130_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_152_store_0_req_1;
      ptr_deref_130_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_152_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup2_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup2_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup2_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup2_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup2_gI: SplitGuardInterface generic map(name => "StoreGroup2_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_130_word_address_0 & ptr_deref_152_word_address_0;
      data_in <= ptr_deref_130_data_0 & ptr_deref_152_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup2 Req ", addr_width => 7,
        data_width => 32,
        num_reqs => 2,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(6 downto 0),
          mdata => memory_space_2_sr_data(31 downto 0),
          mtag => memory_space_2_sr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup2 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 2
    -- shared store operator group (3) : ptr_deref_199_store_0 
    StoreGroup3: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_199_store_0_req_0;
      ptr_deref_199_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_199_store_0_req_1;
      ptr_deref_199_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup3_gI: SplitGuardInterface generic map(name => "StoreGroup3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_199_word_address_0;
      data_in <= ptr_deref_199_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup3 Req ", addr_width => 1,
        data_width => 8,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_8_sr_req(0),
          mack => memory_space_8_sr_ack(0),
          maddr => memory_space_8_sr_addr(0 downto 0),
          mdata => memory_space_8_sr_data(7 downto 0),
          mtag => memory_space_8_sr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup3 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_8_sc_req(0),
          mack => memory_space_8_sc_ack(0),
          mtag => memory_space_8_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 3
    -- shared store operator group (4) : ptr_deref_346_store_0 ptr_deref_376_store_0 ptr_deref_327_store_0 ptr_deref_297_store_0 ptr_deref_278_store_0 ptr_deref_248_store_0 
    StoreGroup4: Block -- 
      signal addr_in: std_logic_vector(41 downto 0);
      signal data_in: std_logic_vector(191 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 5 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 5 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 5 downto 0);
      signal guard_vector : std_logic_vector( 5 downto 0);
      constant inBUFs : IntegerArray(5 downto 0) := (5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(5 downto 0) := (5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(5 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false);
      constant guardBuffering: IntegerArray(5 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2);
      -- 
    begin -- 
      reqL_unguarded(5) <= ptr_deref_346_store_0_req_0;
      reqL_unguarded(4) <= ptr_deref_376_store_0_req_0;
      reqL_unguarded(3) <= ptr_deref_327_store_0_req_0;
      reqL_unguarded(2) <= ptr_deref_297_store_0_req_0;
      reqL_unguarded(1) <= ptr_deref_278_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_248_store_0_req_0;
      ptr_deref_346_store_0_ack_0 <= ackL_unguarded(5);
      ptr_deref_376_store_0_ack_0 <= ackL_unguarded(4);
      ptr_deref_327_store_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_297_store_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_278_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_248_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(5) <= ptr_deref_346_store_0_req_1;
      reqR_unguarded(4) <= ptr_deref_376_store_0_req_1;
      reqR_unguarded(3) <= ptr_deref_327_store_0_req_1;
      reqR_unguarded(2) <= ptr_deref_297_store_0_req_1;
      reqR_unguarded(1) <= ptr_deref_278_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_248_store_0_req_1;
      ptr_deref_346_store_0_ack_1 <= ackR_unguarded(5);
      ptr_deref_376_store_0_ack_1 <= ackR_unguarded(4);
      ptr_deref_327_store_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_297_store_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_278_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_248_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      StoreGroup4_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup4_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup4_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup4_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup4_accessRegulator_2: access_regulator_base generic map (name => "StoreGroup4_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      StoreGroup4_accessRegulator_3: access_regulator_base generic map (name => "StoreGroup4_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      StoreGroup4_accessRegulator_4: access_regulator_base generic map (name => "StoreGroup4_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      StoreGroup4_accessRegulator_5: access_regulator_base generic map (name => "StoreGroup4_accessRegulator_5", num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      StoreGroup4_gI: SplitGuardInterface generic map(name => "StoreGroup4_gI", nreqs => 6, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_346_word_address_0 & ptr_deref_376_word_address_0 & ptr_deref_327_word_address_0 & ptr_deref_297_word_address_0 & ptr_deref_278_word_address_0 & ptr_deref_248_word_address_0;
      data_in <= ptr_deref_346_data_0 & ptr_deref_376_data_0 & ptr_deref_327_data_0 & ptr_deref_297_data_0 & ptr_deref_278_data_0 & ptr_deref_248_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup4 Req ", addr_width => 7,
        data_width => 32,
        num_reqs => 6,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(6 downto 0),
          mdata => memory_space_3_sr_data(31 downto 0),
          mtag => memory_space_3_sr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup4 Complete ",
          num_reqs => 6,
          detailed_buffering_per_output => outBUFs,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 4
    -- shared store operator group (5) : ptr_deref_60_store_0 ptr_deref_82_store_0 
    StoreGroup5: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_60_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_82_store_0_req_0;
      ptr_deref_60_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_82_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_60_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_82_store_0_req_1;
      ptr_deref_60_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_82_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup5_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup5_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup5_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup5_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup5_gI: SplitGuardInterface generic map(name => "StoreGroup5_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_60_word_address_0 & ptr_deref_82_word_address_0;
      data_in <= ptr_deref_60_data_0 & ptr_deref_82_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup5 Req ", addr_width => 7,
        data_width => 32,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(6 downto 0),
          mdata => memory_space_1_sr_data(31 downto 0),
          mtag => memory_space_1_sr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup5 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 5
    -- shared store operator group (6) : ptr_deref_702_store_0 
    StoreGroup6: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_702_store_0_req_0;
      ptr_deref_702_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_702_store_0_req_1;
      ptr_deref_702_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup6_gI: SplitGuardInterface generic map(name => "StoreGroup6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_702_word_address_0;
      data_in <= ptr_deref_702_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup6 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_4_sr_req(0),
          mack => memory_space_4_sr_ack(0),
          maddr => memory_space_4_sr_addr(13 downto 0),
          mdata => memory_space_4_sr_data(63 downto 0),
          mtag => memory_space_4_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup6 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_4_sc_req(0),
          mack => memory_space_4_sc_ack(0),
          mtag => memory_space_4_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 6
    -- shared store operator group (7) : ptr_deref_909_store_0 
    StoreGroup7: Block -- 
      signal addr_in: std_logic_vector(10 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_909_store_0_req_0;
      ptr_deref_909_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_909_store_0_req_1;
      ptr_deref_909_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup7_gI: SplitGuardInterface generic map(name => "StoreGroup7_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_909_word_address_0;
      data_in <= ptr_deref_909_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup7 Req ", addr_width => 11,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 0,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_5_sr_req(0),
          mack => memory_space_5_sr_ack(0),
          maddr => memory_space_5_sr_addr(10 downto 0),
          mdata => memory_space_5_sr_data(63 downto 0),
          mtag => memory_space_5_sr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup7 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_5_sc_req(0),
          mack => memory_space_5_sc_ack(0),
          mtag => memory_space_5_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 7
    -- shared inport operator group (0) : RPIPE_ConvTranspose_input_pipe_307_inst RPIPE_ConvTranspose_input_pipe_776_inst RPIPE_ConvTranspose_input_pipe_690_inst RPIPE_ConvTranspose_input_pipe_582_inst RPIPE_ConvTranspose_input_pipe_807_inst RPIPE_ConvTranspose_input_pipe_600_inst RPIPE_ConvTranspose_input_pipe_879_inst RPIPE_ConvTranspose_input_pipe_618_inst RPIPE_ConvTranspose_input_pipe_636_inst RPIPE_ConvTranspose_input_pipe_861_inst RPIPE_ConvTranspose_input_pipe_331_inst RPIPE_ConvTranspose_input_pipe_356_inst RPIPE_ConvTranspose_input_pipe_569_inst RPIPE_ConvTranspose_input_pipe_654_inst RPIPE_ConvTranspose_input_pipe_897_inst RPIPE_ConvTranspose_input_pipe_825_inst RPIPE_ConvTranspose_input_pipe_789_inst RPIPE_ConvTranspose_input_pipe_843_inst RPIPE_ConvTranspose_input_pipe_672_inst RPIPE_ConvTranspose_input_pipe_53_inst RPIPE_ConvTranspose_input_pipe_70_inst RPIPE_ConvTranspose_input_pipe_123_inst RPIPE_ConvTranspose_input_pipe_140_inst RPIPE_ConvTranspose_input_pipe_175_inst RPIPE_ConvTranspose_input_pipe_203_inst RPIPE_ConvTranspose_input_pipe_233_inst RPIPE_ConvTranspose_input_pipe_282_inst RPIPE_ConvTranspose_input_pipe_258_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(223 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 27 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 27 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 27 downto 0);
      signal guard_vector : std_logic_vector( 27 downto 0);
      constant outBUFs : IntegerArray(27 downto 0) := (27 => 1, 26 => 1, 25 => 1, 24 => 1, 23 => 1, 22 => 1, 21 => 1, 20 => 1, 19 => 1, 18 => 1, 17 => 1, 16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(27 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false, 17 => false, 18 => false, 19 => false, 20 => false, 21 => false, 22 => false, 23 => false, 24 => false, 25 => false, 26 => false, 27 => false);
      constant guardBuffering: IntegerArray(27 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2, 17 => 2, 18 => 2, 19 => 2, 20 => 2, 21 => 2, 22 => 2, 23 => 2, 24 => 2, 25 => 2, 26 => 2, 27 => 2);
      -- 
    begin -- 
      reqL_unguarded(27) <= RPIPE_ConvTranspose_input_pipe_307_inst_req_0;
      reqL_unguarded(26) <= RPIPE_ConvTranspose_input_pipe_776_inst_req_0;
      reqL_unguarded(25) <= RPIPE_ConvTranspose_input_pipe_690_inst_req_0;
      reqL_unguarded(24) <= RPIPE_ConvTranspose_input_pipe_582_inst_req_0;
      reqL_unguarded(23) <= RPIPE_ConvTranspose_input_pipe_807_inst_req_0;
      reqL_unguarded(22) <= RPIPE_ConvTranspose_input_pipe_600_inst_req_0;
      reqL_unguarded(21) <= RPIPE_ConvTranspose_input_pipe_879_inst_req_0;
      reqL_unguarded(20) <= RPIPE_ConvTranspose_input_pipe_618_inst_req_0;
      reqL_unguarded(19) <= RPIPE_ConvTranspose_input_pipe_636_inst_req_0;
      reqL_unguarded(18) <= RPIPE_ConvTranspose_input_pipe_861_inst_req_0;
      reqL_unguarded(17) <= RPIPE_ConvTranspose_input_pipe_331_inst_req_0;
      reqL_unguarded(16) <= RPIPE_ConvTranspose_input_pipe_356_inst_req_0;
      reqL_unguarded(15) <= RPIPE_ConvTranspose_input_pipe_569_inst_req_0;
      reqL_unguarded(14) <= RPIPE_ConvTranspose_input_pipe_654_inst_req_0;
      reqL_unguarded(13) <= RPIPE_ConvTranspose_input_pipe_897_inst_req_0;
      reqL_unguarded(12) <= RPIPE_ConvTranspose_input_pipe_825_inst_req_0;
      reqL_unguarded(11) <= RPIPE_ConvTranspose_input_pipe_789_inst_req_0;
      reqL_unguarded(10) <= RPIPE_ConvTranspose_input_pipe_843_inst_req_0;
      reqL_unguarded(9) <= RPIPE_ConvTranspose_input_pipe_672_inst_req_0;
      reqL_unguarded(8) <= RPIPE_ConvTranspose_input_pipe_53_inst_req_0;
      reqL_unguarded(7) <= RPIPE_ConvTranspose_input_pipe_70_inst_req_0;
      reqL_unguarded(6) <= RPIPE_ConvTranspose_input_pipe_123_inst_req_0;
      reqL_unguarded(5) <= RPIPE_ConvTranspose_input_pipe_140_inst_req_0;
      reqL_unguarded(4) <= RPIPE_ConvTranspose_input_pipe_175_inst_req_0;
      reqL_unguarded(3) <= RPIPE_ConvTranspose_input_pipe_203_inst_req_0;
      reqL_unguarded(2) <= RPIPE_ConvTranspose_input_pipe_233_inst_req_0;
      reqL_unguarded(1) <= RPIPE_ConvTranspose_input_pipe_282_inst_req_0;
      reqL_unguarded(0) <= RPIPE_ConvTranspose_input_pipe_258_inst_req_0;
      RPIPE_ConvTranspose_input_pipe_307_inst_ack_0 <= ackL_unguarded(27);
      RPIPE_ConvTranspose_input_pipe_776_inst_ack_0 <= ackL_unguarded(26);
      RPIPE_ConvTranspose_input_pipe_690_inst_ack_0 <= ackL_unguarded(25);
      RPIPE_ConvTranspose_input_pipe_582_inst_ack_0 <= ackL_unguarded(24);
      RPIPE_ConvTranspose_input_pipe_807_inst_ack_0 <= ackL_unguarded(23);
      RPIPE_ConvTranspose_input_pipe_600_inst_ack_0 <= ackL_unguarded(22);
      RPIPE_ConvTranspose_input_pipe_879_inst_ack_0 <= ackL_unguarded(21);
      RPIPE_ConvTranspose_input_pipe_618_inst_ack_0 <= ackL_unguarded(20);
      RPIPE_ConvTranspose_input_pipe_636_inst_ack_0 <= ackL_unguarded(19);
      RPIPE_ConvTranspose_input_pipe_861_inst_ack_0 <= ackL_unguarded(18);
      RPIPE_ConvTranspose_input_pipe_331_inst_ack_0 <= ackL_unguarded(17);
      RPIPE_ConvTranspose_input_pipe_356_inst_ack_0 <= ackL_unguarded(16);
      RPIPE_ConvTranspose_input_pipe_569_inst_ack_0 <= ackL_unguarded(15);
      RPIPE_ConvTranspose_input_pipe_654_inst_ack_0 <= ackL_unguarded(14);
      RPIPE_ConvTranspose_input_pipe_897_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_ConvTranspose_input_pipe_825_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_ConvTranspose_input_pipe_789_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_ConvTranspose_input_pipe_843_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_ConvTranspose_input_pipe_672_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_ConvTranspose_input_pipe_53_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_ConvTranspose_input_pipe_70_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_ConvTranspose_input_pipe_123_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_ConvTranspose_input_pipe_140_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_ConvTranspose_input_pipe_175_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_ConvTranspose_input_pipe_203_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_ConvTranspose_input_pipe_233_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_ConvTranspose_input_pipe_282_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_ConvTranspose_input_pipe_258_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(27) <= RPIPE_ConvTranspose_input_pipe_307_inst_req_1;
      reqR_unguarded(26) <= RPIPE_ConvTranspose_input_pipe_776_inst_req_1;
      reqR_unguarded(25) <= RPIPE_ConvTranspose_input_pipe_690_inst_req_1;
      reqR_unguarded(24) <= RPIPE_ConvTranspose_input_pipe_582_inst_req_1;
      reqR_unguarded(23) <= RPIPE_ConvTranspose_input_pipe_807_inst_req_1;
      reqR_unguarded(22) <= RPIPE_ConvTranspose_input_pipe_600_inst_req_1;
      reqR_unguarded(21) <= RPIPE_ConvTranspose_input_pipe_879_inst_req_1;
      reqR_unguarded(20) <= RPIPE_ConvTranspose_input_pipe_618_inst_req_1;
      reqR_unguarded(19) <= RPIPE_ConvTranspose_input_pipe_636_inst_req_1;
      reqR_unguarded(18) <= RPIPE_ConvTranspose_input_pipe_861_inst_req_1;
      reqR_unguarded(17) <= RPIPE_ConvTranspose_input_pipe_331_inst_req_1;
      reqR_unguarded(16) <= RPIPE_ConvTranspose_input_pipe_356_inst_req_1;
      reqR_unguarded(15) <= RPIPE_ConvTranspose_input_pipe_569_inst_req_1;
      reqR_unguarded(14) <= RPIPE_ConvTranspose_input_pipe_654_inst_req_1;
      reqR_unguarded(13) <= RPIPE_ConvTranspose_input_pipe_897_inst_req_1;
      reqR_unguarded(12) <= RPIPE_ConvTranspose_input_pipe_825_inst_req_1;
      reqR_unguarded(11) <= RPIPE_ConvTranspose_input_pipe_789_inst_req_1;
      reqR_unguarded(10) <= RPIPE_ConvTranspose_input_pipe_843_inst_req_1;
      reqR_unguarded(9) <= RPIPE_ConvTranspose_input_pipe_672_inst_req_1;
      reqR_unguarded(8) <= RPIPE_ConvTranspose_input_pipe_53_inst_req_1;
      reqR_unguarded(7) <= RPIPE_ConvTranspose_input_pipe_70_inst_req_1;
      reqR_unguarded(6) <= RPIPE_ConvTranspose_input_pipe_123_inst_req_1;
      reqR_unguarded(5) <= RPIPE_ConvTranspose_input_pipe_140_inst_req_1;
      reqR_unguarded(4) <= RPIPE_ConvTranspose_input_pipe_175_inst_req_1;
      reqR_unguarded(3) <= RPIPE_ConvTranspose_input_pipe_203_inst_req_1;
      reqR_unguarded(2) <= RPIPE_ConvTranspose_input_pipe_233_inst_req_1;
      reqR_unguarded(1) <= RPIPE_ConvTranspose_input_pipe_282_inst_req_1;
      reqR_unguarded(0) <= RPIPE_ConvTranspose_input_pipe_258_inst_req_1;
      RPIPE_ConvTranspose_input_pipe_307_inst_ack_1 <= ackR_unguarded(27);
      RPIPE_ConvTranspose_input_pipe_776_inst_ack_1 <= ackR_unguarded(26);
      RPIPE_ConvTranspose_input_pipe_690_inst_ack_1 <= ackR_unguarded(25);
      RPIPE_ConvTranspose_input_pipe_582_inst_ack_1 <= ackR_unguarded(24);
      RPIPE_ConvTranspose_input_pipe_807_inst_ack_1 <= ackR_unguarded(23);
      RPIPE_ConvTranspose_input_pipe_600_inst_ack_1 <= ackR_unguarded(22);
      RPIPE_ConvTranspose_input_pipe_879_inst_ack_1 <= ackR_unguarded(21);
      RPIPE_ConvTranspose_input_pipe_618_inst_ack_1 <= ackR_unguarded(20);
      RPIPE_ConvTranspose_input_pipe_636_inst_ack_1 <= ackR_unguarded(19);
      RPIPE_ConvTranspose_input_pipe_861_inst_ack_1 <= ackR_unguarded(18);
      RPIPE_ConvTranspose_input_pipe_331_inst_ack_1 <= ackR_unguarded(17);
      RPIPE_ConvTranspose_input_pipe_356_inst_ack_1 <= ackR_unguarded(16);
      RPIPE_ConvTranspose_input_pipe_569_inst_ack_1 <= ackR_unguarded(15);
      RPIPE_ConvTranspose_input_pipe_654_inst_ack_1 <= ackR_unguarded(14);
      RPIPE_ConvTranspose_input_pipe_897_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_ConvTranspose_input_pipe_825_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_ConvTranspose_input_pipe_789_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_ConvTranspose_input_pipe_843_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_ConvTranspose_input_pipe_672_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_ConvTranspose_input_pipe_53_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_ConvTranspose_input_pipe_70_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_ConvTranspose_input_pipe_123_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_ConvTranspose_input_pipe_140_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_ConvTranspose_input_pipe_175_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_ConvTranspose_input_pipe_203_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_ConvTranspose_input_pipe_233_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_ConvTranspose_input_pipe_282_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_ConvTranspose_input_pipe_258_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      guard_vector(18)  <=  '1';
      guard_vector(19)  <=  '1';
      guard_vector(20)  <=  '1';
      guard_vector(21)  <=  '1';
      guard_vector(22)  <=  '1';
      guard_vector(23)  <=  '1';
      guard_vector(24)  <=  '1';
      guard_vector(25)  <=  '1';
      guard_vector(26)  <=  '1';
      guard_vector(27)  <=  '1';
      call62_308 <= data_out(223 downto 216);
      call153_777 <= data_out(215 downto 208);
      call132_691 <= data_out(207 downto 200);
      call96_583 <= data_out(199 downto 192);
      call163_808 <= data_out(191 downto 184);
      call102_601 <= data_out(183 downto 176);
      call187_880 <= data_out(175 downto 168);
      call108_619 <= data_out(167 downto 160);
      call114_637 <= data_out(159 downto 152);
      call181_862 <= data_out(151 downto 144);
      call65_332 <= data_out(143 downto 136);
      call69_357 <= data_out(135 downto 128);
      call92_570 <= data_out(127 downto 120);
      call120_655 <= data_out(119 downto 112);
      call193_898 <= data_out(111 downto 104);
      call169_826 <= data_out(103 downto 96);
      call157_790 <= data_out(95 downto 88);
      call175_844 <= data_out(87 downto 80);
      call126_673 <= data_out(79 downto 72);
      call_54 <= data_out(71 downto 64);
      call6_71 <= data_out(63 downto 56);
      call17_124 <= data_out(55 downto 48);
      call27_141 <= data_out(47 downto 40);
      call42237_176 <= data_out(39 downto 32);
      call42_204 <= data_out(31 downto 24);
      call51_234 <= data_out(23 downto 16);
      call58_283 <= data_out(15 downto 8);
      call55_259 <= data_out(7 downto 0);
      ConvTranspose_input_pipe_read_0_gI: SplitGuardInterface generic map(name => "ConvTranspose_input_pipe_read_0_gI", nreqs => 28, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      ConvTranspose_input_pipe_read_0: InputPortRevised -- 
        generic map ( name => "ConvTranspose_input_pipe_read_0", data_width => 8,  num_reqs => 28,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => ConvTranspose_input_pipe_pipe_read_req(0),
          oack => ConvTranspose_input_pipe_pipe_read_ack(0),
          odata => ConvTranspose_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- 
  end Block; -- data_path
  -- 
end testConfigure_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timer is -- 
  generic (tag_length : integer); 
  port ( -- 
    c : out  std_logic_vector(31 downto 0);
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(0 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timer;
architecture timer_arch of timer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 32)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal c_buffer :  std_logic_vector(31 downto 0);
  signal c_update_enable: Boolean;
  signal timer_CP_3083_start: Boolean;
  signal timer_CP_3083_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal LOAD_count_1079_load_0_req_0 : boolean;
  signal LOAD_count_1079_load_0_ack_0 : boolean;
  signal LOAD_count_1079_load_0_req_1 : boolean;
  signal LOAD_count_1079_load_0_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timer_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timer_CP_3083_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timer_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 32) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= c_buffer;
  c <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(tag_length + 31 downto 32) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 31 downto 32);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_3083_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timer_CP_3083_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_3083_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timer_CP_3083: Block -- control-path 
    signal timer_CP_3083_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    timer_CP_3083_elements(0) <= timer_CP_3083_start;
    timer_CP_3083_symbol <= timer_CP_3083_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_1080/$entry
      -- CP-element group 0: 	 assign_stmt_1080/LOAD_count_1079_sample_start_
      -- CP-element group 0: 	 assign_stmt_1080/LOAD_count_1079_update_start_
      -- CP-element group 0: 	 assign_stmt_1080/LOAD_count_1079_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_1080/LOAD_count_1079_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_1080/LOAD_count_1079_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_1080/LOAD_count_1079_Sample/word_access_start/$entry
      -- CP-element group 0: 	 assign_stmt_1080/LOAD_count_1079_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_1080/LOAD_count_1079_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 assign_stmt_1080/LOAD_count_1079_Update/$entry
      -- CP-element group 0: 	 assign_stmt_1080/LOAD_count_1079_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_1080/LOAD_count_1079_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_1080/LOAD_count_1079_Update/word_access_complete/word_0/cr
      -- 
    cr_3115_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3115_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_3083_elements(0), ack => LOAD_count_1079_load_0_req_1); -- 
    rr_3104_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3104_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_3083_elements(0), ack => LOAD_count_1079_load_0_req_0); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (5) 
      -- CP-element group 1: 	 assign_stmt_1080/LOAD_count_1079_sample_completed_
      -- CP-element group 1: 	 assign_stmt_1080/LOAD_count_1079_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_1080/LOAD_count_1079_Sample/word_access_start/$exit
      -- CP-element group 1: 	 assign_stmt_1080/LOAD_count_1079_Sample/word_access_start/word_0/$exit
      -- CP-element group 1: 	 assign_stmt_1080/LOAD_count_1079_Sample/word_access_start/word_0/ra
      -- 
    ra_3105_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_count_1079_load_0_ack_0, ack => timer_CP_3083_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (11) 
      -- CP-element group 2: 	 $exit
      -- CP-element group 2: 	 assign_stmt_1080/$exit
      -- CP-element group 2: 	 assign_stmt_1080/LOAD_count_1079_update_completed_
      -- CP-element group 2: 	 assign_stmt_1080/LOAD_count_1079_Update/$exit
      -- CP-element group 2: 	 assign_stmt_1080/LOAD_count_1079_Update/word_access_complete/$exit
      -- CP-element group 2: 	 assign_stmt_1080/LOAD_count_1079_Update/word_access_complete/word_0/$exit
      -- CP-element group 2: 	 assign_stmt_1080/LOAD_count_1079_Update/word_access_complete/word_0/ca
      -- CP-element group 2: 	 assign_stmt_1080/LOAD_count_1079_Update/LOAD_count_1079_Merge/$entry
      -- CP-element group 2: 	 assign_stmt_1080/LOAD_count_1079_Update/LOAD_count_1079_Merge/$exit
      -- CP-element group 2: 	 assign_stmt_1080/LOAD_count_1079_Update/LOAD_count_1079_Merge/merge_req
      -- CP-element group 2: 	 assign_stmt_1080/LOAD_count_1079_Update/LOAD_count_1079_Merge/merge_ack
      -- 
    ca_3116_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_count_1079_load_0_ack_1, ack => timer_CP_3083_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal LOAD_count_1079_data_0 : std_logic_vector(31 downto 0);
    signal LOAD_count_1079_word_address_0 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    LOAD_count_1079_word_address_0 <= "0";
    -- equivalence LOAD_count_1079_gather_scatter
    process(LOAD_count_1079_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_count_1079_data_0;
      ov(31 downto 0) := iv;
      c_buffer <= ov(31 downto 0);
      --
    end process;
    -- shared load operator group (0) : LOAD_count_1079_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_count_1079_load_0_req_0;
      LOAD_count_1079_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_count_1079_load_0_req_1;
      LOAD_count_1079_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_count_1079_word_address_0;
      LOAD_count_1079_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 0,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(0 downto 0),
          mtag => memory_space_0_lr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(31 downto 0),
          mtag => memory_space_0_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- 
  end Block; -- data_path
  -- 
end timer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    ConvTranspose_input_pipe_pipe_write_data: in std_logic_vector(7 downto 0);
    ConvTranspose_input_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_read_data: out std_logic_vector(7 downto 0);
    ConvTranspose_output_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_read_ack : out std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_read_data: out std_logic_vector(63 downto 0);
    elapsed_time_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(4 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(4 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(34 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(99 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(4 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(4 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(159 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(9 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(6 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(19 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(1 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_lr_req :  std_logic_vector(4 downto 0);
  signal memory_space_2_lr_ack : std_logic_vector(4 downto 0);
  signal memory_space_2_lr_addr : std_logic_vector(34 downto 0);
  signal memory_space_2_lr_tag : std_logic_vector(104 downto 0);
  signal memory_space_2_lc_req : std_logic_vector(4 downto 0);
  signal memory_space_2_lc_ack :  std_logic_vector(4 downto 0);
  signal memory_space_2_lc_data : std_logic_vector(159 downto 0);
  signal memory_space_2_lc_tag :  std_logic_vector(14 downto 0);
  signal memory_space_2_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(6 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(20 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(2 downto 0);
  -- interface signals to connect to memory space memory_space_3
  signal memory_space_3_lr_req :  std_logic_vector(5 downto 0);
  signal memory_space_3_lr_ack : std_logic_vector(5 downto 0);
  signal memory_space_3_lr_addr : std_logic_vector(41 downto 0);
  signal memory_space_3_lr_tag : std_logic_vector(125 downto 0);
  signal memory_space_3_lc_req : std_logic_vector(5 downto 0);
  signal memory_space_3_lc_ack :  std_logic_vector(5 downto 0);
  signal memory_space_3_lc_data : std_logic_vector(191 downto 0);
  signal memory_space_3_lc_tag :  std_logic_vector(17 downto 0);
  signal memory_space_3_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_3_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_3_sr_addr : std_logic_vector(6 downto 0);
  signal memory_space_3_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_3_sr_tag : std_logic_vector(20 downto 0);
  signal memory_space_3_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_3_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_3_sc_tag :  std_logic_vector(2 downto 0);
  -- interface signals to connect to memory space memory_space_4
  signal memory_space_4_lr_req :  std_logic_vector(3 downto 0);
  signal memory_space_4_lr_ack : std_logic_vector(3 downto 0);
  signal memory_space_4_lr_addr : std_logic_vector(55 downto 0);
  signal memory_space_4_lr_tag : std_logic_vector(75 downto 0);
  signal memory_space_4_lc_req : std_logic_vector(3 downto 0);
  signal memory_space_4_lc_ack :  std_logic_vector(3 downto 0);
  signal memory_space_4_lc_data : std_logic_vector(255 downto 0);
  signal memory_space_4_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_4_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_4_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_4_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_4_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_4_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_4_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_4_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_4_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_5
  signal memory_space_5_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_5_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_5_sr_addr : std_logic_vector(10 downto 0);
  signal memory_space_5_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_5_sr_tag : std_logic_vector(0 downto 0);
  signal memory_space_5_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_5_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_5_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_6
  signal memory_space_6_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_6_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_6_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_6_lr_tag : std_logic_vector(18 downto 0);
  signal memory_space_6_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_6_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_6_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_6_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_6_sr_req :  std_logic_vector(4 downto 0);
  signal memory_space_6_sr_ack : std_logic_vector(4 downto 0);
  signal memory_space_6_sr_addr : std_logic_vector(69 downto 0);
  signal memory_space_6_sr_data : std_logic_vector(319 downto 0);
  signal memory_space_6_sr_tag : std_logic_vector(94 downto 0);
  signal memory_space_6_sc_req : std_logic_vector(4 downto 0);
  signal memory_space_6_sc_ack :  std_logic_vector(4 downto 0);
  signal memory_space_6_sc_tag :  std_logic_vector(4 downto 0);
  -- interface signals to connect to memory space memory_space_7
  signal memory_space_7_lr_req :  std_logic_vector(3 downto 0);
  signal memory_space_7_lr_ack : std_logic_vector(3 downto 0);
  signal memory_space_7_lr_addr : std_logic_vector(3 downto 0);
  signal memory_space_7_lr_tag : std_logic_vector(75 downto 0);
  signal memory_space_7_lc_req : std_logic_vector(3 downto 0);
  signal memory_space_7_lc_ack :  std_logic_vector(3 downto 0);
  signal memory_space_7_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_7_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_7_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_7_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_7_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_7_sr_data : std_logic_vector(7 downto 0);
  signal memory_space_7_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_7_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_7_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_7_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_8
  signal memory_space_8_lr_req :  std_logic_vector(3 downto 0);
  signal memory_space_8_lr_ack : std_logic_vector(3 downto 0);
  signal memory_space_8_lr_addr : std_logic_vector(3 downto 0);
  signal memory_space_8_lr_tag : std_logic_vector(79 downto 0);
  signal memory_space_8_lc_req : std_logic_vector(3 downto 0);
  signal memory_space_8_lc_ack :  std_logic_vector(3 downto 0);
  signal memory_space_8_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_8_lc_tag :  std_logic_vector(7 downto 0);
  signal memory_space_8_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_8_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_8_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_8_sr_data : std_logic_vector(7 downto 0);
  signal memory_space_8_sr_tag : std_logic_vector(19 downto 0);
  signal memory_space_8_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_8_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_8_sc_tag :  std_logic_vector(1 downto 0);
  -- declarations related to module convTranspose
  component convTranspose is -- 
    generic (tag_length : integer); 
    port ( -- 
      Block0_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block0_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block0_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block1_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block1_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block1_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block2_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block2_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block2_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block3_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block3_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block3_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block1_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block1_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block1_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      Block0_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block0_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block0_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      Block3_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block3_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block3_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      Block2_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block2_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block2_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      elapsed_time_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      elapsed_time_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      elapsed_time_pipe_pipe_write_data : out  std_logic_vector(63 downto 0);
      testConfigure_call_reqs : out  std_logic_vector(0 downto 0);
      testConfigure_call_acks : in   std_logic_vector(0 downto 0);
      testConfigure_call_tag  :  out  std_logic_vector(0 downto 0);
      testConfigure_return_reqs : out  std_logic_vector(0 downto 0);
      testConfigure_return_acks : in   std_logic_vector(0 downto 0);
      testConfigure_return_data : in   std_logic_vector(15 downto 0);
      testConfigure_return_tag :  in   std_logic_vector(0 downto 0);
      sendOutput_call_reqs : out  std_logic_vector(0 downto 0);
      sendOutput_call_acks : in   std_logic_vector(0 downto 0);
      sendOutput_call_tag  :  out  std_logic_vector(0 downto 0);
      sendOutput_return_reqs : out  std_logic_vector(0 downto 0);
      sendOutput_return_acks : in   std_logic_vector(0 downto 0);
      sendOutput_return_tag :  in   std_logic_vector(0 downto 0);
      timer_call_reqs : out  std_logic_vector(0 downto 0);
      timer_call_acks : in   std_logic_vector(0 downto 0);
      timer_call_tag  :  out  std_logic_vector(1 downto 0);
      timer_return_reqs : out  std_logic_vector(0 downto 0);
      timer_return_acks : in   std_logic_vector(0 downto 0);
      timer_return_data : in   std_logic_vector(31 downto 0);
      timer_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTranspose
  signal convTranspose_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTranspose_tag_out   : std_logic_vector(1 downto 0);
  signal convTranspose_start_req : std_logic;
  signal convTranspose_start_ack : std_logic;
  signal convTranspose_fin_req   : std_logic;
  signal convTranspose_fin_ack : std_logic;
  -- declarations related to module convTransposeA
  component convTransposeA is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_7_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_8_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_8_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_8_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_8_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_8_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_8_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_4_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_4_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_6_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_6_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sc_tag :  in  std_logic_vector(0 downto 0);
      Block0_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block0_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block0_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block0_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block0_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block0_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeA
  signal convTransposeA_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeA_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeA_start_req : std_logic;
  signal convTransposeA_start_ack : std_logic;
  signal convTransposeA_fin_req   : std_logic;
  signal convTransposeA_fin_ack : std_logic;
  -- declarations related to module convTransposeB
  component convTransposeB is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_7_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_8_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_8_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_8_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_8_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_8_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_8_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_4_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_4_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_6_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_6_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sc_tag :  in  std_logic_vector(0 downto 0);
      Block1_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block1_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block1_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block1_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block1_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block1_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeB
  signal convTransposeB_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeB_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeB_start_req : std_logic;
  signal convTransposeB_start_ack : std_logic;
  signal convTransposeB_fin_req   : std_logic;
  signal convTransposeB_fin_ack : std_logic;
  -- declarations related to module convTransposeC
  component convTransposeC is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_7_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_8_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_8_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_8_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_8_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_8_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_8_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_4_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_4_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_6_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_6_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sc_tag :  in  std_logic_vector(0 downto 0);
      Block2_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block2_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block2_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block2_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block2_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block2_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeC
  signal convTransposeC_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeC_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeC_start_req : std_logic;
  signal convTransposeC_start_ack : std_logic;
  signal convTransposeC_fin_req   : std_logic;
  signal convTransposeC_fin_ack : std_logic;
  -- declarations related to module convTransposeD
  component convTransposeD is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_7_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_8_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_8_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_8_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_8_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_8_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_8_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_4_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_4_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_6_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_6_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sc_tag :  in  std_logic_vector(0 downto 0);
      Block3_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block3_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block3_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block3_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block3_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block3_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeD
  signal convTransposeD_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeD_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeD_start_req : std_logic;
  signal convTransposeD_start_ack : std_logic;
  signal convTransposeD_fin_req   : std_logic;
  signal convTransposeD_fin_ack : std_logic;
  -- declarations related to module sendOutput
  component sendOutput is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_6_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_6_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(2 downto 0);
      ConvTranspose_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module sendOutput
  signal sendOutput_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal sendOutput_tag_out   : std_logic_vector(1 downto 0);
  signal sendOutput_start_req : std_logic;
  signal sendOutput_start_ack : std_logic;
  signal sendOutput_fin_req   : std_logic;
  signal sendOutput_fin_ack : std_logic;
  -- caller side aggregated signals for module sendOutput
  signal sendOutput_call_reqs: std_logic_vector(0 downto 0);
  signal sendOutput_call_acks: std_logic_vector(0 downto 0);
  signal sendOutput_return_reqs: std_logic_vector(0 downto 0);
  signal sendOutput_return_acks: std_logic_vector(0 downto 0);
  signal sendOutput_call_tag: std_logic_vector(0 downto 0);
  signal sendOutput_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module testConfigure
  component testConfigure is -- 
    generic (tag_length : integer); 
    port ( -- 
      ret_val_x_x : out  std_logic_vector(15 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sr_addr : out  std_logic_vector(10 downto 0);
      memory_space_5_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_5_sr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_6_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_6_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_7_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_7_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_7_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_8_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_8_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_8_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_8_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_8_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_8_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_8_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_4_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_4_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sc_tag :  in  std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module testConfigure
  signal testConfigure_ret_val_x_x :  std_logic_vector(15 downto 0);
  signal testConfigure_out_args   : std_logic_vector(15 downto 0);
  signal testConfigure_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal testConfigure_tag_out   : std_logic_vector(1 downto 0);
  signal testConfigure_start_req : std_logic;
  signal testConfigure_start_ack : std_logic;
  signal testConfigure_fin_req   : std_logic;
  signal testConfigure_fin_ack : std_logic;
  -- caller side aggregated signals for module testConfigure
  signal testConfigure_call_reqs: std_logic_vector(0 downto 0);
  signal testConfigure_call_acks: std_logic_vector(0 downto 0);
  signal testConfigure_return_reqs: std_logic_vector(0 downto 0);
  signal testConfigure_return_acks: std_logic_vector(0 downto 0);
  signal testConfigure_call_tag: std_logic_vector(0 downto 0);
  signal testConfigure_return_data: std_logic_vector(15 downto 0);
  signal testConfigure_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module timer
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      c : out  std_logic_vector(31 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timer
  signal timer_c :  std_logic_vector(31 downto 0);
  signal timer_out_args   : std_logic_vector(31 downto 0);
  signal timer_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal timer_tag_out   : std_logic_vector(2 downto 0);
  signal timer_start_req : std_logic;
  signal timer_start_ack : std_logic;
  signal timer_fin_req   : std_logic;
  signal timer_fin_ack : std_logic;
  -- caller side aggregated signals for module timer
  signal timer_call_reqs: std_logic_vector(0 downto 0);
  signal timer_call_acks: std_logic_vector(0 downto 0);
  signal timer_return_reqs: std_logic_vector(0 downto 0);
  signal timer_return_acks: std_logic_vector(0 downto 0);
  signal timer_call_tag: std_logic_vector(1 downto 0);
  signal timer_return_data: std_logic_vector(31 downto 0);
  signal timer_return_tag: std_logic_vector(1 downto 0);
  -- aggregate signals for write to pipe Block0_done
  signal Block0_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block0_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block0_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block0_done
  signal Block0_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block0_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block0_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block0_start
  signal Block0_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block0_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block0_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block0_start
  signal Block0_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block0_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block0_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block1_done
  signal Block1_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block1_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block1_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block1_done
  signal Block1_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block1_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block1_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block1_start
  signal Block1_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block1_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block1_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block1_start
  signal Block1_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block1_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block1_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block2_done
  signal Block2_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block2_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block2_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block2_done
  signal Block2_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block2_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block2_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block2_start
  signal Block2_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block2_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block2_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block2_start
  signal Block2_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block2_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block2_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block3_done
  signal Block3_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block3_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block3_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block3_done
  signal Block3_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block3_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block3_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block3_start
  signal Block3_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block3_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block3_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block3_start
  signal Block3_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block3_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block3_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe ConvTranspose_input_pipe
  signal ConvTranspose_input_pipe_pipe_read_data: std_logic_vector(7 downto 0);
  signal ConvTranspose_input_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal ConvTranspose_input_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe ConvTranspose_output_pipe
  signal ConvTranspose_output_pipe_pipe_write_data: std_logic_vector(7 downto 0);
  signal ConvTranspose_output_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal ConvTranspose_output_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe elapsed_time_pipe
  signal elapsed_time_pipe_pipe_write_data: std_logic_vector(63 downto 0);
  signal elapsed_time_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal elapsed_time_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module convTranspose
  convTranspose_instance:convTranspose-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTranspose_start_req,
      start_ack => convTranspose_start_ack,
      fin_req => convTranspose_fin_req,
      fin_ack => convTranspose_fin_ack,
      clk => clk,
      reset => reset,
      Block0_done_pipe_read_req => Block0_done_pipe_read_req(0 downto 0),
      Block0_done_pipe_read_ack => Block0_done_pipe_read_ack(0 downto 0),
      Block0_done_pipe_read_data => Block0_done_pipe_read_data(15 downto 0),
      Block1_done_pipe_read_req => Block1_done_pipe_read_req(0 downto 0),
      Block1_done_pipe_read_ack => Block1_done_pipe_read_ack(0 downto 0),
      Block1_done_pipe_read_data => Block1_done_pipe_read_data(15 downto 0),
      Block2_done_pipe_read_req => Block2_done_pipe_read_req(0 downto 0),
      Block2_done_pipe_read_ack => Block2_done_pipe_read_ack(0 downto 0),
      Block2_done_pipe_read_data => Block2_done_pipe_read_data(15 downto 0),
      Block3_done_pipe_read_req => Block3_done_pipe_read_req(0 downto 0),
      Block3_done_pipe_read_ack => Block3_done_pipe_read_ack(0 downto 0),
      Block3_done_pipe_read_data => Block3_done_pipe_read_data(15 downto 0),
      Block1_start_pipe_write_req => Block1_start_pipe_write_req(0 downto 0),
      Block1_start_pipe_write_ack => Block1_start_pipe_write_ack(0 downto 0),
      Block1_start_pipe_write_data => Block1_start_pipe_write_data(15 downto 0),
      Block0_start_pipe_write_req => Block0_start_pipe_write_req(0 downto 0),
      Block0_start_pipe_write_ack => Block0_start_pipe_write_ack(0 downto 0),
      Block0_start_pipe_write_data => Block0_start_pipe_write_data(15 downto 0),
      Block3_start_pipe_write_req => Block3_start_pipe_write_req(0 downto 0),
      Block3_start_pipe_write_ack => Block3_start_pipe_write_ack(0 downto 0),
      Block3_start_pipe_write_data => Block3_start_pipe_write_data(15 downto 0),
      Block2_start_pipe_write_req => Block2_start_pipe_write_req(0 downto 0),
      Block2_start_pipe_write_ack => Block2_start_pipe_write_ack(0 downto 0),
      Block2_start_pipe_write_data => Block2_start_pipe_write_data(15 downto 0),
      elapsed_time_pipe_pipe_write_req => elapsed_time_pipe_pipe_write_req(0 downto 0),
      elapsed_time_pipe_pipe_write_ack => elapsed_time_pipe_pipe_write_ack(0 downto 0),
      elapsed_time_pipe_pipe_write_data => elapsed_time_pipe_pipe_write_data(63 downto 0),
      testConfigure_call_reqs => testConfigure_call_reqs(0 downto 0),
      testConfigure_call_acks => testConfigure_call_acks(0 downto 0),
      testConfigure_call_tag => testConfigure_call_tag(0 downto 0),
      testConfigure_return_reqs => testConfigure_return_reqs(0 downto 0),
      testConfigure_return_acks => testConfigure_return_acks(0 downto 0),
      testConfigure_return_data => testConfigure_return_data(15 downto 0),
      testConfigure_return_tag => testConfigure_return_tag(0 downto 0),
      timer_call_reqs => timer_call_reqs(0 downto 0),
      timer_call_acks => timer_call_acks(0 downto 0),
      timer_call_tag => timer_call_tag(1 downto 0),
      timer_return_reqs => timer_return_reqs(0 downto 0),
      timer_return_acks => timer_return_acks(0 downto 0),
      timer_return_data => timer_return_data(31 downto 0),
      timer_return_tag => timer_return_tag(1 downto 0),
      sendOutput_call_reqs => sendOutput_call_reqs(0 downto 0),
      sendOutput_call_acks => sendOutput_call_acks(0 downto 0),
      sendOutput_call_tag => sendOutput_call_tag(0 downto 0),
      sendOutput_return_reqs => sendOutput_return_reqs(0 downto 0),
      sendOutput_return_acks => sendOutput_return_acks(0 downto 0),
      sendOutput_return_tag => sendOutput_return_tag(0 downto 0),
      tag_in => convTranspose_tag_in,
      tag_out => convTranspose_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTranspose_tag_in <= (others => '0');
  convTranspose_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTranspose_start_req, start_ack => convTranspose_start_ack,  fin_req => convTranspose_fin_req,  fin_ack => convTranspose_fin_ack);
  -- module convTransposeA
  convTransposeA_instance:convTransposeA-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeA_start_req,
      start_ack => convTransposeA_start_ack,
      fin_req => convTransposeA_fin_req,
      fin_ack => convTransposeA_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(3 downto 3),
      memory_space_1_lr_ack => memory_space_1_lr_ack(3 downto 3),
      memory_space_1_lr_addr => memory_space_1_lr_addr(27 downto 21),
      memory_space_1_lr_tag => memory_space_1_lr_tag(79 downto 60),
      memory_space_1_lc_req => memory_space_1_lc_req(3 downto 3),
      memory_space_1_lc_ack => memory_space_1_lc_ack(3 downto 3),
      memory_space_1_lc_data => memory_space_1_lc_data(127 downto 96),
      memory_space_1_lc_tag => memory_space_1_lc_tag(7 downto 6),
      memory_space_2_lr_req => memory_space_2_lr_req(3 downto 3),
      memory_space_2_lr_ack => memory_space_2_lr_ack(3 downto 3),
      memory_space_2_lr_addr => memory_space_2_lr_addr(27 downto 21),
      memory_space_2_lr_tag => memory_space_2_lr_tag(83 downto 63),
      memory_space_2_lc_req => memory_space_2_lc_req(3 downto 3),
      memory_space_2_lc_ack => memory_space_2_lc_ack(3 downto 3),
      memory_space_2_lc_data => memory_space_2_lc_data(127 downto 96),
      memory_space_2_lc_tag => memory_space_2_lc_tag(11 downto 9),
      memory_space_3_lr_req => memory_space_3_lr_req(3 downto 3),
      memory_space_3_lr_ack => memory_space_3_lr_ack(3 downto 3),
      memory_space_3_lr_addr => memory_space_3_lr_addr(27 downto 21),
      memory_space_3_lr_tag => memory_space_3_lr_tag(83 downto 63),
      memory_space_3_lc_req => memory_space_3_lc_req(3 downto 3),
      memory_space_3_lc_ack => memory_space_3_lc_ack(3 downto 3),
      memory_space_3_lc_data => memory_space_3_lc_data(127 downto 96),
      memory_space_3_lc_tag => memory_space_3_lc_tag(11 downto 9),
      memory_space_4_lr_req => memory_space_4_lr_req(3 downto 3),
      memory_space_4_lr_ack => memory_space_4_lr_ack(3 downto 3),
      memory_space_4_lr_addr => memory_space_4_lr_addr(55 downto 42),
      memory_space_4_lr_tag => memory_space_4_lr_tag(75 downto 57),
      memory_space_4_lc_req => memory_space_4_lc_req(3 downto 3),
      memory_space_4_lc_ack => memory_space_4_lc_ack(3 downto 3),
      memory_space_4_lc_data => memory_space_4_lc_data(255 downto 192),
      memory_space_4_lc_tag => memory_space_4_lc_tag(3 downto 3),
      memory_space_7_lr_req => memory_space_7_lr_req(3 downto 3),
      memory_space_7_lr_ack => memory_space_7_lr_ack(3 downto 3),
      memory_space_7_lr_addr => memory_space_7_lr_addr(3 downto 3),
      memory_space_7_lr_tag => memory_space_7_lr_tag(75 downto 57),
      memory_space_7_lc_req => memory_space_7_lc_req(3 downto 3),
      memory_space_7_lc_ack => memory_space_7_lc_ack(3 downto 3),
      memory_space_7_lc_data => memory_space_7_lc_data(31 downto 24),
      memory_space_7_lc_tag => memory_space_7_lc_tag(3 downto 3),
      memory_space_8_lr_req => memory_space_8_lr_req(3 downto 3),
      memory_space_8_lr_ack => memory_space_8_lr_ack(3 downto 3),
      memory_space_8_lr_addr => memory_space_8_lr_addr(3 downto 3),
      memory_space_8_lr_tag => memory_space_8_lr_tag(79 downto 60),
      memory_space_8_lc_req => memory_space_8_lc_req(3 downto 3),
      memory_space_8_lc_ack => memory_space_8_lc_ack(3 downto 3),
      memory_space_8_lc_data => memory_space_8_lc_data(31 downto 24),
      memory_space_8_lc_tag => memory_space_8_lc_tag(7 downto 6),
      memory_space_6_sr_req => memory_space_6_sr_req(3 downto 3),
      memory_space_6_sr_ack => memory_space_6_sr_ack(3 downto 3),
      memory_space_6_sr_addr => memory_space_6_sr_addr(55 downto 42),
      memory_space_6_sr_data => memory_space_6_sr_data(255 downto 192),
      memory_space_6_sr_tag => memory_space_6_sr_tag(75 downto 57),
      memory_space_6_sc_req => memory_space_6_sc_req(3 downto 3),
      memory_space_6_sc_ack => memory_space_6_sc_ack(3 downto 3),
      memory_space_6_sc_tag => memory_space_6_sc_tag(3 downto 3),
      Block0_start_pipe_read_req => Block0_start_pipe_read_req(0 downto 0),
      Block0_start_pipe_read_ack => Block0_start_pipe_read_ack(0 downto 0),
      Block0_start_pipe_read_data => Block0_start_pipe_read_data(15 downto 0),
      Block0_done_pipe_write_req => Block0_done_pipe_write_req(0 downto 0),
      Block0_done_pipe_write_ack => Block0_done_pipe_write_ack(0 downto 0),
      Block0_done_pipe_write_data => Block0_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeA_tag_in,
      tag_out => convTransposeA_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeA_tag_in <= (others => '0');
  convTransposeA_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeA_start_req, start_ack => convTransposeA_start_ack,  fin_req => convTransposeA_fin_req,  fin_ack => convTransposeA_fin_ack);
  -- module convTransposeB
  convTransposeB_instance:convTransposeB-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeB_start_req,
      start_ack => convTransposeB_start_ack,
      fin_req => convTransposeB_fin_req,
      fin_ack => convTransposeB_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(2 downto 2),
      memory_space_1_lr_ack => memory_space_1_lr_ack(2 downto 2),
      memory_space_1_lr_addr => memory_space_1_lr_addr(20 downto 14),
      memory_space_1_lr_tag => memory_space_1_lr_tag(59 downto 40),
      memory_space_1_lc_req => memory_space_1_lc_req(2 downto 2),
      memory_space_1_lc_ack => memory_space_1_lc_ack(2 downto 2),
      memory_space_1_lc_data => memory_space_1_lc_data(95 downto 64),
      memory_space_1_lc_tag => memory_space_1_lc_tag(5 downto 4),
      memory_space_2_lr_req => memory_space_2_lr_req(2 downto 2),
      memory_space_2_lr_ack => memory_space_2_lr_ack(2 downto 2),
      memory_space_2_lr_addr => memory_space_2_lr_addr(20 downto 14),
      memory_space_2_lr_tag => memory_space_2_lr_tag(62 downto 42),
      memory_space_2_lc_req => memory_space_2_lc_req(2 downto 2),
      memory_space_2_lc_ack => memory_space_2_lc_ack(2 downto 2),
      memory_space_2_lc_data => memory_space_2_lc_data(95 downto 64),
      memory_space_2_lc_tag => memory_space_2_lc_tag(8 downto 6),
      memory_space_3_lr_req => memory_space_3_lr_req(2 downto 2),
      memory_space_3_lr_ack => memory_space_3_lr_ack(2 downto 2),
      memory_space_3_lr_addr => memory_space_3_lr_addr(20 downto 14),
      memory_space_3_lr_tag => memory_space_3_lr_tag(62 downto 42),
      memory_space_3_lc_req => memory_space_3_lc_req(2 downto 2),
      memory_space_3_lc_ack => memory_space_3_lc_ack(2 downto 2),
      memory_space_3_lc_data => memory_space_3_lc_data(95 downto 64),
      memory_space_3_lc_tag => memory_space_3_lc_tag(8 downto 6),
      memory_space_4_lr_req => memory_space_4_lr_req(2 downto 2),
      memory_space_4_lr_ack => memory_space_4_lr_ack(2 downto 2),
      memory_space_4_lr_addr => memory_space_4_lr_addr(41 downto 28),
      memory_space_4_lr_tag => memory_space_4_lr_tag(56 downto 38),
      memory_space_4_lc_req => memory_space_4_lc_req(2 downto 2),
      memory_space_4_lc_ack => memory_space_4_lc_ack(2 downto 2),
      memory_space_4_lc_data => memory_space_4_lc_data(191 downto 128),
      memory_space_4_lc_tag => memory_space_4_lc_tag(2 downto 2),
      memory_space_7_lr_req => memory_space_7_lr_req(2 downto 2),
      memory_space_7_lr_ack => memory_space_7_lr_ack(2 downto 2),
      memory_space_7_lr_addr => memory_space_7_lr_addr(2 downto 2),
      memory_space_7_lr_tag => memory_space_7_lr_tag(56 downto 38),
      memory_space_7_lc_req => memory_space_7_lc_req(2 downto 2),
      memory_space_7_lc_ack => memory_space_7_lc_ack(2 downto 2),
      memory_space_7_lc_data => memory_space_7_lc_data(23 downto 16),
      memory_space_7_lc_tag => memory_space_7_lc_tag(2 downto 2),
      memory_space_8_lr_req => memory_space_8_lr_req(2 downto 2),
      memory_space_8_lr_ack => memory_space_8_lr_ack(2 downto 2),
      memory_space_8_lr_addr => memory_space_8_lr_addr(2 downto 2),
      memory_space_8_lr_tag => memory_space_8_lr_tag(59 downto 40),
      memory_space_8_lc_req => memory_space_8_lc_req(2 downto 2),
      memory_space_8_lc_ack => memory_space_8_lc_ack(2 downto 2),
      memory_space_8_lc_data => memory_space_8_lc_data(23 downto 16),
      memory_space_8_lc_tag => memory_space_8_lc_tag(5 downto 4),
      memory_space_6_sr_req => memory_space_6_sr_req(2 downto 2),
      memory_space_6_sr_ack => memory_space_6_sr_ack(2 downto 2),
      memory_space_6_sr_addr => memory_space_6_sr_addr(41 downto 28),
      memory_space_6_sr_data => memory_space_6_sr_data(191 downto 128),
      memory_space_6_sr_tag => memory_space_6_sr_tag(56 downto 38),
      memory_space_6_sc_req => memory_space_6_sc_req(2 downto 2),
      memory_space_6_sc_ack => memory_space_6_sc_ack(2 downto 2),
      memory_space_6_sc_tag => memory_space_6_sc_tag(2 downto 2),
      Block1_start_pipe_read_req => Block1_start_pipe_read_req(0 downto 0),
      Block1_start_pipe_read_ack => Block1_start_pipe_read_ack(0 downto 0),
      Block1_start_pipe_read_data => Block1_start_pipe_read_data(15 downto 0),
      Block1_done_pipe_write_req => Block1_done_pipe_write_req(0 downto 0),
      Block1_done_pipe_write_ack => Block1_done_pipe_write_ack(0 downto 0),
      Block1_done_pipe_write_data => Block1_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeB_tag_in,
      tag_out => convTransposeB_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeB_tag_in <= (others => '0');
  convTransposeB_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeB_start_req, start_ack => convTransposeB_start_ack,  fin_req => convTransposeB_fin_req,  fin_ack => convTransposeB_fin_ack);
  -- module convTransposeC
  convTransposeC_instance:convTransposeC-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeC_start_req,
      start_ack => convTransposeC_start_ack,
      fin_req => convTransposeC_fin_req,
      fin_ack => convTransposeC_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(1 downto 1),
      memory_space_1_lr_ack => memory_space_1_lr_ack(1 downto 1),
      memory_space_1_lr_addr => memory_space_1_lr_addr(13 downto 7),
      memory_space_1_lr_tag => memory_space_1_lr_tag(39 downto 20),
      memory_space_1_lc_req => memory_space_1_lc_req(1 downto 1),
      memory_space_1_lc_ack => memory_space_1_lc_ack(1 downto 1),
      memory_space_1_lc_data => memory_space_1_lc_data(63 downto 32),
      memory_space_1_lc_tag => memory_space_1_lc_tag(3 downto 2),
      memory_space_2_lr_req => memory_space_2_lr_req(1 downto 1),
      memory_space_2_lr_ack => memory_space_2_lr_ack(1 downto 1),
      memory_space_2_lr_addr => memory_space_2_lr_addr(13 downto 7),
      memory_space_2_lr_tag => memory_space_2_lr_tag(41 downto 21),
      memory_space_2_lc_req => memory_space_2_lc_req(1 downto 1),
      memory_space_2_lc_ack => memory_space_2_lc_ack(1 downto 1),
      memory_space_2_lc_data => memory_space_2_lc_data(63 downto 32),
      memory_space_2_lc_tag => memory_space_2_lc_tag(5 downto 3),
      memory_space_3_lr_req => memory_space_3_lr_req(1 downto 1),
      memory_space_3_lr_ack => memory_space_3_lr_ack(1 downto 1),
      memory_space_3_lr_addr => memory_space_3_lr_addr(13 downto 7),
      memory_space_3_lr_tag => memory_space_3_lr_tag(41 downto 21),
      memory_space_3_lc_req => memory_space_3_lc_req(1 downto 1),
      memory_space_3_lc_ack => memory_space_3_lc_ack(1 downto 1),
      memory_space_3_lc_data => memory_space_3_lc_data(63 downto 32),
      memory_space_3_lc_tag => memory_space_3_lc_tag(5 downto 3),
      memory_space_4_lr_req => memory_space_4_lr_req(1 downto 1),
      memory_space_4_lr_ack => memory_space_4_lr_ack(1 downto 1),
      memory_space_4_lr_addr => memory_space_4_lr_addr(27 downto 14),
      memory_space_4_lr_tag => memory_space_4_lr_tag(37 downto 19),
      memory_space_4_lc_req => memory_space_4_lc_req(1 downto 1),
      memory_space_4_lc_ack => memory_space_4_lc_ack(1 downto 1),
      memory_space_4_lc_data => memory_space_4_lc_data(127 downto 64),
      memory_space_4_lc_tag => memory_space_4_lc_tag(1 downto 1),
      memory_space_7_lr_req => memory_space_7_lr_req(1 downto 1),
      memory_space_7_lr_ack => memory_space_7_lr_ack(1 downto 1),
      memory_space_7_lr_addr => memory_space_7_lr_addr(1 downto 1),
      memory_space_7_lr_tag => memory_space_7_lr_tag(37 downto 19),
      memory_space_7_lc_req => memory_space_7_lc_req(1 downto 1),
      memory_space_7_lc_ack => memory_space_7_lc_ack(1 downto 1),
      memory_space_7_lc_data => memory_space_7_lc_data(15 downto 8),
      memory_space_7_lc_tag => memory_space_7_lc_tag(1 downto 1),
      memory_space_8_lr_req => memory_space_8_lr_req(1 downto 1),
      memory_space_8_lr_ack => memory_space_8_lr_ack(1 downto 1),
      memory_space_8_lr_addr => memory_space_8_lr_addr(1 downto 1),
      memory_space_8_lr_tag => memory_space_8_lr_tag(39 downto 20),
      memory_space_8_lc_req => memory_space_8_lc_req(1 downto 1),
      memory_space_8_lc_ack => memory_space_8_lc_ack(1 downto 1),
      memory_space_8_lc_data => memory_space_8_lc_data(15 downto 8),
      memory_space_8_lc_tag => memory_space_8_lc_tag(3 downto 2),
      memory_space_6_sr_req => memory_space_6_sr_req(1 downto 1),
      memory_space_6_sr_ack => memory_space_6_sr_ack(1 downto 1),
      memory_space_6_sr_addr => memory_space_6_sr_addr(27 downto 14),
      memory_space_6_sr_data => memory_space_6_sr_data(127 downto 64),
      memory_space_6_sr_tag => memory_space_6_sr_tag(37 downto 19),
      memory_space_6_sc_req => memory_space_6_sc_req(1 downto 1),
      memory_space_6_sc_ack => memory_space_6_sc_ack(1 downto 1),
      memory_space_6_sc_tag => memory_space_6_sc_tag(1 downto 1),
      Block2_start_pipe_read_req => Block2_start_pipe_read_req(0 downto 0),
      Block2_start_pipe_read_ack => Block2_start_pipe_read_ack(0 downto 0),
      Block2_start_pipe_read_data => Block2_start_pipe_read_data(15 downto 0),
      Block2_done_pipe_write_req => Block2_done_pipe_write_req(0 downto 0),
      Block2_done_pipe_write_ack => Block2_done_pipe_write_ack(0 downto 0),
      Block2_done_pipe_write_data => Block2_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeC_tag_in,
      tag_out => convTransposeC_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeC_tag_in <= (others => '0');
  convTransposeC_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeC_start_req, start_ack => convTransposeC_start_ack,  fin_req => convTransposeC_fin_req,  fin_ack => convTransposeC_fin_ack);
  -- module convTransposeD
  convTransposeD_instance:convTransposeD-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeD_start_req,
      start_ack => convTransposeD_start_ack,
      fin_req => convTransposeD_fin_req,
      fin_ack => convTransposeD_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(6 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(19 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(31 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(1 downto 0),
      memory_space_2_lr_req => memory_space_2_lr_req(0 downto 0),
      memory_space_2_lr_ack => memory_space_2_lr_ack(0 downto 0),
      memory_space_2_lr_addr => memory_space_2_lr_addr(6 downto 0),
      memory_space_2_lr_tag => memory_space_2_lr_tag(20 downto 0),
      memory_space_2_lc_req => memory_space_2_lc_req(0 downto 0),
      memory_space_2_lc_ack => memory_space_2_lc_ack(0 downto 0),
      memory_space_2_lc_data => memory_space_2_lc_data(31 downto 0),
      memory_space_2_lc_tag => memory_space_2_lc_tag(2 downto 0),
      memory_space_3_lr_req => memory_space_3_lr_req(0 downto 0),
      memory_space_3_lr_ack => memory_space_3_lr_ack(0 downto 0),
      memory_space_3_lr_addr => memory_space_3_lr_addr(6 downto 0),
      memory_space_3_lr_tag => memory_space_3_lr_tag(20 downto 0),
      memory_space_3_lc_req => memory_space_3_lc_req(0 downto 0),
      memory_space_3_lc_ack => memory_space_3_lc_ack(0 downto 0),
      memory_space_3_lc_data => memory_space_3_lc_data(31 downto 0),
      memory_space_3_lc_tag => memory_space_3_lc_tag(2 downto 0),
      memory_space_4_lr_req => memory_space_4_lr_req(0 downto 0),
      memory_space_4_lr_ack => memory_space_4_lr_ack(0 downto 0),
      memory_space_4_lr_addr => memory_space_4_lr_addr(13 downto 0),
      memory_space_4_lr_tag => memory_space_4_lr_tag(18 downto 0),
      memory_space_4_lc_req => memory_space_4_lc_req(0 downto 0),
      memory_space_4_lc_ack => memory_space_4_lc_ack(0 downto 0),
      memory_space_4_lc_data => memory_space_4_lc_data(63 downto 0),
      memory_space_4_lc_tag => memory_space_4_lc_tag(0 downto 0),
      memory_space_7_lr_req => memory_space_7_lr_req(0 downto 0),
      memory_space_7_lr_ack => memory_space_7_lr_ack(0 downto 0),
      memory_space_7_lr_addr => memory_space_7_lr_addr(0 downto 0),
      memory_space_7_lr_tag => memory_space_7_lr_tag(18 downto 0),
      memory_space_7_lc_req => memory_space_7_lc_req(0 downto 0),
      memory_space_7_lc_ack => memory_space_7_lc_ack(0 downto 0),
      memory_space_7_lc_data => memory_space_7_lc_data(7 downto 0),
      memory_space_7_lc_tag => memory_space_7_lc_tag(0 downto 0),
      memory_space_8_lr_req => memory_space_8_lr_req(0 downto 0),
      memory_space_8_lr_ack => memory_space_8_lr_ack(0 downto 0),
      memory_space_8_lr_addr => memory_space_8_lr_addr(0 downto 0),
      memory_space_8_lr_tag => memory_space_8_lr_tag(19 downto 0),
      memory_space_8_lc_req => memory_space_8_lc_req(0 downto 0),
      memory_space_8_lc_ack => memory_space_8_lc_ack(0 downto 0),
      memory_space_8_lc_data => memory_space_8_lc_data(7 downto 0),
      memory_space_8_lc_tag => memory_space_8_lc_tag(1 downto 0),
      memory_space_6_sr_req => memory_space_6_sr_req(0 downto 0),
      memory_space_6_sr_ack => memory_space_6_sr_ack(0 downto 0),
      memory_space_6_sr_addr => memory_space_6_sr_addr(13 downto 0),
      memory_space_6_sr_data => memory_space_6_sr_data(63 downto 0),
      memory_space_6_sr_tag => memory_space_6_sr_tag(18 downto 0),
      memory_space_6_sc_req => memory_space_6_sc_req(0 downto 0),
      memory_space_6_sc_ack => memory_space_6_sc_ack(0 downto 0),
      memory_space_6_sc_tag => memory_space_6_sc_tag(0 downto 0),
      Block3_start_pipe_read_req => Block3_start_pipe_read_req(0 downto 0),
      Block3_start_pipe_read_ack => Block3_start_pipe_read_ack(0 downto 0),
      Block3_start_pipe_read_data => Block3_start_pipe_read_data(15 downto 0),
      Block3_done_pipe_write_req => Block3_done_pipe_write_req(0 downto 0),
      Block3_done_pipe_write_ack => Block3_done_pipe_write_ack(0 downto 0),
      Block3_done_pipe_write_data => Block3_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeD_tag_in,
      tag_out => convTransposeD_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeD_tag_in <= (others => '0');
  convTransposeD_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeD_start_req, start_ack => convTransposeD_start_ack,  fin_req => convTransposeD_fin_req,  fin_ack => convTransposeD_fin_ack);
  -- module sendOutput
  -- call arbiter for module sendOutput
  sendOutput_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargsNoOutargs", num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => sendOutput_call_reqs,
      call_acks => sendOutput_call_acks,
      return_reqs => sendOutput_return_reqs,
      return_acks => sendOutput_return_acks,
      call_tag  => sendOutput_call_tag,
      return_tag  => sendOutput_return_tag,
      call_mtag => sendOutput_tag_in,
      return_mtag => sendOutput_tag_out,
      call_mreq => sendOutput_start_req,
      call_mack => sendOutput_start_ack,
      return_mreq => sendOutput_fin_req,
      return_mack => sendOutput_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  sendOutput_instance:sendOutput-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => sendOutput_start_req,
      start_ack => sendOutput_start_ack,
      fin_req => sendOutput_fin_req,
      fin_ack => sendOutput_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_3_lr_req => memory_space_3_lr_req(4 downto 4),
      memory_space_3_lr_ack => memory_space_3_lr_ack(4 downto 4),
      memory_space_3_lr_addr => memory_space_3_lr_addr(34 downto 28),
      memory_space_3_lr_tag => memory_space_3_lr_tag(104 downto 84),
      memory_space_3_lc_req => memory_space_3_lc_req(4 downto 4),
      memory_space_3_lc_ack => memory_space_3_lc_ack(4 downto 4),
      memory_space_3_lc_data => memory_space_3_lc_data(159 downto 128),
      memory_space_3_lc_tag => memory_space_3_lc_tag(14 downto 12),
      memory_space_6_lr_req => memory_space_6_lr_req(0 downto 0),
      memory_space_6_lr_ack => memory_space_6_lr_ack(0 downto 0),
      memory_space_6_lr_addr => memory_space_6_lr_addr(13 downto 0),
      memory_space_6_lr_tag => memory_space_6_lr_tag(18 downto 0),
      memory_space_6_lc_req => memory_space_6_lc_req(0 downto 0),
      memory_space_6_lc_ack => memory_space_6_lc_ack(0 downto 0),
      memory_space_6_lc_data => memory_space_6_lc_data(63 downto 0),
      memory_space_6_lc_tag => memory_space_6_lc_tag(0 downto 0),
      ConvTranspose_output_pipe_pipe_write_req => ConvTranspose_output_pipe_pipe_write_req(0 downto 0),
      ConvTranspose_output_pipe_pipe_write_ack => ConvTranspose_output_pipe_pipe_write_ack(0 downto 0),
      ConvTranspose_output_pipe_pipe_write_data => ConvTranspose_output_pipe_pipe_write_data(7 downto 0),
      tag_in => sendOutput_tag_in,
      tag_out => sendOutput_tag_out-- 
    ); -- 
  -- module testConfigure
  testConfigure_out_args <= testConfigure_ret_val_x_x ;
  -- call arbiter for module testConfigure
  testConfigure_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargs", num_reqs => 1,
      return_data_width => 16,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => testConfigure_call_reqs,
      call_acks => testConfigure_call_acks,
      return_reqs => testConfigure_return_reqs,
      return_acks => testConfigure_return_acks,
      call_tag  => testConfigure_call_tag,
      return_tag  => testConfigure_return_tag,
      call_mtag => testConfigure_tag_in,
      return_mtag => testConfigure_tag_out,
      return_data =>testConfigure_return_data,
      call_mreq => testConfigure_start_req,
      call_mack => testConfigure_start_ack,
      return_mreq => testConfigure_fin_req,
      return_mack => testConfigure_fin_ack,
      return_mdata => testConfigure_out_args,
      clk => clk, 
      reset => reset --
    ); --
  testConfigure_instance:testConfigure-- 
    generic map(tag_length => 2)
    port map(-- 
      ret_val_x_x => testConfigure_ret_val_x_x,
      start_req => testConfigure_start_req,
      start_ack => testConfigure_start_ack,
      fin_req => testConfigure_fin_req,
      fin_ack => testConfigure_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(4 downto 4),
      memory_space_1_lr_ack => memory_space_1_lr_ack(4 downto 4),
      memory_space_1_lr_addr => memory_space_1_lr_addr(34 downto 28),
      memory_space_1_lr_tag => memory_space_1_lr_tag(99 downto 80),
      memory_space_1_lc_req => memory_space_1_lc_req(4 downto 4),
      memory_space_1_lc_ack => memory_space_1_lc_ack(4 downto 4),
      memory_space_1_lc_data => memory_space_1_lc_data(159 downto 128),
      memory_space_1_lc_tag => memory_space_1_lc_tag(9 downto 8),
      memory_space_2_lr_req => memory_space_2_lr_req(4 downto 4),
      memory_space_2_lr_ack => memory_space_2_lr_ack(4 downto 4),
      memory_space_2_lr_addr => memory_space_2_lr_addr(34 downto 28),
      memory_space_2_lr_tag => memory_space_2_lr_tag(104 downto 84),
      memory_space_2_lc_req => memory_space_2_lc_req(4 downto 4),
      memory_space_2_lc_ack => memory_space_2_lc_ack(4 downto 4),
      memory_space_2_lc_data => memory_space_2_lc_data(159 downto 128),
      memory_space_2_lc_tag => memory_space_2_lc_tag(14 downto 12),
      memory_space_3_lr_req => memory_space_3_lr_req(5 downto 5),
      memory_space_3_lr_ack => memory_space_3_lr_ack(5 downto 5),
      memory_space_3_lr_addr => memory_space_3_lr_addr(41 downto 35),
      memory_space_3_lr_tag => memory_space_3_lr_tag(125 downto 105),
      memory_space_3_lc_req => memory_space_3_lc_req(5 downto 5),
      memory_space_3_lc_ack => memory_space_3_lc_ack(5 downto 5),
      memory_space_3_lc_data => memory_space_3_lc_data(191 downto 160),
      memory_space_3_lc_tag => memory_space_3_lc_tag(17 downto 15),
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(6 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(31 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(19 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(1 downto 0),
      memory_space_2_sr_req => memory_space_2_sr_req(0 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(0 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(6 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(31 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(20 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(0 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(0 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(2 downto 0),
      memory_space_3_sr_req => memory_space_3_sr_req(0 downto 0),
      memory_space_3_sr_ack => memory_space_3_sr_ack(0 downto 0),
      memory_space_3_sr_addr => memory_space_3_sr_addr(6 downto 0),
      memory_space_3_sr_data => memory_space_3_sr_data(31 downto 0),
      memory_space_3_sr_tag => memory_space_3_sr_tag(20 downto 0),
      memory_space_3_sc_req => memory_space_3_sc_req(0 downto 0),
      memory_space_3_sc_ack => memory_space_3_sc_ack(0 downto 0),
      memory_space_3_sc_tag => memory_space_3_sc_tag(2 downto 0),
      memory_space_4_sr_req => memory_space_4_sr_req(0 downto 0),
      memory_space_4_sr_ack => memory_space_4_sr_ack(0 downto 0),
      memory_space_4_sr_addr => memory_space_4_sr_addr(13 downto 0),
      memory_space_4_sr_data => memory_space_4_sr_data(63 downto 0),
      memory_space_4_sr_tag => memory_space_4_sr_tag(18 downto 0),
      memory_space_4_sc_req => memory_space_4_sc_req(0 downto 0),
      memory_space_4_sc_ack => memory_space_4_sc_ack(0 downto 0),
      memory_space_4_sc_tag => memory_space_4_sc_tag(0 downto 0),
      memory_space_5_sr_req => memory_space_5_sr_req(0 downto 0),
      memory_space_5_sr_ack => memory_space_5_sr_ack(0 downto 0),
      memory_space_5_sr_addr => memory_space_5_sr_addr(10 downto 0),
      memory_space_5_sr_data => memory_space_5_sr_data(63 downto 0),
      memory_space_5_sr_tag => memory_space_5_sr_tag(0 downto 0),
      memory_space_5_sc_req => memory_space_5_sc_req(0 downto 0),
      memory_space_5_sc_ack => memory_space_5_sc_ack(0 downto 0),
      memory_space_5_sc_tag => memory_space_5_sc_tag(0 downto 0),
      memory_space_6_sr_req => memory_space_6_sr_req(4 downto 4),
      memory_space_6_sr_ack => memory_space_6_sr_ack(4 downto 4),
      memory_space_6_sr_addr => memory_space_6_sr_addr(69 downto 56),
      memory_space_6_sr_data => memory_space_6_sr_data(319 downto 256),
      memory_space_6_sr_tag => memory_space_6_sr_tag(94 downto 76),
      memory_space_6_sc_req => memory_space_6_sc_req(4 downto 4),
      memory_space_6_sc_ack => memory_space_6_sc_ack(4 downto 4),
      memory_space_6_sc_tag => memory_space_6_sc_tag(4 downto 4),
      memory_space_7_sr_req => memory_space_7_sr_req(0 downto 0),
      memory_space_7_sr_ack => memory_space_7_sr_ack(0 downto 0),
      memory_space_7_sr_addr => memory_space_7_sr_addr(0 downto 0),
      memory_space_7_sr_data => memory_space_7_sr_data(7 downto 0),
      memory_space_7_sr_tag => memory_space_7_sr_tag(18 downto 0),
      memory_space_7_sc_req => memory_space_7_sc_req(0 downto 0),
      memory_space_7_sc_ack => memory_space_7_sc_ack(0 downto 0),
      memory_space_7_sc_tag => memory_space_7_sc_tag(0 downto 0),
      memory_space_8_sr_req => memory_space_8_sr_req(0 downto 0),
      memory_space_8_sr_ack => memory_space_8_sr_ack(0 downto 0),
      memory_space_8_sr_addr => memory_space_8_sr_addr(0 downto 0),
      memory_space_8_sr_data => memory_space_8_sr_data(7 downto 0),
      memory_space_8_sr_tag => memory_space_8_sr_tag(19 downto 0),
      memory_space_8_sc_req => memory_space_8_sc_req(0 downto 0),
      memory_space_8_sc_ack => memory_space_8_sc_ack(0 downto 0),
      memory_space_8_sc_tag => memory_space_8_sc_tag(1 downto 0),
      ConvTranspose_input_pipe_pipe_read_req => ConvTranspose_input_pipe_pipe_read_req(0 downto 0),
      ConvTranspose_input_pipe_pipe_read_ack => ConvTranspose_input_pipe_pipe_read_ack(0 downto 0),
      ConvTranspose_input_pipe_pipe_read_data => ConvTranspose_input_pipe_pipe_read_data(7 downto 0),
      tag_in => testConfigure_tag_in,
      tag_out => testConfigure_tag_out-- 
    ); -- 
  -- module timer
  timer_out_args <= timer_c ;
  -- call arbiter for module timer
  timer_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargs", num_reqs => 1,
      return_data_width => 32,
      callee_tag_length => 1,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => timer_call_reqs,
      call_acks => timer_call_acks,
      return_reqs => timer_return_reqs,
      return_acks => timer_return_acks,
      call_tag  => timer_call_tag,
      return_tag  => timer_return_tag,
      call_mtag => timer_tag_in,
      return_mtag => timer_tag_out,
      return_data =>timer_return_data,
      call_mreq => timer_start_req,
      call_mack => timer_start_ack,
      return_mreq => timer_fin_req,
      return_mack => timer_fin_ack,
      return_mdata => timer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  timer_instance:timer-- 
    generic map(tag_length => 3)
    port map(-- 
      c => timer_c,
      start_req => timer_start_req,
      start_ack => timer_start_ack,
      fin_req => timer_fin_req,
      fin_ack => timer_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(0 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(0 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(31 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(0 downto 0),
      tag_in => timer_tag_in,
      tag_out => timer_tag_out-- 
    ); -- 
  Block0_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block0_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block0_done_pipe_read_req,
      read_ack => Block0_done_pipe_read_ack,
      read_data => Block0_done_pipe_read_data,
      write_req => Block0_done_pipe_write_req,
      write_ack => Block0_done_pipe_write_ack,
      write_data => Block0_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block0_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block0_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block0_start_pipe_read_req,
      read_ack => Block0_start_pipe_read_ack,
      read_data => Block0_start_pipe_read_data,
      write_req => Block0_start_pipe_write_req,
      write_ack => Block0_start_pipe_write_ack,
      write_data => Block0_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block1_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block1_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block1_done_pipe_read_req,
      read_ack => Block1_done_pipe_read_ack,
      read_data => Block1_done_pipe_read_data,
      write_req => Block1_done_pipe_write_req,
      write_ack => Block1_done_pipe_write_ack,
      write_data => Block1_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block1_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block1_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block1_start_pipe_read_req,
      read_ack => Block1_start_pipe_read_ack,
      read_data => Block1_start_pipe_read_data,
      write_req => Block1_start_pipe_write_req,
      write_ack => Block1_start_pipe_write_ack,
      write_data => Block1_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block2_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block2_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block2_done_pipe_read_req,
      read_ack => Block2_done_pipe_read_ack,
      read_data => Block2_done_pipe_read_data,
      write_req => Block2_done_pipe_write_req,
      write_ack => Block2_done_pipe_write_ack,
      write_data => Block2_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block2_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block2_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block2_start_pipe_read_req,
      read_ack => Block2_start_pipe_read_ack,
      read_data => Block2_start_pipe_read_data,
      write_req => Block2_start_pipe_write_req,
      write_ack => Block2_start_pipe_write_ack,
      write_data => Block2_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block3_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block3_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block3_done_pipe_read_req,
      read_ack => Block3_done_pipe_read_ack,
      read_data => Block3_done_pipe_read_data,
      write_req => Block3_done_pipe_write_req,
      write_ack => Block3_done_pipe_write_ack,
      write_data => Block3_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block3_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block3_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block3_start_pipe_read_req,
      read_ack => Block3_start_pipe_read_ack,
      read_data => Block3_start_pipe_read_data,
      write_req => Block3_start_pipe_write_req,
      write_ack => Block3_start_pipe_write_ack,
      write_data => Block3_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  ConvTranspose_input_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe ConvTranspose_input_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => ConvTranspose_input_pipe_pipe_read_req,
      read_ack => ConvTranspose_input_pipe_pipe_read_ack,
      read_data => ConvTranspose_input_pipe_pipe_read_data,
      write_req => ConvTranspose_input_pipe_pipe_write_req,
      write_ack => ConvTranspose_input_pipe_pipe_write_ack,
      write_data => ConvTranspose_input_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  ConvTranspose_output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe ConvTranspose_output_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => ConvTranspose_output_pipe_pipe_read_req,
      read_ack => ConvTranspose_output_pipe_pipe_read_ack,
      read_data => ConvTranspose_output_pipe_pipe_read_data,
      write_req => ConvTranspose_output_pipe_pipe_write_req,
      write_ack => ConvTranspose_output_pipe_pipe_write_ack,
      write_data => ConvTranspose_output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  elapsed_time_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe elapsed_time_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => elapsed_time_pipe_pipe_read_req,
      read_ack => elapsed_time_pipe_pipe_read_ack,
      read_data => elapsed_time_pipe_pipe_read_data,
      write_req => elapsed_time_pipe_pipe_write_req,
      write_ack => elapsed_time_pipe_pipe_write_ack,
      write_data => elapsed_time_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  dummyROM_memory_space_0: dummy_read_only_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 1,
      addr_width => 1,
      data_width => 32,
      tag_width => 1
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_1: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_loads => 5,
      num_stores => 1,
      addr_width => 7,
      data_width => 32,
      tag_width => 2,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 7,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_2: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_2",
      num_loads => 5,
      num_stores => 1,
      addr_width => 7,
      data_width => 32,
      tag_width => 3,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 7,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_2_lr_addr,
      lr_req_in => memory_space_2_lr_req,
      lr_ack_out => memory_space_2_lr_ack,
      lr_tag_in => memory_space_2_lr_tag,
      lc_req_in => memory_space_2_lc_req,
      lc_ack_out => memory_space_2_lc_ack,
      lc_data_out => memory_space_2_lc_data,
      lc_tag_out => memory_space_2_lc_tag,
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_3: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_3",
      num_loads => 6,
      num_stores => 1,
      addr_width => 7,
      data_width => 32,
      tag_width => 3,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 7,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_3_lr_addr,
      lr_req_in => memory_space_3_lr_req,
      lr_ack_out => memory_space_3_lr_ack,
      lr_tag_in => memory_space_3_lr_tag,
      lc_req_in => memory_space_3_lc_req,
      lc_ack_out => memory_space_3_lc_ack,
      lc_data_out => memory_space_3_lc_data,
      lc_tag_out => memory_space_3_lc_tag,
      sr_addr_in => memory_space_3_sr_addr,
      sr_data_in => memory_space_3_sr_data,
      sr_req_in => memory_space_3_sr_req,
      sr_ack_out => memory_space_3_sr_ack,
      sr_tag_in => memory_space_3_sr_tag,
      sc_req_in=> memory_space_3_sc_req,
      sc_ack_out => memory_space_3_sc_ack,
      sc_tag_out => memory_space_3_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_4: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_4",
      num_loads => 4,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_4_lr_addr,
      lr_req_in => memory_space_4_lr_req,
      lr_ack_out => memory_space_4_lr_ack,
      lr_tag_in => memory_space_4_lr_tag,
      lc_req_in => memory_space_4_lc_req,
      lc_ack_out => memory_space_4_lc_ack,
      lc_data_out => memory_space_4_lc_data,
      lc_tag_out => memory_space_4_lc_tag,
      sr_addr_in => memory_space_4_sr_addr,
      sr_data_in => memory_space_4_sr_data,
      sr_req_in => memory_space_4_sr_req,
      sr_ack_out => memory_space_4_sr_ack,
      sr_tag_in => memory_space_4_sr_tag,
      sc_req_in=> memory_space_4_sc_req,
      sc_ack_out => memory_space_4_sc_ack,
      sc_tag_out => memory_space_4_sc_tag,
      clock => clk,
      reset => reset); -- 
  dummyWOM_memory_space_5: dummy_write_only_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_5",
      num_stores => 1,
      addr_width => 11,
      data_width => 64,
      tag_width => 1
      ) -- 
    port map(-- 
      sr_addr_in => memory_space_5_sr_addr,
      sr_data_in => memory_space_5_sr_data,
      sr_req_in => memory_space_5_sr_req,
      sr_ack_out => memory_space_5_sr_ack,
      sr_tag_in => memory_space_5_sr_tag,
      sc_req_in=> memory_space_5_sc_req,
      sc_ack_out => memory_space_5_sc_ack,
      sc_tag_out => memory_space_5_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_6: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_6",
      num_loads => 1,
      num_stores => 5,
      addr_width => 14,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_6_lr_addr,
      lr_req_in => memory_space_6_lr_req,
      lr_ack_out => memory_space_6_lr_ack,
      lr_tag_in => memory_space_6_lr_tag,
      lc_req_in => memory_space_6_lc_req,
      lc_ack_out => memory_space_6_lc_ack,
      lc_data_out => memory_space_6_lc_data,
      lc_tag_out => memory_space_6_lc_tag,
      sr_addr_in => memory_space_6_sr_addr,
      sr_data_in => memory_space_6_sr_data,
      sr_req_in => memory_space_6_sr_req,
      sr_ack_out => memory_space_6_sr_ack,
      sr_tag_in => memory_space_6_sr_tag,
      sc_req_in=> memory_space_6_sc_req,
      sc_ack_out => memory_space_6_sc_ack,
      sc_tag_out => memory_space_6_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_7: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_7",
      num_loads => 4,
      num_stores => 1,
      addr_width => 1,
      data_width => 8,
      tag_width => 1,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 8
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_7_lr_addr,
      lr_req_in => memory_space_7_lr_req,
      lr_ack_out => memory_space_7_lr_ack,
      lr_tag_in => memory_space_7_lr_tag,
      lc_req_in => memory_space_7_lc_req,
      lc_ack_out => memory_space_7_lc_ack,
      lc_data_out => memory_space_7_lc_data,
      lc_tag_out => memory_space_7_lc_tag,
      sr_addr_in => memory_space_7_sr_addr,
      sr_data_in => memory_space_7_sr_data,
      sr_req_in => memory_space_7_sr_req,
      sr_ack_out => memory_space_7_sr_ack,
      sr_tag_in => memory_space_7_sr_tag,
      sc_req_in=> memory_space_7_sc_req,
      sc_ack_out => memory_space_7_sc_ack,
      sc_tag_out => memory_space_7_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_8: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_8",
      num_loads => 4,
      num_stores => 1,
      addr_width => 1,
      data_width => 8,
      tag_width => 2,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 8
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_8_lr_addr,
      lr_req_in => memory_space_8_lr_req,
      lr_ack_out => memory_space_8_lr_ack,
      lr_tag_in => memory_space_8_lr_tag,
      lc_req_in => memory_space_8_lc_req,
      lc_ack_out => memory_space_8_lc_ack,
      lc_data_out => memory_space_8_lc_data,
      lc_tag_out => memory_space_8_lc_tag,
      sr_addr_in => memory_space_8_sr_addr,
      sr_data_in => memory_space_8_sr_data,
      sr_req_in => memory_space_8_sr_req,
      sr_ack_out => memory_space_8_sr_ack,
      sr_tag_in => memory_space_8_sr_tag,
      sc_req_in=> memory_space_8_sc_req,
      sc_ack_out => memory_space_8_sc_ack,
      sc_tag_out => memory_space_8_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
