-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity access_T is -- 
  generic (tag_length : integer); 
  port ( -- 
    num_cont : in  std_logic_vector(15 downto 0);
    row1 : in  std_logic_vector(15 downto 0);
    col1 : in  std_logic_vector(15 downto 0);
    rk1 : in  std_logic_vector(15 downto 0);
    chl_in : in  std_logic_vector(15 downto 0);
    ct : in  std_logic_vector(15 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
    input_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
    input_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
    input_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity access_T;
architecture access_T_arch of access_T is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 96)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal num_cont_buffer :  std_logic_vector(15 downto 0);
  signal num_cont_update_enable: Boolean;
  signal row1_buffer :  std_logic_vector(15 downto 0);
  signal row1_update_enable: Boolean;
  signal col1_buffer :  std_logic_vector(15 downto 0);
  signal col1_update_enable: Boolean;
  signal rk1_buffer :  std_logic_vector(15 downto 0);
  signal rk1_update_enable: Boolean;
  signal chl_in_buffer :  std_logic_vector(15 downto 0);
  signal chl_in_update_enable: Boolean;
  signal ct_buffer :  std_logic_vector(15 downto 0);
  signal ct_update_enable: Boolean;
  -- output port buffer signals
  signal access_T_CP_0_start: Boolean;
  signal access_T_CP_0_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal do_while_stmt_44_branch_req_0 : boolean;
  signal phi_stmt_46_ack_0 : boolean;
  signal phi_stmt_46_req_1 : boolean;
  signal phi_stmt_46_req_0 : boolean;
  signal n_address_280_50_buf_req_0 : boolean;
  signal n_address_280_50_buf_ack_0 : boolean;
  signal n_address_280_50_buf_req_1 : boolean;
  signal n_address_280_50_buf_ack_1 : boolean;
  signal phi_stmt_51_req_1 : boolean;
  signal phi_stmt_51_req_0 : boolean;
  signal phi_stmt_51_ack_0 : boolean;
  signal n_word_start_269_56_buf_req_0 : boolean;
  signal n_word_start_269_56_buf_ack_0 : boolean;
  signal n_word_start_269_56_buf_req_1 : boolean;
  signal n_word_start_269_56_buf_ack_1 : boolean;
  signal n_winr_209_68_buf_req_1 : boolean;
  signal n_winr_209_68_buf_ack_1 : boolean;
  signal phi_stmt_57_req_1 : boolean;
  signal phi_stmt_57_req_0 : boolean;
  signal phi_stmt_57_ack_0 : boolean;
  signal nl_start_35_59_buf_req_0 : boolean;
  signal nl_start_35_59_buf_ack_0 : boolean;
  signal nl_start_35_59_buf_req_1 : boolean;
  signal nl_start_35_59_buf_ack_1 : boolean;
  signal n_left_288_60_buf_req_0 : boolean;
  signal n_left_288_60_buf_ack_0 : boolean;
  signal n_left_288_60_buf_req_1 : boolean;
  signal n_left_288_60_buf_ack_1 : boolean;
  signal phi_stmt_61_req_1 : boolean;
  signal phi_stmt_61_req_0 : boolean;
  signal phi_stmt_61_ack_0 : boolean;
  signal type_cast_64_inst_req_0 : boolean;
  signal type_cast_64_inst_ack_0 : boolean;
  signal type_cast_64_inst_req_1 : boolean;
  signal type_cast_64_inst_ack_1 : boolean;
  signal n_blk_308_65_buf_req_0 : boolean;
  signal n_blk_308_65_buf_ack_0 : boolean;
  signal n_blk_308_65_buf_req_1 : boolean;
  signal n_blk_308_65_buf_ack_1 : boolean;
  signal phi_stmt_66_req_0 : boolean;
  signal phi_stmt_66_req_1 : boolean;
  signal phi_stmt_66_ack_0 : boolean;
  signal n_winr_209_68_buf_req_0 : boolean;
  signal n_winr_209_68_buf_ack_0 : boolean;
  signal WPIPE_input_pipe1_167_inst_ack_0 : boolean;
  signal WPIPE_input_pipe1_167_inst_req_1 : boolean;
  signal WPIPE_input_pipe1_167_inst_ack_1 : boolean;
  signal W_c3_164_delayed_14_0_170_inst_req_0 : boolean;
  signal W_c3_164_delayed_14_0_170_inst_ack_0 : boolean;
  signal W_c3_164_delayed_14_0_170_inst_req_1 : boolean;
  signal W_c3_164_delayed_14_0_170_inst_ack_1 : boolean;
  signal phi_stmt_71_req_0 : boolean;
  signal phi_stmt_71_req_1 : boolean;
  signal phi_stmt_71_ack_0 : boolean;
  signal n_col_222_73_buf_req_0 : boolean;
  signal n_col_222_73_buf_ack_0 : boolean;
  signal n_col_222_73_buf_req_1 : boolean;
  signal n_col_222_73_buf_ack_1 : boolean;
  signal phi_stmt_76_req_1 : boolean;
  signal phi_stmt_76_req_0 : boolean;
  signal phi_stmt_76_ack_0 : boolean;
  signal n_row_234_80_buf_req_0 : boolean;
  signal n_row_234_80_buf_ack_0 : boolean;
  signal n_row_234_80_buf_req_1 : boolean;
  signal n_row_234_80_buf_ack_1 : boolean;
  signal array_obj_ref_133_index_offset_req_0 : boolean;
  signal array_obj_ref_133_index_offset_ack_0 : boolean;
  signal array_obj_ref_133_index_offset_req_1 : boolean;
  signal array_obj_ref_133_index_offset_ack_1 : boolean;
  signal addr_of_134_final_reg_req_0 : boolean;
  signal addr_of_134_final_reg_ack_0 : boolean;
  signal addr_of_134_final_reg_req_1 : boolean;
  signal addr_of_134_final_reg_ack_1 : boolean;
  signal ptr_deref_138_load_0_req_0 : boolean;
  signal ptr_deref_138_load_0_ack_0 : boolean;
  signal ptr_deref_138_load_0_req_1 : boolean;
  signal ptr_deref_138_load_0_ack_1 : boolean;
  signal slice_142_inst_req_0 : boolean;
  signal slice_142_inst_ack_0 : boolean;
  signal slice_142_inst_req_1 : boolean;
  signal slice_142_inst_ack_1 : boolean;
  signal slice_146_inst_req_0 : boolean;
  signal slice_146_inst_ack_0 : boolean;
  signal slice_146_inst_req_1 : boolean;
  signal slice_146_inst_ack_1 : boolean;
  signal slice_150_inst_req_0 : boolean;
  signal slice_150_inst_ack_0 : boolean;
  signal slice_150_inst_req_1 : boolean;
  signal slice_150_inst_ack_1 : boolean;
  signal slice_154_inst_req_0 : boolean;
  signal slice_154_inst_ack_0 : boolean;
  signal slice_154_inst_req_1 : boolean;
  signal slice_154_inst_ack_1 : boolean;
  signal W_c1_156_delayed_14_0_156_inst_req_0 : boolean;
  signal W_c1_156_delayed_14_0_156_inst_ack_0 : boolean;
  signal W_c1_156_delayed_14_0_156_inst_req_1 : boolean;
  signal W_c1_156_delayed_14_0_156_inst_ack_1 : boolean;
  signal WPIPE_input_pipe1_160_inst_req_0 : boolean;
  signal WPIPE_input_pipe1_160_inst_ack_0 : boolean;
  signal WPIPE_input_pipe1_160_inst_req_1 : boolean;
  signal WPIPE_input_pipe1_160_inst_ack_1 : boolean;
  signal W_c2_160_delayed_14_0_163_inst_req_0 : boolean;
  signal W_c2_160_delayed_14_0_163_inst_ack_0 : boolean;
  signal W_c2_160_delayed_14_0_163_inst_req_1 : boolean;
  signal W_c2_160_delayed_14_0_163_inst_ack_1 : boolean;
  signal WPIPE_input_pipe1_167_inst_req_0 : boolean;
  signal WPIPE_input_pipe1_174_inst_req_0 : boolean;
  signal WPIPE_input_pipe1_174_inst_ack_0 : boolean;
  signal WPIPE_input_pipe1_174_inst_req_1 : boolean;
  signal WPIPE_input_pipe1_174_inst_ack_1 : boolean;
  signal W_c4_168_delayed_14_0_177_inst_req_0 : boolean;
  signal W_c4_168_delayed_14_0_177_inst_ack_0 : boolean;
  signal W_c4_168_delayed_14_0_177_inst_req_1 : boolean;
  signal W_c4_168_delayed_14_0_177_inst_ack_1 : boolean;
  signal WPIPE_input_pipe1_181_inst_req_0 : boolean;
  signal WPIPE_input_pipe1_181_inst_ack_0 : boolean;
  signal WPIPE_input_pipe1_181_inst_req_1 : boolean;
  signal WPIPE_input_pipe1_181_inst_ack_1 : boolean;
  signal do_while_stmt_44_branch_ack_0 : boolean;
  signal do_while_stmt_44_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "access_T_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 96) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(15 downto 0) <= num_cont;
  num_cont_buffer <= in_buffer_data_out(15 downto 0);
  in_buffer_data_in(31 downto 16) <= row1;
  row1_buffer <= in_buffer_data_out(31 downto 16);
  in_buffer_data_in(47 downto 32) <= col1;
  col1_buffer <= in_buffer_data_out(47 downto 32);
  in_buffer_data_in(63 downto 48) <= rk1;
  rk1_buffer <= in_buffer_data_out(63 downto 48);
  in_buffer_data_in(79 downto 64) <= chl_in;
  chl_in_buffer <= in_buffer_data_out(79 downto 64);
  in_buffer_data_in(95 downto 80) <= ct;
  ct_buffer <= in_buffer_data_out(95 downto 80);
  in_buffer_data_in(tag_length + 95 downto 96) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 95 downto 96);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  access_T_CP_0_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "access_T_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= access_T_CP_0_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= access_T_CP_0_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= access_T_CP_0_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  access_T_CP_0: Block -- control-path 
    signal access_T_CP_0_elements: BooleanArray(207 downto 0);
    -- 
  begin -- 
    access_T_CP_0_elements(0) <= access_T_CP_0_start;
    access_T_CP_0_symbol <= access_T_CP_0_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_32_to_assign_stmt_43__exit__
      -- CP-element group 0: 	 branch_block_stmt_26/do_while_stmt_44__entry__
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_26/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/branch_block_stmt_26__entry__
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_32_to_assign_stmt_43__entry__
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_32_to_assign_stmt_43/$entry
      -- CP-element group 0: 	 branch_block_stmt_26/assign_stmt_32_to_assign_stmt_43/$exit
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	207 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_26/$exit
      -- CP-element group 1: 	 branch_block_stmt_26/branch_block_stmt_26__exit__
      -- CP-element group 1: 	 branch_block_stmt_26/do_while_stmt_44__exit__
      -- 
    access_T_CP_0_elements(1) <= access_T_CP_0_elements(207);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_26/do_while_stmt_44/$entry
      -- CP-element group 2: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44__entry__
      -- 
    access_T_CP_0_elements(2) <= access_T_CP_0_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	207 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44__exit__
      -- 
    -- Element group access_T_CP_0_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_26/do_while_stmt_44/loop_back
      -- 
    -- Element group access_T_CP_0_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	205 
    -- CP-element group 5: 	206 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_26/do_while_stmt_44/condition_done
      -- CP-element group 5: 	 branch_block_stmt_26/do_while_stmt_44/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_26/do_while_stmt_44/loop_taken/$entry
      -- 
    access_T_CP_0_elements(5) <= access_T_CP_0_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	204 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_26/do_while_stmt_44/loop_body_done
      -- 
    access_T_CP_0_elements(6) <= access_T_CP_0_elements(204);
    -- CP-element group 7:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	116 
    -- CP-element group 7: 	97 
    -- CP-element group 7: 	76 
    -- CP-element group 7: 	135 
    -- CP-element group 7: 	21 
    -- CP-element group 7: 	40 
    -- CP-element group 7: 	59 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/back_edge_to_loop_body
      -- 
    access_T_CP_0_elements(7) <= access_T_CP_0_elements(4);
    -- CP-element group 8:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	99 
    -- CP-element group 8: 	78 
    -- CP-element group 8: 	118 
    -- CP-element group 8: 	137 
    -- CP-element group 8: 	23 
    -- CP-element group 8: 	42 
    -- CP-element group 8: 	61 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/first_time_through_loop_body
      -- 
    access_T_CP_0_elements(8) <= access_T_CP_0_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	149 
    -- CP-element group 9: 	203 
    -- CP-element group 9: 	92 
    -- CP-element group 9: 	110 
    -- CP-element group 9: 	111 
    -- CP-element group 9: 	129 
    -- CP-element group 9: 	73 
    -- CP-element group 9: 	72 
    -- CP-element group 9: 	91 
    -- CP-element group 9: 	130 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	34 
    -- CP-element group 9: 	35 
    -- CP-element group 9: 	150 
    -- CP-element group 9: 	53 
    -- CP-element group 9: 	54 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/loop_body_start
      -- 
    -- Element group access_T_CP_0_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	203 
    -- CP-element group 10: 	14 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/condition_evaluated
      -- 
    condition_evaluated_29_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_29_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(10), ack => do_while_stmt_44_branch_req_0); -- 
    access_T_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(203) & access_T_CP_0_elements(14);
      gj_access_T_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	110 
    -- CP-element group 11: 	129 
    -- CP-element group 11: 	72 
    -- CP-element group 11: 	91 
    -- CP-element group 11: 	15 
    -- CP-element group 11: 	34 
    -- CP-element group 11: 	53 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	112 
    -- CP-element group 11: 	93 
    -- CP-element group 11: 	131 
    -- CP-element group 11: 	17 
    -- CP-element group 11: 	36 
    -- CP-element group 11: 	55 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_61_sample_start__ps
      -- 
    access_T_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= access_T_CP_0_elements(110) & access_T_CP_0_elements(129) & access_T_CP_0_elements(72) & access_T_CP_0_elements(91) & access_T_CP_0_elements(15) & access_T_CP_0_elements(34) & access_T_CP_0_elements(53) & access_T_CP_0_elements(14);
      gj_access_T_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	74 
    -- CP-element group 12: 	94 
    -- CP-element group 12: 	132 
    -- CP-element group 12: 	113 
    -- CP-element group 12: 	18 
    -- CP-element group 12: 	37 
    -- CP-element group 12: 	56 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	204 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	110 
    -- CP-element group 12: 	129 
    -- CP-element group 12: 	72 
    -- CP-element group 12: 	91 
    -- CP-element group 12: 	15 
    -- CP-element group 12: 	34 
    -- CP-element group 12: 	53 
    -- CP-element group 12:  members (8) 
      -- CP-element group 12: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_51_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_57_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_61_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_66_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_71_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_76_sample_completed_
      -- 
    access_T_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= access_T_CP_0_elements(74) & access_T_CP_0_elements(94) & access_T_CP_0_elements(132) & access_T_CP_0_elements(113) & access_T_CP_0_elements(18) & access_T_CP_0_elements(37) & access_T_CP_0_elements(56);
      gj_access_T_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	92 
    -- CP-element group 13: 	111 
    -- CP-element group 13: 	73 
    -- CP-element group 13: 	130 
    -- CP-element group 13: 	16 
    -- CP-element group 13: 	35 
    -- CP-element group 13: 	54 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	114 
    -- CP-element group 13: 	95 
    -- CP-element group 13: 	133 
    -- CP-element group 13: 	19 
    -- CP-element group 13: 	38 
    -- CP-element group 13: 	57 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_61_update_start__ps
      -- 
    access_T_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= access_T_CP_0_elements(92) & access_T_CP_0_elements(111) & access_T_CP_0_elements(73) & access_T_CP_0_elements(130) & access_T_CP_0_elements(16) & access_T_CP_0_elements(35) & access_T_CP_0_elements(54);
      gj_access_T_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	115 
    -- CP-element group 14: 	96 
    -- CP-element group 14: 	134 
    -- CP-element group 14: 	75 
    -- CP-element group 14: 	20 
    -- CP-element group 14: 	39 
    -- CP-element group 14: 	58 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/aggregated_phi_update_ack
      -- 
    access_T_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= access_T_CP_0_elements(115) & access_T_CP_0_elements(96) & access_T_CP_0_elements(134) & access_T_CP_0_elements(75) & access_T_CP_0_elements(20) & access_T_CP_0_elements(39) & access_T_CP_0_elements(58);
      gj_access_T_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_sample_start_
      -- 
    access_T_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	151 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_update_start_
      -- 
    access_T_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(151);
      gj_access_T_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	11 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_sample_start__ps
      -- 
    access_T_CP_0_elements(17) <= access_T_CP_0_elements(11);
    -- CP-element group 18:  join  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	12 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	13 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_update_start__ps
      -- 
    access_T_CP_0_elements(19) <= access_T_CP_0_elements(13);
    -- CP-element group 20:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	14 
    -- CP-element group 20: 	151 
    -- CP-element group 20:  members (15) 
      -- CP-element group 20: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_update_completed__ps
      -- CP-element group 20: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_index_resized_1
      -- CP-element group 20: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_index_scaled_1
      -- CP-element group 20: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_index_computed_1
      -- CP-element group 20: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_index_resize_1/$entry
      -- CP-element group 20: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_index_resize_1/$exit
      -- CP-element group 20: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_index_resize_1/index_resize_req
      -- CP-element group 20: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_index_resize_1/index_resize_ack
      -- CP-element group 20: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_index_scale_1/$entry
      -- CP-element group 20: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_index_scale_1/$exit
      -- CP-element group 20: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_index_scale_1/scale_rename_req
      -- CP-element group 20: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_index_scale_1/scale_rename_ack
      -- CP-element group 20: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_final_index_sum_regn_Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_final_index_sum_regn_Sample/req
      -- 
    req_387_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_387_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(20), ack => array_obj_ref_133_index_offset_req_0); -- 
    -- Element group access_T_CP_0_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	7 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_loopback_trigger
      -- 
    access_T_CP_0_elements(21) <= access_T_CP_0_elements(7);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_loopback_sample_req
      -- CP-element group 22: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_loopback_sample_req_ps
      -- 
    phi_stmt_46_loopback_sample_req_44_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_46_loopback_sample_req_44_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(22), ack => phi_stmt_46_req_1); -- 
    -- Element group access_T_CP_0_elements(22) is bound as output of CP function.
    -- CP-element group 23:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	8 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_entry_trigger
      -- 
    access_T_CP_0_elements(23) <= access_T_CP_0_elements(8);
    -- CP-element group 24:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (2) 
      -- CP-element group 24: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_entry_sample_req
      -- CP-element group 24: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_entry_sample_req_ps
      -- 
    phi_stmt_46_entry_sample_req_47_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_46_entry_sample_req_47_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(24), ack => phi_stmt_46_req_0); -- 
    -- Element group access_T_CP_0_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_phi_mux_ack
      -- CP-element group 25: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_46_phi_mux_ack_ps
      -- 
    phi_stmt_46_phi_mux_ack_50_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_46_ack_0, ack => access_T_CP_0_elements(25)); -- 
    -- CP-element group 26:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (4) 
      -- CP-element group 26: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_49_sample_start__ps
      -- CP-element group 26: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_49_sample_completed__ps
      -- CP-element group 26: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_49_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_49_sample_completed_
      -- 
    -- Element group access_T_CP_0_elements(26) is bound as output of CP function.
    -- CP-element group 27:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (2) 
      -- CP-element group 27: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_49_update_start__ps
      -- CP-element group 27: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_49_update_start_
      -- 
    -- Element group access_T_CP_0_elements(27) is bound as output of CP function.
    -- CP-element group 28:  join  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	29 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_49_update_completed__ps
      -- 
    access_T_CP_0_elements(28) <= access_T_CP_0_elements(29);
    -- CP-element group 29:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	28 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_49_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(29) is a control-delay.
    cp_element_29_delay: control_delay_element  generic map(name => " 29_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(27), ack => access_T_CP_0_elements(29), clk => clk, reset =>reset);
    -- CP-element group 30:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	32 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_address_50_sample_start__ps
      -- CP-element group 30: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_address_50_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_address_50_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_address_50_Sample/req
      -- 
    req_71_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_71_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(30), ack => n_address_280_50_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(30) is bound as output of CP function.
    -- CP-element group 31:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_address_50_update_start__ps
      -- CP-element group 31: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_address_50_update_start_
      -- CP-element group 31: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_address_50_Update/$entry
      -- CP-element group 31: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_address_50_Update/req
      -- 
    req_76_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_76_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(31), ack => n_address_280_50_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(31) is bound as output of CP function.
    -- CP-element group 32:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	30 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (4) 
      -- CP-element group 32: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_address_50_sample_completed__ps
      -- CP-element group 32: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_address_50_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_address_50_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_address_50_Sample/ack
      -- 
    ack_72_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address_280_50_buf_ack_0, ack => access_T_CP_0_elements(32)); -- 
    -- CP-element group 33:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (4) 
      -- CP-element group 33: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_address_50_update_completed__ps
      -- CP-element group 33: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_address_50_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_address_50_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_address_50_Update/ack
      -- 
    ack_77_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address_280_50_buf_ack_1, ack => access_T_CP_0_elements(33)); -- 
    -- CP-element group 34:  join  transition  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	9 
    -- CP-element group 34: marked-predecessors 
    -- CP-element group 34: 	12 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	11 
    -- CP-element group 34:  members (1) 
      -- CP-element group 34: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_51_sample_start_
      -- 
    access_T_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  join  transition  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	9 
    -- CP-element group 35: marked-predecessors 
    -- CP-element group 35: 	191 
    -- CP-element group 35: 	198 
    -- CP-element group 35: 	184 
    -- CP-element group 35: 	177 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	13 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_51_update_start_
      -- 
    access_T_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(191) & access_T_CP_0_elements(198) & access_T_CP_0_elements(184) & access_T_CP_0_elements(177);
      gj_access_T_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	11 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_51_sample_start__ps
      -- 
    access_T_CP_0_elements(36) <= access_T_CP_0_elements(11);
    -- CP-element group 37:  join  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	12 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_51_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(37) is bound as output of CP function.
    -- CP-element group 38:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	13 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_51_update_start__ps
      -- 
    access_T_CP_0_elements(38) <= access_T_CP_0_elements(13);
    -- CP-element group 39:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	14 
    -- CP-element group 39: 	196 
    -- CP-element group 39: 	182 
    -- CP-element group 39: 	189 
    -- CP-element group 39: 	175 
    -- CP-element group 39:  members (2) 
      -- CP-element group 39: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_51_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_51_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(39) is bound as output of CP function.
    -- CP-element group 40:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	7 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_51_loopback_trigger
      -- 
    access_T_CP_0_elements(40) <= access_T_CP_0_elements(7);
    -- CP-element group 41:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (2) 
      -- CP-element group 41: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_51_loopback_sample_req
      -- CP-element group 41: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_51_loopback_sample_req_ps
      -- 
    phi_stmt_51_loopback_sample_req_88_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_51_loopback_sample_req_88_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(41), ack => phi_stmt_51_req_1); -- 
    -- Element group access_T_CP_0_elements(41) is bound as output of CP function.
    -- CP-element group 42:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	8 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_51_entry_trigger
      -- 
    access_T_CP_0_elements(42) <= access_T_CP_0_elements(8);
    -- CP-element group 43:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (2) 
      -- CP-element group 43: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_51_entry_sample_req
      -- CP-element group 43: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_51_entry_sample_req_ps
      -- 
    phi_stmt_51_entry_sample_req_91_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_51_entry_sample_req_91_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(43), ack => phi_stmt_51_req_0); -- 
    -- Element group access_T_CP_0_elements(43) is bound as output of CP function.
    -- CP-element group 44:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_51_phi_mux_ack
      -- CP-element group 44: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_51_phi_mux_ack_ps
      -- 
    phi_stmt_51_phi_mux_ack_94_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_51_ack_0, ack => access_T_CP_0_elements(44)); -- 
    -- CP-element group 45:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (4) 
      -- CP-element group 45: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_55_sample_start__ps
      -- CP-element group 45: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_55_sample_completed__ps
      -- CP-element group 45: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_55_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_55_sample_completed_
      -- 
    -- Element group access_T_CP_0_elements(45) is bound as output of CP function.
    -- CP-element group 46:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	48 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_55_update_start__ps
      -- CP-element group 46: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_55_update_start_
      -- 
    -- Element group access_T_CP_0_elements(46) is bound as output of CP function.
    -- CP-element group 47:  join  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	48 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_55_update_completed__ps
      -- 
    access_T_CP_0_elements(47) <= access_T_CP_0_elements(48);
    -- CP-element group 48:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	46 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	47 
    -- CP-element group 48:  members (1) 
      -- CP-element group 48: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_55_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(48) is a control-delay.
    cp_element_48_delay: control_delay_element  generic map(name => " 48_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(46), ack => access_T_CP_0_elements(48), clk => clk, reset =>reset);
    -- CP-element group 49:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (4) 
      -- CP-element group 49: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_word_start_56_sample_start__ps
      -- CP-element group 49: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_word_start_56_sample_start_
      -- CP-element group 49: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_word_start_56_Sample/$entry
      -- CP-element group 49: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_word_start_56_Sample/req
      -- 
    req_115_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_115_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(49), ack => n_word_start_269_56_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(49) is bound as output of CP function.
    -- CP-element group 50:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (4) 
      -- CP-element group 50: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_word_start_56_update_start__ps
      -- CP-element group 50: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_word_start_56_update_start_
      -- CP-element group 50: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_word_start_56_Update/$entry
      -- CP-element group 50: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_word_start_56_Update/req
      -- 
    req_120_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_120_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(50), ack => n_word_start_269_56_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(50) is bound as output of CP function.
    -- CP-element group 51:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (4) 
      -- CP-element group 51: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_word_start_56_sample_completed__ps
      -- CP-element group 51: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_word_start_56_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_word_start_56_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_word_start_56_Sample/ack
      -- 
    ack_116_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_word_start_269_56_buf_ack_0, ack => access_T_CP_0_elements(51)); -- 
    -- CP-element group 52:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (4) 
      -- CP-element group 52: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_word_start_56_update_completed__ps
      -- CP-element group 52: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_word_start_56_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_word_start_56_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_word_start_56_Update/ack
      -- 
    ack_121_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_word_start_269_56_buf_ack_1, ack => access_T_CP_0_elements(52)); -- 
    -- CP-element group 53:  join  transition  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	9 
    -- CP-element group 53: marked-predecessors 
    -- CP-element group 53: 	12 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	11 
    -- CP-element group 53:  members (1) 
      -- CP-element group 53: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_57_sample_start_
      -- 
    access_T_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  join  transition  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	9 
    -- CP-element group 54: marked-predecessors 
    -- CP-element group 54: 	58 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	13 
    -- CP-element group 54:  members (1) 
      -- CP-element group 54: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_57_update_start_
      -- 
    access_T_cp_element_group_54: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_54"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(58);
      gj_access_T_cp_element_group_54 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(54), clk => clk, reset => reset); --
    end block;
    -- CP-element group 55:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	11 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (1) 
      -- CP-element group 55: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_57_sample_start__ps
      -- 
    access_T_CP_0_elements(55) <= access_T_CP_0_elements(11);
    -- CP-element group 56:  join  transition  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	12 
    -- CP-element group 56:  members (1) 
      -- CP-element group 56: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_57_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(56) is bound as output of CP function.
    -- CP-element group 57:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	13 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (1) 
      -- CP-element group 57: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_57_update_start__ps
      -- 
    access_T_CP_0_elements(57) <= access_T_CP_0_elements(13);
    -- CP-element group 58:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	14 
    -- CP-element group 58: marked-successors 
    -- CP-element group 58: 	54 
    -- CP-element group 58:  members (2) 
      -- CP-element group 58: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_57_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_57_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(58) is bound as output of CP function.
    -- CP-element group 59:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	7 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_57_loopback_trigger
      -- 
    access_T_CP_0_elements(59) <= access_T_CP_0_elements(7);
    -- CP-element group 60:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: successors 
    -- CP-element group 60:  members (2) 
      -- CP-element group 60: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_57_loopback_sample_req
      -- CP-element group 60: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_57_loopback_sample_req_ps
      -- 
    phi_stmt_57_loopback_sample_req_132_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_57_loopback_sample_req_132_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(60), ack => phi_stmt_57_req_1); -- 
    -- Element group access_T_CP_0_elements(60) is bound as output of CP function.
    -- CP-element group 61:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	8 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (1) 
      -- CP-element group 61: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_57_entry_trigger
      -- 
    access_T_CP_0_elements(61) <= access_T_CP_0_elements(8);
    -- CP-element group 62:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (2) 
      -- CP-element group 62: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_57_entry_sample_req
      -- CP-element group 62: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_57_entry_sample_req_ps
      -- 
    phi_stmt_57_entry_sample_req_135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_57_entry_sample_req_135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(62), ack => phi_stmt_57_req_0); -- 
    -- Element group access_T_CP_0_elements(62) is bound as output of CP function.
    -- CP-element group 63:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (2) 
      -- CP-element group 63: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_57_phi_mux_ack
      -- CP-element group 63: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_57_phi_mux_ack_ps
      -- 
    phi_stmt_57_phi_mux_ack_138_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_57_ack_0, ack => access_T_CP_0_elements(63)); -- 
    -- CP-element group 64:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	66 
    -- CP-element group 64:  members (4) 
      -- CP-element group 64: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_nl_start_59_sample_start__ps
      -- CP-element group 64: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_nl_start_59_sample_start_
      -- CP-element group 64: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_nl_start_59_Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_nl_start_59_Sample/req
      -- 
    req_151_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_151_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(64), ack => nl_start_35_59_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(64) is bound as output of CP function.
    -- CP-element group 65:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	67 
    -- CP-element group 65:  members (4) 
      -- CP-element group 65: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_nl_start_59_update_start__ps
      -- CP-element group 65: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_nl_start_59_update_start_
      -- CP-element group 65: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_nl_start_59_Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_nl_start_59_Update/req
      -- 
    req_156_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_156_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(65), ack => nl_start_35_59_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(65) is bound as output of CP function.
    -- CP-element group 66:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	64 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (4) 
      -- CP-element group 66: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_nl_start_59_sample_completed__ps
      -- CP-element group 66: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_nl_start_59_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_nl_start_59_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_nl_start_59_Sample/ack
      -- 
    ack_152_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nl_start_35_59_buf_ack_0, ack => access_T_CP_0_elements(66)); -- 
    -- CP-element group 67:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	65 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (4) 
      -- CP-element group 67: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_nl_start_59_update_completed__ps
      -- CP-element group 67: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_nl_start_59_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_nl_start_59_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_nl_start_59_Update/ack
      -- 
    ack_157_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nl_start_35_59_buf_ack_1, ack => access_T_CP_0_elements(67)); -- 
    -- CP-element group 68:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (4) 
      -- CP-element group 68: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_left_60_sample_start__ps
      -- CP-element group 68: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_left_60_sample_start_
      -- CP-element group 68: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_left_60_Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_left_60_Sample/req
      -- 
    req_169_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_169_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(68), ack => n_left_288_60_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(68) is bound as output of CP function.
    -- CP-element group 69:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	71 
    -- CP-element group 69:  members (4) 
      -- CP-element group 69: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_left_60_update_start__ps
      -- CP-element group 69: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_left_60_update_start_
      -- CP-element group 69: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_left_60_Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_left_60_Update/req
      -- 
    req_174_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_174_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(69), ack => n_left_288_60_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(69) is bound as output of CP function.
    -- CP-element group 70:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (4) 
      -- CP-element group 70: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_left_60_sample_completed__ps
      -- CP-element group 70: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_left_60_sample_completed_
      -- CP-element group 70: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_left_60_Sample/$exit
      -- CP-element group 70: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_left_60_Sample/ack
      -- 
    ack_170_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_left_288_60_buf_ack_0, ack => access_T_CP_0_elements(70)); -- 
    -- CP-element group 71:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	69 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (4) 
      -- CP-element group 71: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_left_60_update_completed__ps
      -- CP-element group 71: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_left_60_update_completed_
      -- CP-element group 71: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_left_60_Update/$exit
      -- CP-element group 71: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_left_60_Update/ack
      -- 
    ack_175_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_left_288_60_buf_ack_1, ack => access_T_CP_0_elements(71)); -- 
    -- CP-element group 72:  join  transition  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	9 
    -- CP-element group 72: marked-predecessors 
    -- CP-element group 72: 	12 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	11 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_61_sample_start_
      -- 
    access_T_cp_element_group_72: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_72"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_72 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(72), clk => clk, reset => reset); --
    end block;
    -- CP-element group 73:  join  transition  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	9 
    -- CP-element group 73: marked-predecessors 
    -- CP-element group 73: 	191 
    -- CP-element group 73: 	198 
    -- CP-element group 73: 	184 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	13 
    -- CP-element group 73:  members (1) 
      -- CP-element group 73: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_61_update_start_
      -- 
    access_T_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(191) & access_T_CP_0_elements(198) & access_T_CP_0_elements(184);
      gj_access_T_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  join  transition  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	12 
    -- CP-element group 74:  members (1) 
      -- CP-element group 74: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_61_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(74) is bound as output of CP function.
    -- CP-element group 75:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	14 
    -- CP-element group 75: 	196 
    -- CP-element group 75: 	182 
    -- CP-element group 75: 	189 
    -- CP-element group 75:  members (2) 
      -- CP-element group 75: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_61_update_completed_
      -- CP-element group 75: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_61_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(75) is bound as output of CP function.
    -- CP-element group 76:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	7 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (1) 
      -- CP-element group 76: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_61_loopback_trigger
      -- 
    access_T_CP_0_elements(76) <= access_T_CP_0_elements(7);
    -- CP-element group 77:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: successors 
    -- CP-element group 77:  members (2) 
      -- CP-element group 77: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_61_loopback_sample_req
      -- CP-element group 77: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_61_loopback_sample_req_ps
      -- 
    phi_stmt_61_loopback_sample_req_186_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_61_loopback_sample_req_186_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(77), ack => phi_stmt_61_req_1); -- 
    -- Element group access_T_CP_0_elements(77) is bound as output of CP function.
    -- CP-element group 78:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	8 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_61_entry_trigger
      -- 
    access_T_CP_0_elements(78) <= access_T_CP_0_elements(8);
    -- CP-element group 79:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_61_entry_sample_req
      -- CP-element group 79: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_61_entry_sample_req_ps
      -- 
    phi_stmt_61_entry_sample_req_189_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_61_entry_sample_req_189_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(79), ack => phi_stmt_61_req_0); -- 
    -- Element group access_T_CP_0_elements(79) is bound as output of CP function.
    -- CP-element group 80:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (2) 
      -- CP-element group 80: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_61_phi_mux_ack
      -- CP-element group 80: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_61_phi_mux_ack_ps
      -- 
    phi_stmt_61_phi_mux_ack_192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_61_ack_0, ack => access_T_CP_0_elements(80)); -- 
    -- CP-element group 81:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	83 
    -- CP-element group 81:  members (1) 
      -- CP-element group 81: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_64_sample_start__ps
      -- 
    -- Element group access_T_CP_0_elements(81) is bound as output of CP function.
    -- CP-element group 82:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	84 
    -- CP-element group 82:  members (1) 
      -- CP-element group 82: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_64_update_start__ps
      -- 
    -- Element group access_T_CP_0_elements(82) is bound as output of CP function.
    -- CP-element group 83:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	81 
    -- CP-element group 83: marked-predecessors 
    -- CP-element group 83: 	85 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	85 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_64_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_64_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_64_Sample/rr
      -- 
    rr_205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(83), ack => type_cast_64_inst_req_0); -- 
    access_T_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(81) & access_T_CP_0_elements(85);
      gj_access_T_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: marked-predecessors 
    -- CP-element group 84: 	86 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_64_update_start_
      -- CP-element group 84: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_64_Update/$entry
      -- CP-element group 84: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_64_Update/cr
      -- 
    cr_210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(84), ack => type_cast_64_inst_req_1); -- 
    access_T_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(82) & access_T_CP_0_elements(86);
      gj_access_T_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	83 
    -- CP-element group 85: successors 
    -- CP-element group 85: marked-successors 
    -- CP-element group 85: 	83 
    -- CP-element group 85:  members (4) 
      -- CP-element group 85: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_64_sample_completed__ps
      -- CP-element group 85: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_64_sample_completed_
      -- CP-element group 85: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_64_Sample/$exit
      -- CP-element group 85: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_64_Sample/ra
      -- 
    ra_206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_64_inst_ack_0, ack => access_T_CP_0_elements(85)); -- 
    -- CP-element group 86:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: successors 
    -- CP-element group 86: marked-successors 
    -- CP-element group 86: 	84 
    -- CP-element group 86:  members (4) 
      -- CP-element group 86: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_64_update_completed__ps
      -- CP-element group 86: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_64_update_completed_
      -- CP-element group 86: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_64_Update/$exit
      -- CP-element group 86: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_64_Update/ca
      -- 
    ca_211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_64_inst_ack_1, ack => access_T_CP_0_elements(86)); -- 
    -- CP-element group 87:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	89 
    -- CP-element group 87:  members (4) 
      -- CP-element group 87: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_blk_65_sample_start__ps
      -- CP-element group 87: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_blk_65_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_blk_65_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_blk_65_Sample/req
      -- 
    req_223_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_223_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(87), ack => n_blk_308_65_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(87) is bound as output of CP function.
    -- CP-element group 88:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	90 
    -- CP-element group 88:  members (4) 
      -- CP-element group 88: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_blk_65_update_start__ps
      -- CP-element group 88: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_blk_65_update_start_
      -- CP-element group 88: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_blk_65_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_blk_65_Update/req
      -- 
    req_228_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_228_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(88), ack => n_blk_308_65_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(88) is bound as output of CP function.
    -- CP-element group 89:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	87 
    -- CP-element group 89: successors 
    -- CP-element group 89:  members (4) 
      -- CP-element group 89: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_blk_65_sample_completed__ps
      -- CP-element group 89: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_blk_65_sample_completed_
      -- CP-element group 89: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_blk_65_Sample/$exit
      -- CP-element group 89: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_blk_65_Sample/ack
      -- 
    ack_224_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_blk_308_65_buf_ack_0, ack => access_T_CP_0_elements(89)); -- 
    -- CP-element group 90:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	88 
    -- CP-element group 90: successors 
    -- CP-element group 90:  members (4) 
      -- CP-element group 90: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_blk_65_update_completed__ps
      -- CP-element group 90: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_blk_65_update_completed_
      -- CP-element group 90: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_blk_65_Update/$exit
      -- CP-element group 90: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_blk_65_Update/ack
      -- 
    ack_229_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_blk_308_65_buf_ack_1, ack => access_T_CP_0_elements(90)); -- 
    -- CP-element group 91:  join  transition  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	9 
    -- CP-element group 91: marked-predecessors 
    -- CP-element group 91: 	12 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	11 
    -- CP-element group 91:  members (1) 
      -- CP-element group 91: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_66_sample_start_
      -- 
    access_T_cp_element_group_91: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_91"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_91 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(91), clk => clk, reset => reset); --
    end block;
    -- CP-element group 92:  join  transition  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	9 
    -- CP-element group 92: marked-predecessors 
    -- CP-element group 92: 	96 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	13 
    -- CP-element group 92:  members (1) 
      -- CP-element group 92: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_66_update_start_
      -- 
    access_T_cp_element_group_92: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_92"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(96);
      gj_access_T_cp_element_group_92 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(92), clk => clk, reset => reset); --
    end block;
    -- CP-element group 93:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	11 
    -- CP-element group 93: successors 
    -- CP-element group 93:  members (1) 
      -- CP-element group 93: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_66_sample_start__ps
      -- 
    access_T_CP_0_elements(93) <= access_T_CP_0_elements(11);
    -- CP-element group 94:  join  transition  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	12 
    -- CP-element group 94:  members (1) 
      -- CP-element group 94: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_66_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(94) is bound as output of CP function.
    -- CP-element group 95:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	13 
    -- CP-element group 95: successors 
    -- CP-element group 95:  members (1) 
      -- CP-element group 95: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_66_update_start__ps
      -- 
    access_T_CP_0_elements(95) <= access_T_CP_0_elements(13);
    -- CP-element group 96:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	14 
    -- CP-element group 96: marked-successors 
    -- CP-element group 96: 	92 
    -- CP-element group 96:  members (2) 
      -- CP-element group 96: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_66_update_completed_
      -- CP-element group 96: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_66_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(96) is bound as output of CP function.
    -- CP-element group 97:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	7 
    -- CP-element group 97: successors 
    -- CP-element group 97:  members (1) 
      -- CP-element group 97: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_66_loopback_trigger
      -- 
    access_T_CP_0_elements(97) <= access_T_CP_0_elements(7);
    -- CP-element group 98:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: successors 
    -- CP-element group 98:  members (2) 
      -- CP-element group 98: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_66_loopback_sample_req
      -- CP-element group 98: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_66_loopback_sample_req_ps
      -- 
    phi_stmt_66_loopback_sample_req_240_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_66_loopback_sample_req_240_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(98), ack => phi_stmt_66_req_0); -- 
    -- Element group access_T_CP_0_elements(98) is bound as output of CP function.
    -- CP-element group 99:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	8 
    -- CP-element group 99: successors 
    -- CP-element group 99:  members (1) 
      -- CP-element group 99: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_66_entry_trigger
      -- 
    access_T_CP_0_elements(99) <= access_T_CP_0_elements(8);
    -- CP-element group 100:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: successors 
    -- CP-element group 100:  members (2) 
      -- CP-element group 100: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_66_entry_sample_req
      -- CP-element group 100: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_66_entry_sample_req_ps
      -- 
    phi_stmt_66_entry_sample_req_243_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_66_entry_sample_req_243_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(100), ack => phi_stmt_66_req_1); -- 
    -- Element group access_T_CP_0_elements(100) is bound as output of CP function.
    -- CP-element group 101:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (2) 
      -- CP-element group 101: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_66_phi_mux_ack
      -- CP-element group 101: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_66_phi_mux_ack_ps
      -- 
    phi_stmt_66_phi_mux_ack_246_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_66_ack_0, ack => access_T_CP_0_elements(101)); -- 
    -- CP-element group 102:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	104 
    -- CP-element group 102:  members (4) 
      -- CP-element group 102: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_winr_68_sample_start__ps
      -- CP-element group 102: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_winr_68_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_winr_68_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_winr_68_Sample/req
      -- 
    req_259_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_259_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(102), ack => n_winr_209_68_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(102) is bound as output of CP function.
    -- CP-element group 103:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	105 
    -- CP-element group 103:  members (4) 
      -- CP-element group 103: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_winr_68_Update/$entry
      -- CP-element group 103: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_winr_68_Update/req
      -- CP-element group 103: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_winr_68_update_start__ps
      -- CP-element group 103: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_winr_68_update_start_
      -- 
    req_264_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_264_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(103), ack => n_winr_209_68_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(103) is bound as output of CP function.
    -- CP-element group 104:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	102 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (4) 
      -- CP-element group 104: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_winr_68_sample_completed__ps
      -- CP-element group 104: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_winr_68_sample_completed_
      -- CP-element group 104: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_winr_68_Sample/$exit
      -- CP-element group 104: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_winr_68_Sample/ack
      -- 
    ack_260_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_winr_209_68_buf_ack_0, ack => access_T_CP_0_elements(104)); -- 
    -- CP-element group 105:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	103 
    -- CP-element group 105: successors 
    -- CP-element group 105:  members (4) 
      -- CP-element group 105: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_winr_68_Update/$exit
      -- CP-element group 105: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_winr_68_Update/ack
      -- CP-element group 105: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_winr_68_update_completed__ps
      -- CP-element group 105: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_winr_68_update_completed_
      -- 
    ack_265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_winr_209_68_buf_ack_1, ack => access_T_CP_0_elements(105)); -- 
    -- CP-element group 106:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: successors 
    -- CP-element group 106:  members (4) 
      -- CP-element group 106: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_70_sample_start__ps
      -- CP-element group 106: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_70_sample_completed__ps
      -- CP-element group 106: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_70_sample_start_
      -- CP-element group 106: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_70_sample_completed_
      -- 
    -- Element group access_T_CP_0_elements(106) is bound as output of CP function.
    -- CP-element group 107:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	109 
    -- CP-element group 107:  members (2) 
      -- CP-element group 107: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_70_update_start__ps
      -- CP-element group 107: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_70_update_start_
      -- 
    -- Element group access_T_CP_0_elements(107) is bound as output of CP function.
    -- CP-element group 108:  join  transition  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	109 
    -- CP-element group 108: successors 
    -- CP-element group 108:  members (1) 
      -- CP-element group 108: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_70_update_completed__ps
      -- 
    access_T_CP_0_elements(108) <= access_T_CP_0_elements(109);
    -- CP-element group 109:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	107 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	108 
    -- CP-element group 109:  members (1) 
      -- CP-element group 109: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_70_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(109) is a control-delay.
    cp_element_109_delay: control_delay_element  generic map(name => " 109_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(107), ack => access_T_CP_0_elements(109), clk => clk, reset =>reset);
    -- CP-element group 110:  join  transition  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	9 
    -- CP-element group 110: marked-predecessors 
    -- CP-element group 110: 	12 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	11 
    -- CP-element group 110:  members (1) 
      -- CP-element group 110: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_71_sample_start_
      -- 
    access_T_cp_element_group_110: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_110"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_110 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(110), clk => clk, reset => reset); --
    end block;
    -- CP-element group 111:  join  transition  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	9 
    -- CP-element group 111: marked-predecessors 
    -- CP-element group 111: 	115 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	13 
    -- CP-element group 111:  members (1) 
      -- CP-element group 111: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_71_update_start_
      -- 
    access_T_cp_element_group_111: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_111"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(115);
      gj_access_T_cp_element_group_111 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(111), clk => clk, reset => reset); --
    end block;
    -- CP-element group 112:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	11 
    -- CP-element group 112: successors 
    -- CP-element group 112:  members (1) 
      -- CP-element group 112: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_71_sample_start__ps
      -- 
    access_T_CP_0_elements(112) <= access_T_CP_0_elements(11);
    -- CP-element group 113:  join  transition  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	12 
    -- CP-element group 113:  members (1) 
      -- CP-element group 113: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_71_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(113) is bound as output of CP function.
    -- CP-element group 114:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	13 
    -- CP-element group 114: successors 
    -- CP-element group 114:  members (1) 
      -- CP-element group 114: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_71_update_start__ps
      -- 
    access_T_CP_0_elements(114) <= access_T_CP_0_elements(13);
    -- CP-element group 115:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	14 
    -- CP-element group 115: marked-successors 
    -- CP-element group 115: 	111 
    -- CP-element group 115:  members (2) 
      -- CP-element group 115: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_71_update_completed_
      -- CP-element group 115: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_71_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(115) is bound as output of CP function.
    -- CP-element group 116:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	7 
    -- CP-element group 116: successors 
    -- CP-element group 116:  members (1) 
      -- CP-element group 116: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_71_loopback_trigger
      -- 
    access_T_CP_0_elements(116) <= access_T_CP_0_elements(7);
    -- CP-element group 117:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: successors 
    -- CP-element group 117:  members (2) 
      -- CP-element group 117: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_71_loopback_sample_req
      -- CP-element group 117: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_71_loopback_sample_req_ps
      -- 
    phi_stmt_71_loopback_sample_req_284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_71_loopback_sample_req_284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(117), ack => phi_stmt_71_req_0); -- 
    -- Element group access_T_CP_0_elements(117) is bound as output of CP function.
    -- CP-element group 118:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	8 
    -- CP-element group 118: successors 
    -- CP-element group 118:  members (1) 
      -- CP-element group 118: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_71_entry_trigger
      -- 
    access_T_CP_0_elements(118) <= access_T_CP_0_elements(8);
    -- CP-element group 119:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: successors 
    -- CP-element group 119:  members (2) 
      -- CP-element group 119: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_71_entry_sample_req
      -- CP-element group 119: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_71_entry_sample_req_ps
      -- 
    phi_stmt_71_entry_sample_req_287_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_71_entry_sample_req_287_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(119), ack => phi_stmt_71_req_1); -- 
    -- Element group access_T_CP_0_elements(119) is bound as output of CP function.
    -- CP-element group 120:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: successors 
    -- CP-element group 120:  members (2) 
      -- CP-element group 120: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_71_phi_mux_ack
      -- CP-element group 120: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_71_phi_mux_ack_ps
      -- 
    phi_stmt_71_phi_mux_ack_290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_71_ack_0, ack => access_T_CP_0_elements(120)); -- 
    -- CP-element group 121:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	123 
    -- CP-element group 121:  members (4) 
      -- CP-element group 121: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_col_73_sample_start__ps
      -- CP-element group 121: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_col_73_sample_start_
      -- CP-element group 121: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_col_73_Sample/$entry
      -- CP-element group 121: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_col_73_Sample/req
      -- 
    req_303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(121), ack => n_col_222_73_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(121) is bound as output of CP function.
    -- CP-element group 122:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	124 
    -- CP-element group 122:  members (4) 
      -- CP-element group 122: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_col_73_update_start__ps
      -- CP-element group 122: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_col_73_update_start_
      -- CP-element group 122: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_col_73_Update/$entry
      -- CP-element group 122: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_col_73_Update/req
      -- 
    req_308_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_308_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(122), ack => n_col_222_73_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(122) is bound as output of CP function.
    -- CP-element group 123:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	121 
    -- CP-element group 123: successors 
    -- CP-element group 123:  members (4) 
      -- CP-element group 123: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_col_73_sample_completed__ps
      -- CP-element group 123: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_col_73_sample_completed_
      -- CP-element group 123: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_col_73_Sample/$exit
      -- CP-element group 123: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_col_73_Sample/ack
      -- 
    ack_304_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_col_222_73_buf_ack_0, ack => access_T_CP_0_elements(123)); -- 
    -- CP-element group 124:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	122 
    -- CP-element group 124: successors 
    -- CP-element group 124:  members (4) 
      -- CP-element group 124: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_col_73_update_completed__ps
      -- CP-element group 124: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_col_73_update_completed_
      -- CP-element group 124: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_col_73_Update/$exit
      -- CP-element group 124: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_col_73_Update/ack
      -- 
    ack_309_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_col_222_73_buf_ack_1, ack => access_T_CP_0_elements(124)); -- 
    -- CP-element group 125:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: successors 
    -- CP-element group 125:  members (4) 
      -- CP-element group 125: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_75_sample_start__ps
      -- CP-element group 125: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_75_sample_completed__ps
      -- CP-element group 125: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_75_sample_start_
      -- CP-element group 125: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_75_sample_completed_
      -- 
    -- Element group access_T_CP_0_elements(125) is bound as output of CP function.
    -- CP-element group 126:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	128 
    -- CP-element group 126:  members (2) 
      -- CP-element group 126: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_75_update_start__ps
      -- CP-element group 126: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_75_update_start_
      -- 
    -- Element group access_T_CP_0_elements(126) is bound as output of CP function.
    -- CP-element group 127:  join  transition  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	128 
    -- CP-element group 127: successors 
    -- CP-element group 127:  members (1) 
      -- CP-element group 127: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_75_update_completed__ps
      -- 
    access_T_CP_0_elements(127) <= access_T_CP_0_elements(128);
    -- CP-element group 128:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	126 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	127 
    -- CP-element group 128:  members (1) 
      -- CP-element group 128: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_75_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(128) is a control-delay.
    cp_element_128_delay: control_delay_element  generic map(name => " 128_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(126), ack => access_T_CP_0_elements(128), clk => clk, reset =>reset);
    -- CP-element group 129:  join  transition  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	9 
    -- CP-element group 129: marked-predecessors 
    -- CP-element group 129: 	12 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	11 
    -- CP-element group 129:  members (1) 
      -- CP-element group 129: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_76_sample_start_
      -- 
    access_T_cp_element_group_129: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_129"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_129 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(129), clk => clk, reset => reset); --
    end block;
    -- CP-element group 130:  join  transition  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	9 
    -- CP-element group 130: marked-predecessors 
    -- CP-element group 130: 	134 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	13 
    -- CP-element group 130:  members (1) 
      -- CP-element group 130: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_76_update_start_
      -- 
    access_T_cp_element_group_130: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_130"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(134);
      gj_access_T_cp_element_group_130 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(130), clk => clk, reset => reset); --
    end block;
    -- CP-element group 131:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	11 
    -- CP-element group 131: successors 
    -- CP-element group 131:  members (1) 
      -- CP-element group 131: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_76_sample_start__ps
      -- 
    access_T_CP_0_elements(131) <= access_T_CP_0_elements(11);
    -- CP-element group 132:  join  transition  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	12 
    -- CP-element group 132:  members (1) 
      -- CP-element group 132: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_76_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(132) is bound as output of CP function.
    -- CP-element group 133:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	13 
    -- CP-element group 133: successors 
    -- CP-element group 133:  members (1) 
      -- CP-element group 133: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_76_update_start__ps
      -- 
    access_T_CP_0_elements(133) <= access_T_CP_0_elements(13);
    -- CP-element group 134:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	14 
    -- CP-element group 134: marked-successors 
    -- CP-element group 134: 	130 
    -- CP-element group 134:  members (2) 
      -- CP-element group 134: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_76_update_completed_
      -- CP-element group 134: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_76_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(134) is bound as output of CP function.
    -- CP-element group 135:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	7 
    -- CP-element group 135: successors 
    -- CP-element group 135:  members (1) 
      -- CP-element group 135: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_76_loopback_trigger
      -- 
    access_T_CP_0_elements(135) <= access_T_CP_0_elements(7);
    -- CP-element group 136:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: successors 
    -- CP-element group 136:  members (2) 
      -- CP-element group 136: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_76_loopback_sample_req
      -- CP-element group 136: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_76_loopback_sample_req_ps
      -- 
    phi_stmt_76_loopback_sample_req_328_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_76_loopback_sample_req_328_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(136), ack => phi_stmt_76_req_1); -- 
    -- Element group access_T_CP_0_elements(136) is bound as output of CP function.
    -- CP-element group 137:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	8 
    -- CP-element group 137: successors 
    -- CP-element group 137:  members (1) 
      -- CP-element group 137: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_76_entry_trigger
      -- 
    access_T_CP_0_elements(137) <= access_T_CP_0_elements(8);
    -- CP-element group 138:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: successors 
    -- CP-element group 138:  members (2) 
      -- CP-element group 138: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_76_entry_sample_req
      -- CP-element group 138: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_76_entry_sample_req_ps
      -- 
    phi_stmt_76_entry_sample_req_331_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_76_entry_sample_req_331_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(138), ack => phi_stmt_76_req_0); -- 
    -- Element group access_T_CP_0_elements(138) is bound as output of CP function.
    -- CP-element group 139:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: successors 
    -- CP-element group 139:  members (2) 
      -- CP-element group 139: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_76_phi_mux_ack
      -- CP-element group 139: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/phi_stmt_76_phi_mux_ack_ps
      -- 
    phi_stmt_76_phi_mux_ack_334_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_76_ack_0, ack => access_T_CP_0_elements(139)); -- 
    -- CP-element group 140:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: successors 
    -- CP-element group 140:  members (4) 
      -- CP-element group 140: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_79_sample_start__ps
      -- CP-element group 140: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_79_sample_completed__ps
      -- CP-element group 140: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_79_sample_start_
      -- CP-element group 140: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_79_sample_completed_
      -- 
    -- Element group access_T_CP_0_elements(140) is bound as output of CP function.
    -- CP-element group 141:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	143 
    -- CP-element group 141:  members (2) 
      -- CP-element group 141: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_79_update_start__ps
      -- CP-element group 141: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_79_update_start_
      -- 
    -- Element group access_T_CP_0_elements(141) is bound as output of CP function.
    -- CP-element group 142:  join  transition  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	143 
    -- CP-element group 142: successors 
    -- CP-element group 142:  members (1) 
      -- CP-element group 142: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_79_update_completed__ps
      -- 
    access_T_CP_0_elements(142) <= access_T_CP_0_elements(143);
    -- CP-element group 143:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	141 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	142 
    -- CP-element group 143:  members (1) 
      -- CP-element group 143: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/type_cast_79_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(143) is a control-delay.
    cp_element_143_delay: control_delay_element  generic map(name => " 143_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(141), ack => access_T_CP_0_elements(143), clk => clk, reset =>reset);
    -- CP-element group 144:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	146 
    -- CP-element group 144:  members (4) 
      -- CP-element group 144: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_row_80_sample_start__ps
      -- CP-element group 144: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_row_80_sample_start_
      -- CP-element group 144: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_row_80_Sample/$entry
      -- CP-element group 144: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_row_80_Sample/req
      -- 
    req_355_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_355_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(144), ack => n_row_234_80_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(144) is bound as output of CP function.
    -- CP-element group 145:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	147 
    -- CP-element group 145:  members (4) 
      -- CP-element group 145: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_row_80_update_start__ps
      -- CP-element group 145: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_row_80_update_start_
      -- CP-element group 145: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_row_80_Update/$entry
      -- CP-element group 145: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_row_80_Update/req
      -- 
    req_360_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_360_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(145), ack => n_row_234_80_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(145) is bound as output of CP function.
    -- CP-element group 146:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	144 
    -- CP-element group 146: successors 
    -- CP-element group 146:  members (4) 
      -- CP-element group 146: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_row_80_sample_completed__ps
      -- CP-element group 146: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_row_80_sample_completed_
      -- CP-element group 146: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_row_80_Sample/$exit
      -- CP-element group 146: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_row_80_Sample/ack
      -- 
    ack_356_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row_234_80_buf_ack_0, ack => access_T_CP_0_elements(146)); -- 
    -- CP-element group 147:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	145 
    -- CP-element group 147: successors 
    -- CP-element group 147:  members (4) 
      -- CP-element group 147: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_row_80_update_completed__ps
      -- CP-element group 147: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_row_80_update_completed_
      -- CP-element group 147: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_row_80_Update/$exit
      -- CP-element group 147: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/R_n_row_80_Update/ack
      -- 
    ack_361_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row_234_80_buf_ack_1, ack => access_T_CP_0_elements(147)); -- 
    -- CP-element group 148:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	152 
    -- CP-element group 148: marked-predecessors 
    -- CP-element group 148: 	153 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	153 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/addr_of_134_sample_start_
      -- CP-element group 148: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/addr_of_134_request/$entry
      -- CP-element group 148: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/addr_of_134_request/req
      -- 
    req_402_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_402_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(148), ack => addr_of_134_final_reg_req_0); -- 
    access_T_cp_element_group_148: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_148"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(152) & access_T_CP_0_elements(153);
      gj_access_T_cp_element_group_148 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(148), clk => clk, reset => reset); --
    end block;
    -- CP-element group 149:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	9 
    -- CP-element group 149: marked-predecessors 
    -- CP-element group 149: 	157 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	154 
    -- CP-element group 149:  members (3) 
      -- CP-element group 149: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/addr_of_134_update_start_
      -- CP-element group 149: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/addr_of_134_complete/$entry
      -- CP-element group 149: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/addr_of_134_complete/req
      -- 
    req_407_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_407_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(149), ack => addr_of_134_final_reg_req_1); -- 
    access_T_cp_element_group_149: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_149"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(157);
      gj_access_T_cp_element_group_149 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(149), clk => clk, reset => reset); --
    end block;
    -- CP-element group 150:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	9 
    -- CP-element group 150: marked-predecessors 
    -- CP-element group 150: 	153 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	152 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_final_index_sum_regn_update_start
      -- CP-element group 150: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_final_index_sum_regn_Update/$entry
      -- CP-element group 150: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_final_index_sum_regn_Update/req
      -- 
    req_392_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_392_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(150), ack => array_obj_ref_133_index_offset_req_1); -- 
    access_T_cp_element_group_150: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_150"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(153);
      gj_access_T_cp_element_group_150 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(150), clk => clk, reset => reset); --
    end block;
    -- CP-element group 151:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	20 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	204 
    -- CP-element group 151: marked-successors 
    -- CP-element group 151: 	16 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_final_index_sum_regn_sample_complete
      -- CP-element group 151: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_final_index_sum_regn_Sample/$exit
      -- CP-element group 151: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_final_index_sum_regn_Sample/ack
      -- 
    ack_388_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_133_index_offset_ack_0, ack => access_T_CP_0_elements(151)); -- 
    -- CP-element group 152:  transition  input  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	150 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	148 
    -- CP-element group 152:  members (8) 
      -- CP-element group 152: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_root_address_calculated
      -- CP-element group 152: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_offset_calculated
      -- CP-element group 152: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_final_index_sum_regn_Update/$exit
      -- CP-element group 152: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_final_index_sum_regn_Update/ack
      -- CP-element group 152: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_base_plus_offset/$entry
      -- CP-element group 152: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_base_plus_offset/$exit
      -- CP-element group 152: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_base_plus_offset/sum_rename_req
      -- CP-element group 152: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/array_obj_ref_133_base_plus_offset/sum_rename_ack
      -- 
    ack_393_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_133_index_offset_ack_1, ack => access_T_CP_0_elements(152)); -- 
    -- CP-element group 153:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	148 
    -- CP-element group 153: successors 
    -- CP-element group 153: marked-successors 
    -- CP-element group 153: 	148 
    -- CP-element group 153: 	150 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/addr_of_134_sample_completed_
      -- CP-element group 153: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/addr_of_134_request/$exit
      -- CP-element group 153: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/addr_of_134_request/ack
      -- 
    ack_403_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_134_final_reg_ack_0, ack => access_T_CP_0_elements(153)); -- 
    -- CP-element group 154:  transition  input  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	149 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	155 
    -- CP-element group 154:  members (19) 
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/addr_of_134_update_completed_
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/addr_of_134_complete/$exit
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/addr_of_134_complete/ack
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_base_address_calculated
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_word_address_calculated
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_root_address_calculated
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_base_address_resized
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_base_addr_resize/$entry
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_base_addr_resize/$exit
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_base_addr_resize/base_resize_req
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_base_addr_resize/base_resize_ack
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_base_plus_offset/$entry
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_base_plus_offset/$exit
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_base_plus_offset/sum_rename_req
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_base_plus_offset/sum_rename_ack
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_word_addrgen/$entry
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_word_addrgen/$exit
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_word_addrgen/root_register_req
      -- CP-element group 154: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_word_addrgen/root_register_ack
      -- 
    ack_408_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_134_final_reg_ack_1, ack => access_T_CP_0_elements(154)); -- 
    -- CP-element group 155:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	154 
    -- CP-element group 155: marked-predecessors 
    -- CP-element group 155: 	157 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	157 
    -- CP-element group 155:  members (5) 
      -- CP-element group 155: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_sample_start_
      -- CP-element group 155: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Sample/$entry
      -- CP-element group 155: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Sample/word_access_start/$entry
      -- CP-element group 155: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Sample/word_access_start/word_0/$entry
      -- CP-element group 155: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Sample/word_access_start/word_0/rr
      -- 
    rr_441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(155), ack => ptr_deref_138_load_0_req_0); -- 
    access_T_cp_element_group_155: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_155"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(154) & access_T_CP_0_elements(157);
      gj_access_T_cp_element_group_155 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(155), clk => clk, reset => reset); --
    end block;
    -- CP-element group 156:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: marked-predecessors 
    -- CP-element group 156: 	161 
    -- CP-element group 156: 	165 
    -- CP-element group 156: 	169 
    -- CP-element group 156: 	173 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	158 
    -- CP-element group 156:  members (5) 
      -- CP-element group 156: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_update_start_
      -- CP-element group 156: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Update/$entry
      -- CP-element group 156: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Update/word_access_complete/$entry
      -- CP-element group 156: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Update/word_access_complete/word_0/$entry
      -- CP-element group 156: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Update/word_access_complete/word_0/cr
      -- 
    cr_452_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_452_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(156), ack => ptr_deref_138_load_0_req_1); -- 
    access_T_cp_element_group_156: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_156"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(161) & access_T_CP_0_elements(165) & access_T_CP_0_elements(169) & access_T_CP_0_elements(173);
      gj_access_T_cp_element_group_156 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(156), clk => clk, reset => reset); --
    end block;
    -- CP-element group 157:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	155 
    -- CP-element group 157: successors 
    -- CP-element group 157: marked-successors 
    -- CP-element group 157: 	149 
    -- CP-element group 157: 	155 
    -- CP-element group 157:  members (5) 
      -- CP-element group 157: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_sample_completed_
      -- CP-element group 157: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Sample/$exit
      -- CP-element group 157: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Sample/word_access_start/$exit
      -- CP-element group 157: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Sample/word_access_start/word_0/$exit
      -- CP-element group 157: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Sample/word_access_start/word_0/ra
      -- 
    ra_442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_138_load_0_ack_0, ack => access_T_CP_0_elements(157)); -- 
    -- CP-element group 158:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	156 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	159 
    -- CP-element group 158: 	163 
    -- CP-element group 158: 	167 
    -- CP-element group 158: 	171 
    -- CP-element group 158:  members (9) 
      -- CP-element group 158: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_update_completed_
      -- CP-element group 158: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Update/$exit
      -- CP-element group 158: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Update/word_access_complete/$exit
      -- CP-element group 158: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Update/word_access_complete/word_0/$exit
      -- CP-element group 158: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Update/word_access_complete/word_0/ca
      -- CP-element group 158: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Update/ptr_deref_138_Merge/$entry
      -- CP-element group 158: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Update/ptr_deref_138_Merge/$exit
      -- CP-element group 158: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Update/ptr_deref_138_Merge/merge_req
      -- CP-element group 158: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/ptr_deref_138_Update/ptr_deref_138_Merge/merge_ack
      -- 
    ca_453_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_138_load_0_ack_1, ack => access_T_CP_0_elements(158)); -- 
    -- CP-element group 159:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	158 
    -- CP-element group 159: marked-predecessors 
    -- CP-element group 159: 	161 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	161 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_142_sample_start_
      -- CP-element group 159: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_142_Sample/$entry
      -- CP-element group 159: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_142_Sample/rr
      -- 
    rr_466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(159), ack => slice_142_inst_req_0); -- 
    access_T_cp_element_group_159: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_159"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(158) & access_T_CP_0_elements(161);
      gj_access_T_cp_element_group_159 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(159), clk => clk, reset => reset); --
    end block;
    -- CP-element group 160:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: marked-predecessors 
    -- CP-element group 160: 	180 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	162 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_142_update_start_
      -- CP-element group 160: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_142_Update/$entry
      -- CP-element group 160: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_142_Update/cr
      -- 
    cr_471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(160), ack => slice_142_inst_req_1); -- 
    access_T_cp_element_group_160: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_160"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(180);
      gj_access_T_cp_element_group_160 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(160), clk => clk, reset => reset); --
    end block;
    -- CP-element group 161:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	159 
    -- CP-element group 161: successors 
    -- CP-element group 161: marked-successors 
    -- CP-element group 161: 	156 
    -- CP-element group 161: 	159 
    -- CP-element group 161:  members (3) 
      -- CP-element group 161: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_142_sample_completed_
      -- CP-element group 161: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_142_Sample/$exit
      -- CP-element group 161: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_142_Sample/ra
      -- 
    ra_467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_142_inst_ack_0, ack => access_T_CP_0_elements(161)); -- 
    -- CP-element group 162:  transition  input  bypass  pipeline-parent 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	160 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	179 
    -- CP-element group 162:  members (3) 
      -- CP-element group 162: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_142_update_completed_
      -- CP-element group 162: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_142_Update/$exit
      -- CP-element group 162: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_142_Update/ca
      -- 
    ca_472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_142_inst_ack_1, ack => access_T_CP_0_elements(162)); -- 
    -- CP-element group 163:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	158 
    -- CP-element group 163: marked-predecessors 
    -- CP-element group 163: 	165 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	165 
    -- CP-element group 163:  members (3) 
      -- CP-element group 163: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_146_sample_start_
      -- CP-element group 163: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_146_Sample/$entry
      -- CP-element group 163: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_146_Sample/rr
      -- 
    rr_480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(163), ack => slice_146_inst_req_0); -- 
    access_T_cp_element_group_163: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_163"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(158) & access_T_CP_0_elements(165);
      gj_access_T_cp_element_group_163 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(163), clk => clk, reset => reset); --
    end block;
    -- CP-element group 164:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: marked-predecessors 
    -- CP-element group 164: 	187 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	166 
    -- CP-element group 164:  members (3) 
      -- CP-element group 164: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_146_update_start_
      -- CP-element group 164: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_146_Update/$entry
      -- CP-element group 164: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_146_Update/cr
      -- 
    cr_485_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_485_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(164), ack => slice_146_inst_req_1); -- 
    access_T_cp_element_group_164: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_164"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(187);
      gj_access_T_cp_element_group_164 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(164), clk => clk, reset => reset); --
    end block;
    -- CP-element group 165:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	163 
    -- CP-element group 165: successors 
    -- CP-element group 165: marked-successors 
    -- CP-element group 165: 	156 
    -- CP-element group 165: 	163 
    -- CP-element group 165:  members (3) 
      -- CP-element group 165: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_146_sample_completed_
      -- CP-element group 165: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_146_Sample/$exit
      -- CP-element group 165: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_146_Sample/ra
      -- 
    ra_481_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_146_inst_ack_0, ack => access_T_CP_0_elements(165)); -- 
    -- CP-element group 166:  transition  input  bypass  pipeline-parent 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	164 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	186 
    -- CP-element group 166:  members (3) 
      -- CP-element group 166: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_146_update_completed_
      -- CP-element group 166: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_146_Update/$exit
      -- CP-element group 166: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_146_Update/ca
      -- 
    ca_486_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_146_inst_ack_1, ack => access_T_CP_0_elements(166)); -- 
    -- CP-element group 167:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	158 
    -- CP-element group 167: marked-predecessors 
    -- CP-element group 167: 	169 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	169 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_150_sample_start_
      -- CP-element group 167: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_150_Sample/$entry
      -- CP-element group 167: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_150_Sample/rr
      -- 
    rr_494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(167), ack => slice_150_inst_req_0); -- 
    access_T_cp_element_group_167: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_167"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(158) & access_T_CP_0_elements(169);
      gj_access_T_cp_element_group_167 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(167), clk => clk, reset => reset); --
    end block;
    -- CP-element group 168:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: marked-predecessors 
    -- CP-element group 168: 	194 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	170 
    -- CP-element group 168:  members (3) 
      -- CP-element group 168: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_150_update_start_
      -- CP-element group 168: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_150_Update/$entry
      -- CP-element group 168: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_150_Update/cr
      -- 
    cr_499_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_499_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(168), ack => slice_150_inst_req_1); -- 
    access_T_cp_element_group_168: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_168"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(194);
      gj_access_T_cp_element_group_168 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(168), clk => clk, reset => reset); --
    end block;
    -- CP-element group 169:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	167 
    -- CP-element group 169: successors 
    -- CP-element group 169: marked-successors 
    -- CP-element group 169: 	156 
    -- CP-element group 169: 	167 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_150_sample_completed_
      -- CP-element group 169: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_150_Sample/$exit
      -- CP-element group 169: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_150_Sample/ra
      -- 
    ra_495_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_150_inst_ack_0, ack => access_T_CP_0_elements(169)); -- 
    -- CP-element group 170:  transition  input  bypass  pipeline-parent 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	168 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	193 
    -- CP-element group 170:  members (3) 
      -- CP-element group 170: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_150_update_completed_
      -- CP-element group 170: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_150_Update/$exit
      -- CP-element group 170: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_150_Update/ca
      -- 
    ca_500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_150_inst_ack_1, ack => access_T_CP_0_elements(170)); -- 
    -- CP-element group 171:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	158 
    -- CP-element group 171: marked-predecessors 
    -- CP-element group 171: 	173 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	173 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_154_sample_start_
      -- CP-element group 171: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_154_Sample/$entry
      -- CP-element group 171: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_154_Sample/rr
      -- 
    rr_508_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_508_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(171), ack => slice_154_inst_req_0); -- 
    access_T_cp_element_group_171: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_171"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(158) & access_T_CP_0_elements(173);
      gj_access_T_cp_element_group_171 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(171), clk => clk, reset => reset); --
    end block;
    -- CP-element group 172:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: marked-predecessors 
    -- CP-element group 172: 	201 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	174 
    -- CP-element group 172:  members (3) 
      -- CP-element group 172: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_154_update_start_
      -- CP-element group 172: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_154_Update/$entry
      -- CP-element group 172: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_154_Update/cr
      -- 
    cr_513_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_513_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(172), ack => slice_154_inst_req_1); -- 
    access_T_cp_element_group_172: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_172"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(201);
      gj_access_T_cp_element_group_172 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(172), clk => clk, reset => reset); --
    end block;
    -- CP-element group 173:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	171 
    -- CP-element group 173: successors 
    -- CP-element group 173: marked-successors 
    -- CP-element group 173: 	156 
    -- CP-element group 173: 	171 
    -- CP-element group 173:  members (3) 
      -- CP-element group 173: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_154_sample_completed_
      -- CP-element group 173: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_154_Sample/$exit
      -- CP-element group 173: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_154_Sample/ra
      -- 
    ra_509_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_154_inst_ack_0, ack => access_T_CP_0_elements(173)); -- 
    -- CP-element group 174:  transition  input  bypass  pipeline-parent 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	172 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	200 
    -- CP-element group 174:  members (3) 
      -- CP-element group 174: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_154_update_completed_
      -- CP-element group 174: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_154_Update/$exit
      -- CP-element group 174: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/slice_154_Update/ca
      -- 
    ca_514_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_154_inst_ack_1, ack => access_T_CP_0_elements(174)); -- 
    -- CP-element group 175:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	39 
    -- CP-element group 175: marked-predecessors 
    -- CP-element group 175: 	177 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	177 
    -- CP-element group 175:  members (3) 
      -- CP-element group 175: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_158_sample_start_
      -- CP-element group 175: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_158_Sample/$entry
      -- CP-element group 175: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_158_Sample/req
      -- 
    req_522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(175), ack => W_c1_156_delayed_14_0_156_inst_req_0); -- 
    access_T_cp_element_group_175: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_175"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(39) & access_T_CP_0_elements(177);
      gj_access_T_cp_element_group_175 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(175), clk => clk, reset => reset); --
    end block;
    -- CP-element group 176:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: marked-predecessors 
    -- CP-element group 176: 	180 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	178 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_158_update_start_
      -- CP-element group 176: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_158_Update/$entry
      -- CP-element group 176: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_158_Update/req
      -- 
    req_527_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_527_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(176), ack => W_c1_156_delayed_14_0_156_inst_req_1); -- 
    access_T_cp_element_group_176: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_176"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(180);
      gj_access_T_cp_element_group_176 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(176), clk => clk, reset => reset); --
    end block;
    -- CP-element group 177:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	175 
    -- CP-element group 177: successors 
    -- CP-element group 177: marked-successors 
    -- CP-element group 177: 	35 
    -- CP-element group 177: 	175 
    -- CP-element group 177:  members (3) 
      -- CP-element group 177: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_158_sample_completed_
      -- CP-element group 177: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_158_Sample/$exit
      -- CP-element group 177: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_158_Sample/ack
      -- 
    ack_523_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_c1_156_delayed_14_0_156_inst_ack_0, ack => access_T_CP_0_elements(177)); -- 
    -- CP-element group 178:  transition  input  bypass  pipeline-parent 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	176 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	179 
    -- CP-element group 178:  members (3) 
      -- CP-element group 178: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_158_update_completed_
      -- CP-element group 178: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_158_Update/$exit
      -- CP-element group 178: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_158_Update/ack
      -- 
    ack_528_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_c1_156_delayed_14_0_156_inst_ack_1, ack => access_T_CP_0_elements(178)); -- 
    -- CP-element group 179:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	162 
    -- CP-element group 179: 	178 
    -- CP-element group 179: marked-predecessors 
    -- CP-element group 179: 	202 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	180 
    -- CP-element group 179:  members (3) 
      -- CP-element group 179: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_160_sample_start_
      -- CP-element group 179: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_160_Sample/$entry
      -- CP-element group 179: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_160_Sample/req
      -- 
    req_536_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_536_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(179), ack => WPIPE_input_pipe1_160_inst_req_0); -- 
    access_T_cp_element_group_179: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_179"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(162) & access_T_CP_0_elements(178) & access_T_CP_0_elements(202);
      gj_access_T_cp_element_group_179 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(179), clk => clk, reset => reset); --
    end block;
    -- CP-element group 180:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	179 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	181 
    -- CP-element group 180: marked-successors 
    -- CP-element group 180: 	160 
    -- CP-element group 180: 	176 
    -- CP-element group 180:  members (6) 
      -- CP-element group 180: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_160_sample_completed_
      -- CP-element group 180: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_160_update_start_
      -- CP-element group 180: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_160_Sample/$exit
      -- CP-element group 180: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_160_Sample/ack
      -- CP-element group 180: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_160_Update/$entry
      -- CP-element group 180: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_160_Update/req
      -- 
    ack_537_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_160_inst_ack_0, ack => access_T_CP_0_elements(180)); -- 
    req_541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(180), ack => WPIPE_input_pipe1_160_inst_req_1); -- 
    -- CP-element group 181:  transition  input  bypass  pipeline-parent 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	180 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	186 
    -- CP-element group 181:  members (3) 
      -- CP-element group 181: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_160_update_completed_
      -- CP-element group 181: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_160_Update/$exit
      -- CP-element group 181: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_160_Update/ack
      -- 
    ack_542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_160_inst_ack_1, ack => access_T_CP_0_elements(181)); -- 
    -- CP-element group 182:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	75 
    -- CP-element group 182: 	39 
    -- CP-element group 182: marked-predecessors 
    -- CP-element group 182: 	184 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	184 
    -- CP-element group 182:  members (3) 
      -- CP-element group 182: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_165_sample_start_
      -- CP-element group 182: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_165_Sample/$entry
      -- CP-element group 182: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_165_Sample/req
      -- 
    req_550_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_550_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(182), ack => W_c2_160_delayed_14_0_163_inst_req_0); -- 
    access_T_cp_element_group_182: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_182"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(75) & access_T_CP_0_elements(39) & access_T_CP_0_elements(184);
      gj_access_T_cp_element_group_182 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(182), clk => clk, reset => reset); --
    end block;
    -- CP-element group 183:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: marked-predecessors 
    -- CP-element group 183: 	187 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	185 
    -- CP-element group 183:  members (3) 
      -- CP-element group 183: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_165_update_start_
      -- CP-element group 183: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_165_Update/$entry
      -- CP-element group 183: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_165_Update/req
      -- 
    req_555_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_555_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(183), ack => W_c2_160_delayed_14_0_163_inst_req_1); -- 
    access_T_cp_element_group_183: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_183"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(187);
      gj_access_T_cp_element_group_183 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(183), clk => clk, reset => reset); --
    end block;
    -- CP-element group 184:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	182 
    -- CP-element group 184: successors 
    -- CP-element group 184: marked-successors 
    -- CP-element group 184: 	73 
    -- CP-element group 184: 	35 
    -- CP-element group 184: 	182 
    -- CP-element group 184:  members (3) 
      -- CP-element group 184: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_165_sample_completed_
      -- CP-element group 184: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_165_Sample/$exit
      -- CP-element group 184: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_165_Sample/ack
      -- 
    ack_551_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_c2_160_delayed_14_0_163_inst_ack_0, ack => access_T_CP_0_elements(184)); -- 
    -- CP-element group 185:  transition  input  bypass  pipeline-parent 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	183 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	186 
    -- CP-element group 185:  members (3) 
      -- CP-element group 185: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_165_update_completed_
      -- CP-element group 185: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_165_Update/$exit
      -- CP-element group 185: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_165_Update/ack
      -- 
    ack_556_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_c2_160_delayed_14_0_163_inst_ack_1, ack => access_T_CP_0_elements(185)); -- 
    -- CP-element group 186:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	181 
    -- CP-element group 186: 	185 
    -- CP-element group 186: 	166 
    -- CP-element group 186: marked-predecessors 
    -- CP-element group 186: 	188 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	187 
    -- CP-element group 186:  members (3) 
      -- CP-element group 186: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_167_sample_start_
      -- CP-element group 186: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_167_Sample/$entry
      -- CP-element group 186: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_167_Sample/req
      -- 
    req_564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(186), ack => WPIPE_input_pipe1_167_inst_req_0); -- 
    access_T_cp_element_group_186: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_186"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(181) & access_T_CP_0_elements(185) & access_T_CP_0_elements(166) & access_T_CP_0_elements(188);
      gj_access_T_cp_element_group_186 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(186), clk => clk, reset => reset); --
    end block;
    -- CP-element group 187:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	186 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	188 
    -- CP-element group 187: marked-successors 
    -- CP-element group 187: 	183 
    -- CP-element group 187: 	164 
    -- CP-element group 187:  members (6) 
      -- CP-element group 187: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_167_Sample/ack
      -- CP-element group 187: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_167_Update/$entry
      -- CP-element group 187: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_167_Update/req
      -- CP-element group 187: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_167_sample_completed_
      -- CP-element group 187: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_167_update_start_
      -- CP-element group 187: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_167_Sample/$exit
      -- 
    ack_565_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_167_inst_ack_0, ack => access_T_CP_0_elements(187)); -- 
    req_569_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_569_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(187), ack => WPIPE_input_pipe1_167_inst_req_1); -- 
    -- CP-element group 188:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	187 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	193 
    -- CP-element group 188: marked-successors 
    -- CP-element group 188: 	186 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_167_Update/$exit
      -- CP-element group 188: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_167_Update/ack
      -- CP-element group 188: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_167_update_completed_
      -- 
    ack_570_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_167_inst_ack_1, ack => access_T_CP_0_elements(188)); -- 
    -- CP-element group 189:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	75 
    -- CP-element group 189: 	39 
    -- CP-element group 189: marked-predecessors 
    -- CP-element group 189: 	191 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	191 
    -- CP-element group 189:  members (3) 
      -- CP-element group 189: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_172_sample_start_
      -- CP-element group 189: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_172_Sample/$entry
      -- CP-element group 189: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_172_Sample/req
      -- 
    req_578_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_578_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(189), ack => W_c3_164_delayed_14_0_170_inst_req_0); -- 
    access_T_cp_element_group_189: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_189"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(75) & access_T_CP_0_elements(39) & access_T_CP_0_elements(191);
      gj_access_T_cp_element_group_189 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(189), clk => clk, reset => reset); --
    end block;
    -- CP-element group 190:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: marked-predecessors 
    -- CP-element group 190: 	194 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	192 
    -- CP-element group 190:  members (3) 
      -- CP-element group 190: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_172_update_start_
      -- CP-element group 190: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_172_Update/$entry
      -- CP-element group 190: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_172_Update/req
      -- 
    req_583_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_583_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(190), ack => W_c3_164_delayed_14_0_170_inst_req_1); -- 
    access_T_cp_element_group_190: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_190"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(194);
      gj_access_T_cp_element_group_190 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(190), clk => clk, reset => reset); --
    end block;
    -- CP-element group 191:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	189 
    -- CP-element group 191: successors 
    -- CP-element group 191: marked-successors 
    -- CP-element group 191: 	73 
    -- CP-element group 191: 	35 
    -- CP-element group 191: 	189 
    -- CP-element group 191:  members (3) 
      -- CP-element group 191: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_172_sample_completed_
      -- CP-element group 191: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_172_Sample/$exit
      -- CP-element group 191: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_172_Sample/ack
      -- 
    ack_579_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_c3_164_delayed_14_0_170_inst_ack_0, ack => access_T_CP_0_elements(191)); -- 
    -- CP-element group 192:  transition  input  bypass  pipeline-parent 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	190 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	193 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_172_update_completed_
      -- CP-element group 192: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_172_Update/$exit
      -- CP-element group 192: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_172_Update/ack
      -- 
    ack_584_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_c3_164_delayed_14_0_170_inst_ack_1, ack => access_T_CP_0_elements(192)); -- 
    -- CP-element group 193:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	192 
    -- CP-element group 193: 	188 
    -- CP-element group 193: 	170 
    -- CP-element group 193: marked-predecessors 
    -- CP-element group 193: 	195 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	194 
    -- CP-element group 193:  members (3) 
      -- CP-element group 193: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_174_sample_start_
      -- CP-element group 193: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_174_Sample/$entry
      -- CP-element group 193: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_174_Sample/req
      -- 
    req_592_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_592_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(193), ack => WPIPE_input_pipe1_174_inst_req_0); -- 
    access_T_cp_element_group_193: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_193"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(192) & access_T_CP_0_elements(188) & access_T_CP_0_elements(170) & access_T_CP_0_elements(195);
      gj_access_T_cp_element_group_193 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(193), clk => clk, reset => reset); --
    end block;
    -- CP-element group 194:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	193 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	195 
    -- CP-element group 194: marked-successors 
    -- CP-element group 194: 	190 
    -- CP-element group 194: 	168 
    -- CP-element group 194:  members (6) 
      -- CP-element group 194: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_174_sample_completed_
      -- CP-element group 194: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_174_update_start_
      -- CP-element group 194: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_174_Sample/$exit
      -- CP-element group 194: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_174_Sample/ack
      -- CP-element group 194: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_174_Update/$entry
      -- CP-element group 194: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_174_Update/req
      -- 
    ack_593_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_174_inst_ack_0, ack => access_T_CP_0_elements(194)); -- 
    req_597_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_597_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(194), ack => WPIPE_input_pipe1_174_inst_req_1); -- 
    -- CP-element group 195:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	194 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	200 
    -- CP-element group 195: marked-successors 
    -- CP-element group 195: 	193 
    -- CP-element group 195:  members (3) 
      -- CP-element group 195: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_174_update_completed_
      -- CP-element group 195: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_174_Update/$exit
      -- CP-element group 195: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_174_Update/ack
      -- 
    ack_598_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_174_inst_ack_1, ack => access_T_CP_0_elements(195)); -- 
    -- CP-element group 196:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	75 
    -- CP-element group 196: 	39 
    -- CP-element group 196: marked-predecessors 
    -- CP-element group 196: 	198 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	198 
    -- CP-element group 196:  members (3) 
      -- CP-element group 196: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_179_sample_start_
      -- CP-element group 196: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_179_Sample/$entry
      -- CP-element group 196: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_179_Sample/req
      -- 
    req_606_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_606_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(196), ack => W_c4_168_delayed_14_0_177_inst_req_0); -- 
    access_T_cp_element_group_196: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_196"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(75) & access_T_CP_0_elements(39) & access_T_CP_0_elements(198);
      gj_access_T_cp_element_group_196 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(196), clk => clk, reset => reset); --
    end block;
    -- CP-element group 197:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: marked-predecessors 
    -- CP-element group 197: 	201 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	199 
    -- CP-element group 197:  members (3) 
      -- CP-element group 197: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_179_update_start_
      -- CP-element group 197: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_179_Update/$entry
      -- CP-element group 197: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_179_Update/req
      -- 
    req_611_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_611_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(197), ack => W_c4_168_delayed_14_0_177_inst_req_1); -- 
    access_T_cp_element_group_197: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_197"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(201);
      gj_access_T_cp_element_group_197 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(197), clk => clk, reset => reset); --
    end block;
    -- CP-element group 198:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	196 
    -- CP-element group 198: successors 
    -- CP-element group 198: marked-successors 
    -- CP-element group 198: 	73 
    -- CP-element group 198: 	35 
    -- CP-element group 198: 	196 
    -- CP-element group 198:  members (3) 
      -- CP-element group 198: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_179_sample_completed_
      -- CP-element group 198: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_179_Sample/$exit
      -- CP-element group 198: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_179_Sample/ack
      -- 
    ack_607_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_c4_168_delayed_14_0_177_inst_ack_0, ack => access_T_CP_0_elements(198)); -- 
    -- CP-element group 199:  transition  input  bypass  pipeline-parent 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	197 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	200 
    -- CP-element group 199:  members (3) 
      -- CP-element group 199: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_179_update_completed_
      -- CP-element group 199: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_179_Update/$exit
      -- CP-element group 199: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/assign_stmt_179_Update/ack
      -- 
    ack_612_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_c4_168_delayed_14_0_177_inst_ack_1, ack => access_T_CP_0_elements(199)); -- 
    -- CP-element group 200:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	195 
    -- CP-element group 200: 	199 
    -- CP-element group 200: 	174 
    -- CP-element group 200: marked-predecessors 
    -- CP-element group 200: 	202 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	201 
    -- CP-element group 200:  members (3) 
      -- CP-element group 200: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_181_sample_start_
      -- CP-element group 200: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_181_Sample/$entry
      -- CP-element group 200: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_181_Sample/req
      -- 
    req_620_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_620_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(200), ack => WPIPE_input_pipe1_181_inst_req_0); -- 
    access_T_cp_element_group_200: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_200"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(195) & access_T_CP_0_elements(199) & access_T_CP_0_elements(174) & access_T_CP_0_elements(202);
      gj_access_T_cp_element_group_200 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(200), clk => clk, reset => reset); --
    end block;
    -- CP-element group 201:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	200 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	202 
    -- CP-element group 201: marked-successors 
    -- CP-element group 201: 	197 
    -- CP-element group 201: 	172 
    -- CP-element group 201:  members (6) 
      -- CP-element group 201: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_181_sample_completed_
      -- CP-element group 201: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_181_update_start_
      -- CP-element group 201: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_181_Sample/$exit
      -- CP-element group 201: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_181_Sample/ack
      -- CP-element group 201: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_181_Update/$entry
      -- CP-element group 201: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_181_Update/req
      -- 
    ack_621_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_181_inst_ack_0, ack => access_T_CP_0_elements(201)); -- 
    req_625_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_625_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(201), ack => WPIPE_input_pipe1_181_inst_req_1); -- 
    -- CP-element group 202:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	201 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	204 
    -- CP-element group 202: marked-successors 
    -- CP-element group 202: 	200 
    -- CP-element group 202: 	179 
    -- CP-element group 202:  members (3) 
      -- CP-element group 202: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_181_update_completed_
      -- CP-element group 202: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_181_Update/$exit
      -- CP-element group 202: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/WPIPE_input_pipe1_181_Update/ack
      -- 
    ack_626_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_181_inst_ack_1, ack => access_T_CP_0_elements(202)); -- 
    -- CP-element group 203:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	9 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	10 
    -- CP-element group 203:  members (1) 
      -- CP-element group 203: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group access_T_CP_0_elements(203) is a control-delay.
    cp_element_203_delay: control_delay_element  generic map(name => " 203_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(9), ack => access_T_CP_0_elements(203), clk => clk, reset =>reset);
    -- CP-element group 204:  join  transition  bypass  pipeline-parent 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	202 
    -- CP-element group 204: 	12 
    -- CP-element group 204: 	151 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	6 
    -- CP-element group 204:  members (1) 
      -- CP-element group 204: 	 branch_block_stmt_26/do_while_stmt_44/do_while_stmt_44_loop_body/$exit
      -- 
    access_T_cp_element_group_204: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_204"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(202) & access_T_CP_0_elements(12) & access_T_CP_0_elements(151);
      gj_access_T_cp_element_group_204 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(204), clk => clk, reset => reset); --
    end block;
    -- CP-element group 205:  transition  input  bypass  pipeline-parent 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	5 
    -- CP-element group 205: successors 
    -- CP-element group 205:  members (2) 
      -- CP-element group 205: 	 branch_block_stmt_26/do_while_stmt_44/loop_exit/$exit
      -- CP-element group 205: 	 branch_block_stmt_26/do_while_stmt_44/loop_exit/ack
      -- 
    ack_631_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_44_branch_ack_0, ack => access_T_CP_0_elements(205)); -- 
    -- CP-element group 206:  transition  input  bypass  pipeline-parent 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	5 
    -- CP-element group 206: successors 
    -- CP-element group 206:  members (2) 
      -- CP-element group 206: 	 branch_block_stmt_26/do_while_stmt_44/loop_taken/$exit
      -- CP-element group 206: 	 branch_block_stmt_26/do_while_stmt_44/loop_taken/ack
      -- 
    ack_635_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 206_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_44_branch_ack_1, ack => access_T_CP_0_elements(206)); -- 
    -- CP-element group 207:  transition  bypass  pipeline-parent 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	3 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	1 
    -- CP-element group 207:  members (1) 
      -- CP-element group 207: 	 branch_block_stmt_26/do_while_stmt_44/$exit
      -- 
    access_T_CP_0_elements(207) <= access_T_CP_0_elements(3);
    access_T_do_while_stmt_44_terminator_636: loop_terminator -- 
      generic map (name => " access_T_do_while_stmt_44_terminator_636", max_iterations_in_flight =>15) 
      port map(loop_body_exit => access_T_CP_0_elements(6),loop_continue => access_T_CP_0_elements(206),loop_terminate => access_T_CP_0_elements(205),loop_back => access_T_CP_0_elements(4),loop_exit => access_T_CP_0_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_46_phi_seq_78_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(23);
      access_T_CP_0_elements(26)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(26);
      access_T_CP_0_elements(27)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(28);
      access_T_CP_0_elements(24) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(21);
      access_T_CP_0_elements(30)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(32);
      access_T_CP_0_elements(31)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(33);
      access_T_CP_0_elements(22) <= phi_mux_reqs(1);
      phi_stmt_46_phi_seq_78 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_46_phi_seq_78") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(17), 
          phi_sample_ack => access_T_CP_0_elements(18), 
          phi_update_req => access_T_CP_0_elements(19), 
          phi_update_ack => access_T_CP_0_elements(20), 
          phi_mux_ack => access_T_CP_0_elements(25), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_51_phi_seq_122_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(42);
      access_T_CP_0_elements(45)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(45);
      access_T_CP_0_elements(46)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(47);
      access_T_CP_0_elements(43) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(40);
      access_T_CP_0_elements(49)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(51);
      access_T_CP_0_elements(50)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(52);
      access_T_CP_0_elements(41) <= phi_mux_reqs(1);
      phi_stmt_51_phi_seq_122 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_51_phi_seq_122") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(36), 
          phi_sample_ack => access_T_CP_0_elements(37), 
          phi_update_req => access_T_CP_0_elements(38), 
          phi_update_ack => access_T_CP_0_elements(39), 
          phi_mux_ack => access_T_CP_0_elements(44), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_57_phi_seq_176_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(61);
      access_T_CP_0_elements(64)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(66);
      access_T_CP_0_elements(65)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(67);
      access_T_CP_0_elements(62) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(59);
      access_T_CP_0_elements(68)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(70);
      access_T_CP_0_elements(69)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(71);
      access_T_CP_0_elements(60) <= phi_mux_reqs(1);
      phi_stmt_57_phi_seq_176 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_57_phi_seq_176") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(55), 
          phi_sample_ack => access_T_CP_0_elements(56), 
          phi_update_req => access_T_CP_0_elements(57), 
          phi_update_ack => access_T_CP_0_elements(58), 
          phi_mux_ack => access_T_CP_0_elements(63), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_61_phi_seq_230_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(78);
      access_T_CP_0_elements(81)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(85);
      access_T_CP_0_elements(82)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(86);
      access_T_CP_0_elements(79) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(76);
      access_T_CP_0_elements(87)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(89);
      access_T_CP_0_elements(88)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(90);
      access_T_CP_0_elements(77) <= phi_mux_reqs(1);
      phi_stmt_61_phi_seq_230 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_61_phi_seq_230") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(11), 
          phi_sample_ack => access_T_CP_0_elements(74), 
          phi_update_req => access_T_CP_0_elements(13), 
          phi_update_ack => access_T_CP_0_elements(75), 
          phi_mux_ack => access_T_CP_0_elements(80), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_66_phi_seq_274_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(97);
      access_T_CP_0_elements(102)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(104);
      access_T_CP_0_elements(103)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(105);
      access_T_CP_0_elements(98) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(99);
      access_T_CP_0_elements(106)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(106);
      access_T_CP_0_elements(107)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(108);
      access_T_CP_0_elements(100) <= phi_mux_reqs(1);
      phi_stmt_66_phi_seq_274 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_66_phi_seq_274") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(93), 
          phi_sample_ack => access_T_CP_0_elements(94), 
          phi_update_req => access_T_CP_0_elements(95), 
          phi_update_ack => access_T_CP_0_elements(96), 
          phi_mux_ack => access_T_CP_0_elements(101), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_71_phi_seq_318_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(116);
      access_T_CP_0_elements(121)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(123);
      access_T_CP_0_elements(122)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(124);
      access_T_CP_0_elements(117) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(118);
      access_T_CP_0_elements(125)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(125);
      access_T_CP_0_elements(126)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(127);
      access_T_CP_0_elements(119) <= phi_mux_reqs(1);
      phi_stmt_71_phi_seq_318 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_71_phi_seq_318") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(112), 
          phi_sample_ack => access_T_CP_0_elements(113), 
          phi_update_req => access_T_CP_0_elements(114), 
          phi_update_ack => access_T_CP_0_elements(115), 
          phi_mux_ack => access_T_CP_0_elements(120), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_76_phi_seq_362_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(137);
      access_T_CP_0_elements(140)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(140);
      access_T_CP_0_elements(141)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(142);
      access_T_CP_0_elements(138) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(135);
      access_T_CP_0_elements(144)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(146);
      access_T_CP_0_elements(145)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(147);
      access_T_CP_0_elements(136) <= phi_mux_reqs(1);
      phi_stmt_76_phi_seq_362 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_76_phi_seq_362") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(131), 
          phi_sample_ack => access_T_CP_0_elements(132), 
          phi_update_req => access_T_CP_0_elements(133), 
          phi_update_ack => access_T_CP_0_elements(134), 
          phi_mux_ack => access_T_CP_0_elements(139), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_30_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= access_T_CP_0_elements(7);
        preds(1)  <= access_T_CP_0_elements(8);
        entry_tmerge_30 : transition_merge -- 
          generic map(name => " entry_tmerge_30")
          port map (preds => preds, symbol_out => access_T_CP_0_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u16_u16_125_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_205_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_218_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_231_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_241_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_293_wire : std_logic_vector(15 downto 0);
    signal ADD_u64_u64_278_wire : std_logic_vector(63 downto 0);
    signal AND_u1_u1_107_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_114_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_213_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_227_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_228_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_94_wire : std_logic_vector(0 downto 0);
    signal AND_u32_u32_260_wire : std_logic_vector(31 downto 0);
    signal EQ_u2_u1_103_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_110_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_117_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_90_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_97_wire : std_logic_vector(0 downto 0);
    signal LSHR_u32_u32_274_wire : std_logic_vector(31 downto 0);
    signal MUL_u16_u16_240_wire : std_logic_vector(15 downto 0);
    signal MUL_u16_u16_242_wire : std_logic_vector(15 downto 0);
    signal MUL_u16_u16_30_wire : std_logic_vector(15 downto 0);
    signal MUL_u32_u32_249_wire : std_logic_vector(31 downto 0);
    signal MUX_206_wire : std_logic_vector(15 downto 0);
    signal MUX_219_wire : std_logic_vector(15 downto 0);
    signal MUX_300_wire : std_logic_vector(15 downto 0);
    signal MUX_306_wire : std_logic_vector(15 downto 0);
    signal NEQ_u16_u1_312_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_118_wire : std_logic_vector(0 downto 0);
    signal R_address_132_resized : std_logic_vector(13 downto 0);
    signal R_address_132_scaled : std_logic_vector(13 downto 0);
    signal SUB_u16_u16_286_wire : std_logic_vector(15 downto 0);
    signal SUB_u16_u16_298_wire : std_logic_vector(15 downto 0);
    signal UGT_u16_u1_106_wire : std_logic_vector(0 downto 0);
    signal UGT_u16_u1_113_wire : std_logic_vector(0 downto 0);
    signal UGT_u16_u1_295_wire : std_logic_vector(0 downto 0);
    signal UGT_u16_u1_93_wire : std_logic_vector(0 downto 0);
    signal ULT_u16_u1_303_wire : std_logic_vector(0 downto 0);
    signal ULT_u16_u1_39_wire : std_logic_vector(0 downto 0);
    signal address_46 : std_logic_vector(63 downto 0);
    signal array_obj_ref_133_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_133_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_133_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_133_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_133_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_133_root_address : std_logic_vector(13 downto 0);
    signal c1_156_delayed_14_0_158 : std_logic_vector(0 downto 0);
    signal c1_86 : std_logic_vector(0 downto 0);
    signal c2_160_delayed_14_0_165 : std_logic_vector(0 downto 0);
    signal c2_99 : std_logic_vector(0 downto 0);
    signal c3_120 : std_logic_vector(0 downto 0);
    signal c3_164_delayed_14_0_172 : std_logic_vector(0 downto 0);
    signal c4_128 : std_logic_vector(0 downto 0);
    signal c4_168_delayed_14_0_179 : std_logic_vector(0 downto 0);
    signal col_71 : std_logic_vector(15 downto 0);
    signal col_done_198 : std_logic_vector(0 downto 0);
    signal fetch_addr_135 : std_logic_vector(31 downto 0);
    signal flag1_188 : std_logic_vector(0 downto 0);
    signal fn_blk_43 : std_logic_vector(15 downto 0);
    signal konst_102_wire_constant : std_logic_vector(1 downto 0);
    signal konst_105_wire_constant : std_logic_vector(15 downto 0);
    signal konst_109_wire_constant : std_logic_vector(1 downto 0);
    signal konst_112_wire_constant : std_logic_vector(15 downto 0);
    signal konst_116_wire_constant : std_logic_vector(1 downto 0);
    signal konst_126_wire_constant : std_logic_vector(15 downto 0);
    signal konst_202_wire_constant : std_logic_vector(15 downto 0);
    signal konst_204_wire_constant : std_logic_vector(15 downto 0);
    signal konst_215_wire_constant : std_logic_vector(15 downto 0);
    signal konst_217_wire_constant : std_logic_vector(15 downto 0);
    signal konst_230_wire_constant : std_logic_vector(15 downto 0);
    signal konst_259_wire_constant : std_logic_vector(31 downto 0);
    signal konst_267_wire_constant : std_logic_vector(1 downto 0);
    signal konst_273_wire_constant : std_logic_vector(31 downto 0);
    signal konst_277_wire_constant : std_logic_vector(63 downto 0);
    signal konst_294_wire_constant : std_logic_vector(15 downto 0);
    signal konst_296_wire_constant : std_logic_vector(15 downto 0);
    signal konst_302_wire_constant : std_logic_vector(15 downto 0);
    signal konst_305_wire_constant : std_logic_vector(15 downto 0);
    signal konst_38_wire_constant : std_logic_vector(15 downto 0);
    signal konst_41_wire_constant : std_logic_vector(15 downto 0);
    signal konst_84_wire_constant : std_logic_vector(1 downto 0);
    signal konst_89_wire_constant : std_logic_vector(1 downto 0);
    signal konst_92_wire_constant : std_logic_vector(15 downto 0);
    signal konst_96_wire_constant : std_logic_vector(1 downto 0);
    signal m_factor_32 : std_logic_vector(31 downto 0);
    signal n_address_280 : std_logic_vector(63 downto 0);
    signal n_address_280_50_buffered : std_logic_vector(63 downto 0);
    signal n_blk_308 : std_logic_vector(15 downto 0);
    signal n_blk_308_65_buffered : std_logic_vector(15 downto 0);
    signal n_col_222 : std_logic_vector(15 downto 0);
    signal n_col_222_73_buffered : std_logic_vector(15 downto 0);
    signal n_left_288 : std_logic_vector(15 downto 0);
    signal n_left_288_60_buffered : std_logic_vector(15 downto 0);
    signal n_row_234 : std_logic_vector(15 downto 0);
    signal n_row_234_80_buffered : std_logic_vector(15 downto 0);
    signal n_winr_209 : std_logic_vector(15 downto 0);
    signal n_winr_209_68_buffered : std_logic_vector(15 downto 0);
    signal n_word_start_269 : std_logic_vector(1 downto 0);
    signal n_word_start_269_56_buffered : std_logic_vector(1 downto 0);
    signal na1_244 : std_logic_vector(31 downto 0);
    signal na2_251 : std_logic_vector(31 downto 0);
    signal na3_256 : std_logic_vector(31 downto 0);
    signal na4_262 : std_logic_vector(15 downto 0);
    signal nl_start_35 : std_logic_vector(15 downto 0);
    signal nl_start_35_59_buffered : std_logic_vector(15 downto 0);
    signal num_blk_61 : std_logic_vector(15 downto 0);
    signal num_left_57 : std_logic_vector(15 downto 0);
    signal ptr_deref_138_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_138_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_138_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_138_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_138_word_offset_0 : std_logic_vector(13 downto 0);
    signal row_76 : std_logic_vector(15 downto 0);
    signal type_cast_124_wire : std_logic_vector(15 downto 0);
    signal type_cast_248_wire : std_logic_vector(31 downto 0);
    signal type_cast_266_wire : std_logic_vector(1 downto 0);
    signal type_cast_275_wire : std_logic_vector(63 downto 0);
    signal type_cast_49_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_55_wire_constant : std_logic_vector(1 downto 0);
    signal type_cast_64_wire : std_logic_vector(15 downto 0);
    signal type_cast_70_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_75_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_79_wire_constant : std_logic_vector(15 downto 0);
    signal w1_143 : std_logic_vector(15 downto 0);
    signal w2_147 : std_logic_vector(15 downto 0);
    signal w3_151 : std_logic_vector(15 downto 0);
    signal w4_155 : std_logic_vector(15 downto 0);
    signal winr_66 : std_logic_vector(15 downto 0);
    signal winr_done_193 : std_logic_vector(0 downto 0);
    signal word_read_139 : std_logic_vector(63 downto 0);
    signal word_start_51 : std_logic_vector(1 downto 0);
    -- 
  begin -- 
    array_obj_ref_133_constant_part_of_offset <= "00000000000000";
    array_obj_ref_133_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_133_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_133_resized_base_address <= "00000000000000";
    konst_102_wire_constant <= "00";
    konst_105_wire_constant <= "0000000000000010";
    konst_109_wire_constant <= "01";
    konst_112_wire_constant <= "0000000000000001";
    konst_116_wire_constant <= "10";
    konst_126_wire_constant <= "0000000000000011";
    konst_202_wire_constant <= "0000000000000000";
    konst_204_wire_constant <= "0000000000000001";
    konst_215_wire_constant <= "0000000000000000";
    konst_217_wire_constant <= "0000000000000001";
    konst_230_wire_constant <= "0000000000000001";
    konst_259_wire_constant <= "00000000000000000000000000000011";
    konst_267_wire_constant <= "00";
    konst_273_wire_constant <= "00000000000000000000000000000010";
    konst_277_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    konst_294_wire_constant <= "0000000000000100";
    konst_296_wire_constant <= "0000000000000100";
    konst_302_wire_constant <= "0000000000000100";
    konst_305_wire_constant <= "0000000000000100";
    konst_38_wire_constant <= "0000000000000100";
    konst_41_wire_constant <= "0000000000000100";
    konst_84_wire_constant <= "00";
    konst_89_wire_constant <= "00";
    konst_92_wire_constant <= "0000000000000001";
    konst_96_wire_constant <= "01";
    ptr_deref_138_word_offset_0 <= "00000000000000";
    type_cast_49_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_55_wire_constant <= "00";
    type_cast_70_wire_constant <= "0000000000000000";
    type_cast_75_wire_constant <= "0000000000000000";
    type_cast_79_wire_constant <= "0000000000000000";
    phi_stmt_46: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_49_wire_constant & n_address_280_50_buffered;
      req <= phi_stmt_46_req_0 & phi_stmt_46_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_46",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_46_ack_0,
          idata => idata,
          odata => address_46,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_46
    phi_stmt_51: Block -- phi operator 
      signal idata: std_logic_vector(3 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_55_wire_constant & n_word_start_269_56_buffered;
      req <= phi_stmt_51_req_0 & phi_stmt_51_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_51",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 2) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_51_ack_0,
          idata => idata,
          odata => word_start_51,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_51
    phi_stmt_57: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= nl_start_35_59_buffered & n_left_288_60_buffered;
      req <= phi_stmt_57_req_0 & phi_stmt_57_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_57",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_57_ack_0,
          idata => idata,
          odata => num_left_57,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_57
    phi_stmt_61: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_64_wire & n_blk_308_65_buffered;
      req <= phi_stmt_61_req_0 & phi_stmt_61_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_61",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_61_ack_0,
          idata => idata,
          odata => num_blk_61,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_61
    phi_stmt_66: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= n_winr_209_68_buffered & type_cast_70_wire_constant;
      req <= phi_stmt_66_req_0 & phi_stmt_66_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_66",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_66_ack_0,
          idata => idata,
          odata => winr_66,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_66
    phi_stmt_71: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= n_col_222_73_buffered & type_cast_75_wire_constant;
      req <= phi_stmt_71_req_0 & phi_stmt_71_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_71",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_71_ack_0,
          idata => idata,
          odata => col_71,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_71
    phi_stmt_76: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_79_wire_constant & n_row_234_80_buffered;
      req <= phi_stmt_76_req_0 & phi_stmt_76_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_76",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_76_ack_0,
          idata => idata,
          odata => row_76,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_76
    -- flow-through select operator MUX_206_inst
    MUX_206_wire <= konst_202_wire_constant when (winr_done_193(0) /=  '0') else ADD_u16_u16_205_wire;
    -- flow-through select operator MUX_208_inst
    n_winr_209 <= MUX_206_wire when (flag1_188(0) /=  '0') else winr_66;
    -- flow-through select operator MUX_219_inst
    MUX_219_wire <= konst_215_wire_constant when (col_done_198(0) /=  '0') else ADD_u16_u16_218_wire;
    -- flow-through select operator MUX_221_inst
    n_col_222 <= MUX_219_wire when (AND_u1_u1_213_wire(0) /=  '0') else col_71;
    -- flow-through select operator MUX_233_inst
    n_row_234 <= ADD_u16_u16_231_wire when (AND_u1_u1_228_wire(0) /=  '0') else row_76;
    -- flow-through select operator MUX_268_inst
    n_word_start_269 <= type_cast_266_wire when (flag1_188(0) /=  '0') else konst_267_wire_constant;
    -- flow-through select operator MUX_279_inst
    n_address_280 <= type_cast_275_wire when (flag1_188(0) /=  '0') else ADD_u64_u64_278_wire;
    -- flow-through select operator MUX_287_inst
    n_left_288 <= nl_start_35 when (flag1_188(0) /=  '0') else SUB_u16_u16_286_wire;
    -- flow-through select operator MUX_300_inst
    MUX_300_wire <= SUB_u16_u16_298_wire when (UGT_u16_u1_295_wire(0) /=  '0') else fn_blk_43;
    -- flow-through select operator MUX_306_inst
    MUX_306_wire <= n_left_288 when (ULT_u16_u1_303_wire(0) /=  '0') else konst_305_wire_constant;
    -- flow-through select operator MUX_307_inst
    n_blk_308 <= MUX_300_wire when (flag1_188(0) /=  '0') else MUX_306_wire;
    -- flow-through select operator MUX_42_inst
    fn_blk_43 <= num_cont_buffer when (ULT_u16_u1_39_wire(0) /=  '0') else konst_41_wire_constant;
    slice_142_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_142_inst_req_0;
      slice_142_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_142_inst_req_1;
      slice_142_inst_ack_1<= update_ack(0);
      slice_142_inst: SliceSplitProtocol generic map(name => "slice_142_inst", in_data_width => 64, high_index => 63, low_index => 48, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => word_read_139, dout => w1_143, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_146_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_146_inst_req_0;
      slice_146_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_146_inst_req_1;
      slice_146_inst_ack_1<= update_ack(0);
      slice_146_inst: SliceSplitProtocol generic map(name => "slice_146_inst", in_data_width => 64, high_index => 47, low_index => 32, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => word_read_139, dout => w2_147, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_150_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_150_inst_req_0;
      slice_150_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_150_inst_req_1;
      slice_150_inst_ack_1<= update_ack(0);
      slice_150_inst: SliceSplitProtocol generic map(name => "slice_150_inst", in_data_width => 64, high_index => 31, low_index => 16, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => word_read_139, dout => w3_151, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_154_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_154_inst_req_0;
      slice_154_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_154_inst_req_1;
      slice_154_inst_ack_1<= update_ack(0);
      slice_154_inst: SliceSplitProtocol generic map(name => "slice_154_inst", in_data_width => 64, high_index => 15, low_index => 0, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => word_read_139, dout => w4_155, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    W_c1_156_delayed_14_0_156_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_c1_156_delayed_14_0_156_inst_req_0;
      W_c1_156_delayed_14_0_156_inst_ack_0<= wack(0);
      rreq(0) <= W_c1_156_delayed_14_0_156_inst_req_1;
      W_c1_156_delayed_14_0_156_inst_ack_1<= rack(0);
      W_c1_156_delayed_14_0_156_inst : InterlockBuffer generic map ( -- 
        name => "W_c1_156_delayed_14_0_156_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => c1_86,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => c1_156_delayed_14_0_158,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_c2_160_delayed_14_0_163_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_c2_160_delayed_14_0_163_inst_req_0;
      W_c2_160_delayed_14_0_163_inst_ack_0<= wack(0);
      rreq(0) <= W_c2_160_delayed_14_0_163_inst_req_1;
      W_c2_160_delayed_14_0_163_inst_ack_1<= rack(0);
      W_c2_160_delayed_14_0_163_inst : InterlockBuffer generic map ( -- 
        name => "W_c2_160_delayed_14_0_163_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => c2_99,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => c2_160_delayed_14_0_165,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_c3_164_delayed_14_0_170_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_c3_164_delayed_14_0_170_inst_req_0;
      W_c3_164_delayed_14_0_170_inst_ack_0<= wack(0);
      rreq(0) <= W_c3_164_delayed_14_0_170_inst_req_1;
      W_c3_164_delayed_14_0_170_inst_ack_1<= rack(0);
      W_c3_164_delayed_14_0_170_inst : InterlockBuffer generic map ( -- 
        name => "W_c3_164_delayed_14_0_170_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => c3_120,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => c3_164_delayed_14_0_172,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_c4_168_delayed_14_0_177_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_c4_168_delayed_14_0_177_inst_req_0;
      W_c4_168_delayed_14_0_177_inst_ack_0<= wack(0);
      rreq(0) <= W_c4_168_delayed_14_0_177_inst_req_1;
      W_c4_168_delayed_14_0_177_inst_ack_1<= rack(0);
      W_c4_168_delayed_14_0_177_inst : InterlockBuffer generic map ( -- 
        name => "W_c4_168_delayed_14_0_177_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => c4_128,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => c4_168_delayed_14_0_179,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock W_nl_start_33_inst
    process(num_cont_buffer) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := num_cont_buffer(15 downto 0);
      nl_start_35 <= tmp_var; -- 
    end process;
    addr_of_134_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_134_final_reg_req_0;
      addr_of_134_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_134_final_reg_req_1;
      addr_of_134_final_reg_ack_1<= rack(0);
      addr_of_134_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_134_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_133_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr_135,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_address_280_50_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_address_280_50_buf_req_0;
      n_address_280_50_buf_ack_0<= wack(0);
      rreq(0) <= n_address_280_50_buf_req_1;
      n_address_280_50_buf_ack_1<= rack(0);
      n_address_280_50_buf : InterlockBuffer generic map ( -- 
        name => "n_address_280_50_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_address_280,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_address_280_50_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_blk_308_65_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_blk_308_65_buf_req_0;
      n_blk_308_65_buf_ack_0<= wack(0);
      rreq(0) <= n_blk_308_65_buf_req_1;
      n_blk_308_65_buf_ack_1<= rack(0);
      n_blk_308_65_buf : InterlockBuffer generic map ( -- 
        name => "n_blk_308_65_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_blk_308,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_blk_308_65_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_col_222_73_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_col_222_73_buf_req_0;
      n_col_222_73_buf_ack_0<= wack(0);
      rreq(0) <= n_col_222_73_buf_req_1;
      n_col_222_73_buf_ack_1<= rack(0);
      n_col_222_73_buf : InterlockBuffer generic map ( -- 
        name => "n_col_222_73_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_col_222,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_col_222_73_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_left_288_60_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_left_288_60_buf_req_0;
      n_left_288_60_buf_ack_0<= wack(0);
      rreq(0) <= n_left_288_60_buf_req_1;
      n_left_288_60_buf_ack_1<= rack(0);
      n_left_288_60_buf : InterlockBuffer generic map ( -- 
        name => "n_left_288_60_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_left_288,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_left_288_60_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_row_234_80_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_row_234_80_buf_req_0;
      n_row_234_80_buf_ack_0<= wack(0);
      rreq(0) <= n_row_234_80_buf_req_1;
      n_row_234_80_buf_ack_1<= rack(0);
      n_row_234_80_buf : InterlockBuffer generic map ( -- 
        name => "n_row_234_80_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_row_234,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_row_234_80_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_winr_209_68_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_winr_209_68_buf_req_0;
      n_winr_209_68_buf_ack_0<= wack(0);
      rreq(0) <= n_winr_209_68_buf_req_1;
      n_winr_209_68_buf_ack_1<= rack(0);
      n_winr_209_68_buf : InterlockBuffer generic map ( -- 
        name => "n_winr_209_68_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_winr_209,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_winr_209_68_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_word_start_269_56_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_word_start_269_56_buf_req_0;
      n_word_start_269_56_buf_ack_0<= wack(0);
      rreq(0) <= n_word_start_269_56_buf_req_1;
      n_word_start_269_56_buf_ack_1<= rack(0);
      n_word_start_269_56_buf : InterlockBuffer generic map ( -- 
        name => "n_word_start_269_56_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 2,
        out_data_width => 2,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_word_start_269,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_word_start_269_56_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nl_start_35_59_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nl_start_35_59_buf_req_0;
      nl_start_35_59_buf_ack_0<= wack(0);
      rreq(0) <= nl_start_35_59_buf_req_1;
      nl_start_35_59_buf_ack_1<= rack(0);
      nl_start_35_59_buf : InterlockBuffer generic map ( -- 
        name => "nl_start_35_59_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nl_start_35,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nl_start_35_59_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_124_inst
    process(word_start_51) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 1 downto 0) := word_start_51(1 downto 0);
      type_cast_124_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_243_inst
    process(MUL_u16_u16_242_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := MUL_u16_u16_242_wire(15 downto 0);
      na1_244 <= tmp_var; -- 
    end process;
    -- interlock type_cast_248_inst
    process(n_winr_209) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := n_winr_209(15 downto 0);
      type_cast_248_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_250_inst
    process(MUL_u32_u32_249_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := MUL_u32_u32_249_wire(31 downto 0);
      na2_251 <= tmp_var; -- 
    end process;
    -- interlock type_cast_261_inst
    process(AND_u32_u32_260_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := AND_u32_u32_260_wire(15 downto 0);
      na4_262 <= tmp_var; -- 
    end process;
    -- interlock type_cast_266_inst
    process(na4_262) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 1 downto 0) := na4_262(1 downto 0);
      type_cast_266_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_275_inst
    process(LSHR_u32_u32_274_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := LSHR_u32_u32_274_wire(31 downto 0);
      type_cast_275_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_31_inst
    process(MUL_u16_u16_30_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := MUL_u16_u16_30_wire(15 downto 0);
      m_factor_32 <= tmp_var; -- 
    end process;
    type_cast_64_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_64_inst_req_0;
      type_cast_64_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_64_inst_req_1;
      type_cast_64_inst_ack_1<= rack(0);
      type_cast_64_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_64_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fn_blk_43,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_64_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_133_index_1_rename
    process(R_address_132_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_address_132_resized;
      ov(13 downto 0) := iv;
      R_address_132_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_133_index_1_resize
    process(address_46) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := address_46;
      ov := iv(13 downto 0);
      R_address_132_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_133_root_address_inst
    process(array_obj_ref_133_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_133_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_133_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_138_addr_0
    process(ptr_deref_138_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_138_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_138_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_138_base_resize
    process(fetch_addr_135) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr_135;
      ov := iv(13 downto 0);
      ptr_deref_138_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_138_gather_scatter
    process(ptr_deref_138_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_138_data_0;
      ov(63 downto 0) := iv;
      word_read_139 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_138_root_address_inst
    process(ptr_deref_138_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_138_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_138_root_address <= ov(13 downto 0);
      --
    end process;
    do_while_stmt_44_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NEQ_u16_u1_312_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_44_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_44_branch_req_0,
          ack0 => do_while_stmt_44_branch_ack_0,
          ack1 => do_while_stmt_44_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_125_inst
    process(num_blk_61, type_cast_124_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(num_blk_61, type_cast_124_wire, tmp_var);
      ADD_u16_u16_125_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_205_inst
    process(winr_66) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(winr_66, konst_204_wire_constant, tmp_var);
      ADD_u16_u16_205_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_218_inst
    process(col_71) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(col_71, konst_217_wire_constant, tmp_var);
      ADD_u16_u16_218_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_231_inst
    process(row_76) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(row_76, konst_230_wire_constant, tmp_var);
      ADD_u16_u16_231_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_241_inst
    process(n_col_222, MUL_u16_u16_240_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(n_col_222, MUL_u16_u16_240_wire, tmp_var);
      ADD_u16_u16_241_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_293_inst
    process(fn_blk_43, na4_262) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(fn_blk_43, na4_262, tmp_var);
      ADD_u16_u16_293_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_255_inst
    process(na1_244, na2_251) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(na1_244, na2_251, tmp_var);
      na3_256 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_278_inst
    process(address_46) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(address_46, konst_277_wire_constant, tmp_var);
      ADD_u64_u64_278_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_107_inst
    process(EQ_u2_u1_103_wire, UGT_u16_u1_106_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u2_u1_103_wire, UGT_u16_u1_106_wire, tmp_var);
      AND_u1_u1_107_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_114_inst
    process(EQ_u2_u1_110_wire, UGT_u16_u1_113_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u2_u1_110_wire, UGT_u16_u1_113_wire, tmp_var);
      AND_u1_u1_114_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_213_inst
    process(winr_done_193, flag1_188) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(winr_done_193, flag1_188, tmp_var);
      AND_u1_u1_213_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_227_inst
    process(col_done_198, flag1_188) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(col_done_198, flag1_188, tmp_var);
      AND_u1_u1_227_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_228_inst
    process(winr_done_193, AND_u1_u1_227_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(winr_done_193, AND_u1_u1_227_wire, tmp_var);
      AND_u1_u1_228_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_94_inst
    process(EQ_u2_u1_90_wire, UGT_u16_u1_93_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u2_u1_90_wire, UGT_u16_u1_93_wire, tmp_var);
      AND_u1_u1_94_wire <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_260_inst
    process(na3_256) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(na3_256, konst_259_wire_constant, tmp_var);
      AND_u32_u32_260_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_187_inst
    process(num_left_57, num_blk_61) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(num_left_57, num_blk_61, tmp_var);
      flag1_188 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_192_inst
    process(winr_66, rk1_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(winr_66, rk1_buffer, tmp_var);
      winr_done_193 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_197_inst
    process(col_71, col1_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(col_71, col1_buffer, tmp_var);
      col_done_198 <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_103_inst
    process(word_start_51) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(word_start_51, konst_102_wire_constant, tmp_var);
      EQ_u2_u1_103_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_110_inst
    process(word_start_51) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(word_start_51, konst_109_wire_constant, tmp_var);
      EQ_u2_u1_110_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_117_inst
    process(word_start_51) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(word_start_51, konst_116_wire_constant, tmp_var);
      EQ_u2_u1_117_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_85_inst
    process(word_start_51) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(word_start_51, konst_84_wire_constant, tmp_var);
      c1_86 <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_90_inst
    process(word_start_51) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(word_start_51, konst_89_wire_constant, tmp_var);
      EQ_u2_u1_90_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_97_inst
    process(word_start_51) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(word_start_51, konst_96_wire_constant, tmp_var);
      EQ_u2_u1_97_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_274_inst
    process(na3_256) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(na3_256, konst_273_wire_constant, tmp_var);
      LSHR_u32_u32_274_wire <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_240_inst
    process(ct_buffer, n_row_234) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(ct_buffer, n_row_234, tmp_var);
      MUL_u16_u16_240_wire <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_242_inst
    process(chl_in_buffer, ADD_u16_u16_241_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(chl_in_buffer, ADD_u16_u16_241_wire, tmp_var);
      MUL_u16_u16_242_wire <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_30_inst
    process(ct_buffer, chl_in_buffer) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(ct_buffer, chl_in_buffer, tmp_var);
      MUL_u16_u16_30_wire <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_249_inst
    process(m_factor_32, type_cast_248_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(m_factor_32, type_cast_248_wire, tmp_var);
      MUL_u32_u32_249_wire <= tmp_var; --
    end process;
    -- binary operator NEQ_u16_u1_312_inst
    process(n_row_234, row1_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntNe_proc(n_row_234, row1_buffer, tmp_var);
      NEQ_u16_u1_312_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_118_inst
    process(AND_u1_u1_114_wire, EQ_u2_u1_117_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(AND_u1_u1_114_wire, EQ_u2_u1_117_wire, tmp_var);
      OR_u1_u1_118_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_119_inst
    process(AND_u1_u1_107_wire, OR_u1_u1_118_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(AND_u1_u1_107_wire, OR_u1_u1_118_wire, tmp_var);
      c3_120 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_98_inst
    process(AND_u1_u1_94_wire, EQ_u2_u1_97_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(AND_u1_u1_94_wire, EQ_u2_u1_97_wire, tmp_var);
      c2_99 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_286_inst
    process(num_left_57, num_blk_61) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(num_left_57, num_blk_61, tmp_var);
      SUB_u16_u16_286_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_298_inst
    process(konst_296_wire_constant, na4_262) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(konst_296_wire_constant, na4_262, tmp_var);
      SUB_u16_u16_298_wire <= tmp_var; --
    end process;
    -- binary operator UGT_u16_u1_106_inst
    process(num_blk_61) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(num_blk_61, konst_105_wire_constant, tmp_var);
      UGT_u16_u1_106_wire <= tmp_var; --
    end process;
    -- binary operator UGT_u16_u1_113_inst
    process(num_blk_61) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(num_blk_61, konst_112_wire_constant, tmp_var);
      UGT_u16_u1_113_wire <= tmp_var; --
    end process;
    -- binary operator UGT_u16_u1_127_inst
    process(ADD_u16_u16_125_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(ADD_u16_u16_125_wire, konst_126_wire_constant, tmp_var);
      c4_128 <= tmp_var; --
    end process;
    -- binary operator UGT_u16_u1_295_inst
    process(ADD_u16_u16_293_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(ADD_u16_u16_293_wire, konst_294_wire_constant, tmp_var);
      UGT_u16_u1_295_wire <= tmp_var; --
    end process;
    -- binary operator UGT_u16_u1_93_inst
    process(num_blk_61) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(num_blk_61, konst_92_wire_constant, tmp_var);
      UGT_u16_u1_93_wire <= tmp_var; --
    end process;
    -- binary operator ULT_u16_u1_303_inst
    process(n_left_288) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(n_left_288, konst_302_wire_constant, tmp_var);
      ULT_u16_u1_303_wire <= tmp_var; --
    end process;
    -- binary operator ULT_u16_u1_39_inst
    process(num_cont_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(num_cont_buffer, konst_38_wire_constant, tmp_var);
      ULT_u16_u1_39_wire <= tmp_var; --
    end process;
    -- shared split operator group (42) : array_obj_ref_133_index_offset 
    ApIntAdd_group_42: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_address_132_scaled;
      array_obj_ref_133_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_133_index_offset_req_0;
      array_obj_ref_133_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_133_index_offset_req_1;
      array_obj_ref_133_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_42_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_42_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_42",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 42
    -- shared load operator group (0) : ptr_deref_138_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 6);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_138_load_0_req_0;
      ptr_deref_138_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_138_load_0_req_1;
      ptr_deref_138_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_138_word_address_0;
      ptr_deref_138_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared outport operator group (0) : WPIPE_input_pipe1_174_inst WPIPE_input_pipe1_167_inst WPIPE_input_pipe1_160_inst WPIPE_input_pipe1_181_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 3 downto 0);
      signal update_req, update_ack : BooleanArray( 3 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 3 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 3 downto 0);
      signal guard_vector : std_logic_vector( 3 downto 0);
      constant inBUFs : IntegerArray(3 downto 0) := (3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(3 downto 0) := (0 => true, 1 => true, 2 => true, 3 => true);
      constant guardBuffering: IntegerArray(3 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2);
      -- 
    begin -- 
      sample_req_unguarded(3) <= WPIPE_input_pipe1_174_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_input_pipe1_167_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_input_pipe1_160_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_input_pipe1_181_inst_req_0;
      WPIPE_input_pipe1_174_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_input_pipe1_167_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_input_pipe1_160_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_input_pipe1_181_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(3) <= WPIPE_input_pipe1_174_inst_req_1;
      update_req_unguarded(2) <= WPIPE_input_pipe1_167_inst_req_1;
      update_req_unguarded(1) <= WPIPE_input_pipe1_160_inst_req_1;
      update_req_unguarded(0) <= WPIPE_input_pipe1_181_inst_req_1;
      WPIPE_input_pipe1_174_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_input_pipe1_167_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_input_pipe1_160_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_input_pipe1_181_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= c4_168_delayed_14_0_179(0);
      guard_vector(1)  <= c1_156_delayed_14_0_158(0);
      guard_vector(2)  <= c2_160_delayed_14_0_165(0);
      guard_vector(3)  <= c3_164_delayed_14_0_172(0);
      data_in <= w3_151 & w2_147 & w1_143 & w4_155;
      input_pipe1_write_0_gI: SplitGuardInterface generic map(name => "input_pipe1_write_0_gI", nreqs => 4, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      input_pipe1_write_0: OutputPortRevised -- 
        generic map ( name => "input_pipe1", data_width => 16, num_reqs => 4, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => input_pipe1_pipe_write_req(0),
          oack => input_pipe1_pipe_write_ack(0),
          odata => input_pipe1_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end access_T_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convolution3D is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(1 downto 0);
    maxpool_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    elapsed_time_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_write_data : out  std_logic_vector(63 downto 0);
    maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    num_out_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    num_out_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    num_out_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
    access_T_call_reqs : out  std_logic_vector(0 downto 0);
    access_T_call_acks : in   std_logic_vector(0 downto 0);
    access_T_call_data : out  std_logic_vector(95 downto 0);
    access_T_call_tag  :  out  std_logic_vector(0 downto 0);
    access_T_return_reqs : out  std_logic_vector(0 downto 0);
    access_T_return_acks : in   std_logic_vector(0 downto 0);
    access_T_return_tag :  in   std_logic_vector(0 downto 0);
    timer_call_reqs : out  std_logic_vector(0 downto 0);
    timer_call_acks : in   std_logic_vector(0 downto 0);
    timer_call_tag  :  out  std_logic_vector(1 downto 0);
    timer_return_reqs : out  std_logic_vector(0 downto 0);
    timer_return_acks : in   std_logic_vector(0 downto 0);
    timer_return_data : in   std_logic_vector(63 downto 0);
    timer_return_tag :  in   std_logic_vector(1 downto 0);
    loadKernelChannel_call_reqs : out  std_logic_vector(0 downto 0);
    loadKernelChannel_call_acks : in   std_logic_vector(0 downto 0);
    loadKernelChannel_call_data : out  std_logic_vector(127 downto 0);
    loadKernelChannel_call_tag  :  out  std_logic_vector(0 downto 0);
    loadKernelChannel_return_reqs : out  std_logic_vector(0 downto 0);
    loadKernelChannel_return_acks : in   std_logic_vector(0 downto 0);
    loadKernelChannel_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convolution3D;
architecture convolution3D_arch of convolution3D is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convolution3D_CP_1120_start: Boolean;
  signal convolution3D_CP_1120_symbol: Boolean;
  -- volatile/operator module components. 
  component access_T is -- 
    generic (tag_length : integer); 
    port ( -- 
      num_cont : in  std_logic_vector(15 downto 0);
      row1 : in  std_logic_vector(15 downto 0);
      col1 : in  std_logic_vector(15 downto 0);
      rk1 : in  std_logic_vector(15 downto 0);
      chl_in : in  std_logic_vector(15 downto 0);
      ct : in  std_logic_vector(15 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
      input_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      c : out  std_logic_vector(63 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component loadKernelChannel is -- 
    generic (tag_length : integer); 
    port ( -- 
      start_add : in  std_logic_vector(63 downto 0);
      end_add : in  std_logic_vector(63 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
      input_done_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_data : in   std_logic_vector(0 downto 0);
      size_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      size_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      size_pipe_pipe_write_data : out  std_logic_vector(31 downto 0);
      kernel_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal WPIPE_maxpool_output_pipe_611_inst_req_1 : boolean;
  signal type_cast_616_inst_ack_0 : boolean;
  signal type_cast_569_inst_ack_1 : boolean;
  signal type_cast_492_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_564_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_593_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_593_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_518_inst_ack_0 : boolean;
  signal type_cast_492_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_609_inst_ack_1 : boolean;
  signal type_cast_600_inst_ack_0 : boolean;
  signal type_cast_600_inst_req_1 : boolean;
  signal type_cast_569_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_518_inst_req_0 : boolean;
  signal type_cast_569_inst_req_0 : boolean;
  signal type_cast_492_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_580_inst_req_0 : boolean;
  signal type_cast_600_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_531_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_531_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_533_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_547_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_593_inst_req_1 : boolean;
  signal type_cast_1102_inst_ack_1 : boolean;
  signal type_cast_1159_inst_ack_1 : boolean;
  signal type_cast_1159_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_564_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_564_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_531_inst_req_1 : boolean;
  signal type_cast_554_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_611_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_593_inst_ack_0 : boolean;
  signal type_cast_538_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_516_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_533_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_502_inst_ack_1 : boolean;
  signal type_cast_554_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_533_inst_ack_1 : boolean;
  signal type_cast_554_inst_req_0 : boolean;
  signal type_cast_1159_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_516_inst_req_1 : boolean;
  signal type_cast_523_inst_ack_0 : boolean;
  signal type_cast_554_inst_req_1 : boolean;
  signal type_cast_538_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_533_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_516_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_562_inst_ack_1 : boolean;
  signal type_cast_569_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_562_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_549_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_578_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_516_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_502_inst_req_1 : boolean;
  signal type_cast_507_inst_ack_1 : boolean;
  signal type_cast_492_inst_ack_1 : boolean;
  signal type_cast_600_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_609_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_580_inst_ack_1 : boolean;
  signal type_cast_616_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_487_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_487_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_930_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_564_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_562_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_549_inst_ack_0 : boolean;
  signal type_cast_538_inst_req_1 : boolean;
  signal type_cast_523_inst_req_0 : boolean;
  signal type_cast_538_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_500_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_531_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_562_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_500_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_609_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_580_inst_ack_0 : boolean;
  signal type_cast_585_inst_req_0 : boolean;
  signal type_cast_585_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_518_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_518_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_500_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_500_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_951_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_611_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_626_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_626_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_609_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_595_inst_ack_1 : boolean;
  signal type_cast_631_inst_ack_1 : boolean;
  signal type_cast_616_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_626_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_626_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_951_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_580_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_578_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_595_inst_req_1 : boolean;
  signal type_cast_616_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_640_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_640_inst_ack_0 : boolean;
  signal type_cast_1163_inst_ack_1 : boolean;
  signal type_cast_1171_inst_req_1 : boolean;
  signal call_stmt_1761_call_ack_0 : boolean;
  signal type_cast_1163_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_547_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_595_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_549_inst_ack_1 : boolean;
  signal type_cast_1159_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_624_inst_ack_1 : boolean;
  signal type_cast_631_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_502_inst_ack_0 : boolean;
  signal type_cast_631_inst_ack_0 : boolean;
  signal type_cast_631_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_502_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_624_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_624_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_611_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_640_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_640_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_624_inst_ack_0 : boolean;
  signal type_cast_1102_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_547_inst_req_1 : boolean;
  signal type_cast_507_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_595_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_578_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_930_inst_ack_1 : boolean;
  signal type_cast_523_inst_ack_1 : boolean;
  signal type_cast_585_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_578_inst_req_0 : boolean;
  signal type_cast_523_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_549_inst_req_1 : boolean;
  signal type_cast_507_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_547_inst_ack_0 : boolean;
  signal type_cast_507_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_932_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_953_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_932_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_932_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_932_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_953_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_951_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_438_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_438_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_438_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_438_inst_ack_1 : boolean;
  signal ptr_deref_966_store_0_req_0 : boolean;
  signal ptr_deref_966_store_0_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_440_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_440_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_440_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_440_inst_ack_1 : boolean;
  signal array_obj_ref_1148_index_offset_req_0 : boolean;
  signal type_cast_445_inst_req_0 : boolean;
  signal type_cast_445_inst_ack_0 : boolean;
  signal type_cast_445_inst_req_1 : boolean;
  signal type_cast_445_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_454_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_454_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_454_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_454_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_456_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_456_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_456_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_456_inst_ack_1 : boolean;
  signal type_cast_585_inst_req_1 : boolean;
  signal type_cast_461_inst_req_0 : boolean;
  signal type_cast_461_inst_ack_0 : boolean;
  signal type_cast_461_inst_req_1 : boolean;
  signal type_cast_461_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_469_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_469_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_469_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_469_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_471_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_471_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_471_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_471_inst_ack_1 : boolean;
  signal type_cast_476_inst_req_0 : boolean;
  signal type_cast_476_inst_ack_0 : boolean;
  signal type_cast_476_inst_req_1 : boolean;
  signal type_cast_476_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_485_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_485_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_485_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_485_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_487_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_487_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1080_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_642_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1080_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_642_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_642_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_642_inst_ack_1 : boolean;
  signal type_cast_1102_inst_ack_0 : boolean;
  signal type_cast_1102_inst_req_0 : boolean;
  signal array_obj_ref_1148_index_offset_ack_1 : boolean;
  signal type_cast_647_inst_req_0 : boolean;
  signal type_cast_647_inst_ack_0 : boolean;
  signal type_cast_647_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1080_inst_ack_0 : boolean;
  signal type_cast_647_inst_ack_1 : boolean;
  signal array_obj_ref_1648_index_offset_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_655_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1080_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_655_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_655_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_951_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_655_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_657_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_657_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_657_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_657_inst_ack_1 : boolean;
  signal array_obj_ref_1148_index_offset_req_1 : boolean;
  signal type_cast_662_inst_req_0 : boolean;
  signal type_cast_662_inst_ack_0 : boolean;
  signal type_cast_662_inst_req_1 : boolean;
  signal type_cast_662_inst_ack_1 : boolean;
  signal type_cast_1167_inst_ack_1 : boolean;
  signal type_cast_1163_inst_ack_0 : boolean;
  signal type_cast_1163_inst_req_0 : boolean;
  signal if_stmt_1109_branch_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_671_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_671_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_671_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_671_inst_ack_1 : boolean;
  signal type_cast_1167_inst_ack_0 : boolean;
  signal if_stmt_1109_branch_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_673_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_673_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_673_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_673_inst_ack_1 : boolean;
  signal type_cast_1087_inst_ack_1 : boolean;
  signal type_cast_678_inst_req_0 : boolean;
  signal type_cast_678_inst_ack_0 : boolean;
  signal type_cast_678_inst_req_1 : boolean;
  signal type_cast_678_inst_ack_1 : boolean;
  signal type_cast_1167_inst_req_1 : boolean;
  signal type_cast_1171_inst_ack_0 : boolean;
  signal type_cast_1087_inst_req_1 : boolean;
  signal type_cast_1087_inst_ack_0 : boolean;
  signal type_cast_687_inst_req_0 : boolean;
  signal if_stmt_1031_branch_ack_0 : boolean;
  signal type_cast_687_inst_ack_0 : boolean;
  signal ptr_deref_966_store_0_ack_1 : boolean;
  signal type_cast_687_inst_req_1 : boolean;
  signal type_cast_687_inst_ack_1 : boolean;
  signal type_cast_1171_inst_ack_1 : boolean;
  signal type_cast_1087_inst_req_0 : boolean;
  signal type_cast_691_inst_req_0 : boolean;
  signal if_stmt_1031_branch_ack_1 : boolean;
  signal type_cast_691_inst_ack_0 : boolean;
  signal type_cast_691_inst_req_1 : boolean;
  signal type_cast_691_inst_ack_1 : boolean;
  signal ptr_deref_1152_store_0_ack_1 : boolean;
  signal type_cast_707_inst_req_0 : boolean;
  signal if_stmt_1031_branch_req_0 : boolean;
  signal type_cast_707_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_930_inst_ack_0 : boolean;
  signal type_cast_707_inst_req_1 : boolean;
  signal type_cast_707_inst_ack_1 : boolean;
  signal type_cast_937_inst_ack_1 : boolean;
  signal ptr_deref_1152_store_0_req_1 : boolean;
  signal ptr_deref_1152_store_0_ack_0 : boolean;
  signal ptr_deref_1152_store_0_req_0 : boolean;
  signal type_cast_937_inst_req_1 : boolean;
  signal ptr_deref_966_store_0_req_1 : boolean;
  signal if_stmt_715_branch_req_0 : boolean;
  signal if_stmt_715_branch_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_930_inst_req_0 : boolean;
  signal if_stmt_715_branch_ack_0 : boolean;
  signal addr_of_1149_final_reg_ack_1 : boolean;
  signal type_cast_735_inst_req_0 : boolean;
  signal type_cast_735_inst_ack_0 : boolean;
  signal addr_of_1149_final_reg_req_1 : boolean;
  signal type_cast_735_inst_req_1 : boolean;
  signal type_cast_735_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1082_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1082_inst_req_1 : boolean;
  signal if_stmt_1109_branch_req_0 : boolean;
  signal type_cast_751_inst_req_0 : boolean;
  signal type_cast_751_inst_ack_0 : boolean;
  signal type_cast_751_inst_req_1 : boolean;
  signal type_cast_751_inst_ack_1 : boolean;
  signal type_cast_937_inst_ack_0 : boolean;
  signal type_cast_937_inst_req_0 : boolean;
  signal type_cast_958_inst_ack_1 : boolean;
  signal addr_of_1149_final_reg_ack_0 : boolean;
  signal type_cast_760_inst_req_0 : boolean;
  signal type_cast_760_inst_ack_0 : boolean;
  signal addr_of_1149_final_reg_req_0 : boolean;
  signal type_cast_760_inst_req_1 : boolean;
  signal type_cast_760_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1082_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1082_inst_req_0 : boolean;
  signal type_cast_958_inst_req_1 : boolean;
  signal type_cast_958_inst_ack_0 : boolean;
  signal type_cast_770_inst_req_0 : boolean;
  signal if_stmt_980_branch_ack_0 : boolean;
  signal type_cast_770_inst_ack_0 : boolean;
  signal type_cast_770_inst_req_1 : boolean;
  signal type_cast_770_inst_ack_1 : boolean;
  signal type_cast_958_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_953_inst_ack_1 : boolean;
  signal type_cast_1167_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_953_inst_req_1 : boolean;
  signal array_obj_ref_805_index_offset_req_0 : boolean;
  signal if_stmt_980_branch_ack_1 : boolean;
  signal array_obj_ref_805_index_offset_ack_0 : boolean;
  signal array_obj_ref_805_index_offset_req_1 : boolean;
  signal array_obj_ref_805_index_offset_ack_1 : boolean;
  signal array_obj_ref_1148_index_offset_ack_0 : boolean;
  signal if_stmt_980_branch_req_0 : boolean;
  signal addr_of_806_final_reg_req_0 : boolean;
  signal addr_of_806_final_reg_ack_0 : boolean;
  signal addr_of_806_final_reg_req_1 : boolean;
  signal addr_of_806_final_reg_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_809_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_809_inst_ack_0 : boolean;
  signal ptr_deref_1652_store_0_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_809_inst_req_1 : boolean;
  signal ptr_deref_1652_store_0_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_809_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_811_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_811_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_811_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_811_inst_ack_1 : boolean;
  signal type_cast_1698_inst_req_0 : boolean;
  signal type_cast_816_inst_req_0 : boolean;
  signal type_cast_816_inst_ack_0 : boolean;
  signal type_cast_816_inst_req_1 : boolean;
  signal type_cast_816_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_825_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_825_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_825_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_825_inst_ack_1 : boolean;
  signal type_cast_1698_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_827_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_827_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_827_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_827_inst_ack_1 : boolean;
  signal type_cast_832_inst_req_0 : boolean;
  signal type_cast_832_inst_ack_0 : boolean;
  signal type_cast_832_inst_req_1 : boolean;
  signal type_cast_832_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1580_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_846_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_846_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_846_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_846_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1580_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_848_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_848_inst_ack_0 : boolean;
  signal type_cast_1171_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_848_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_848_inst_ack_1 : boolean;
  signal type_cast_1698_inst_req_1 : boolean;
  signal type_cast_1746_inst_req_0 : boolean;
  signal type_cast_853_inst_req_0 : boolean;
  signal type_cast_853_inst_ack_0 : boolean;
  signal type_cast_853_inst_req_1 : boolean;
  signal type_cast_853_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1580_inst_req_1 : boolean;
  signal type_cast_1698_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_867_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_867_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1580_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_867_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_867_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_869_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_869_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_869_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_869_inst_ack_1 : boolean;
  signal type_cast_874_inst_req_0 : boolean;
  signal type_cast_874_inst_ack_0 : boolean;
  signal type_cast_874_inst_req_1 : boolean;
  signal type_cast_874_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_888_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_888_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_888_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_888_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_890_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_890_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_890_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_890_inst_ack_1 : boolean;
  signal type_cast_895_inst_req_0 : boolean;
  signal type_cast_895_inst_ack_0 : boolean;
  signal type_cast_895_inst_req_1 : boolean;
  signal type_cast_895_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_909_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_909_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_909_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_909_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_911_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_911_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_911_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_911_inst_ack_1 : boolean;
  signal type_cast_916_inst_req_0 : boolean;
  signal type_cast_916_inst_ack_0 : boolean;
  signal type_cast_916_inst_req_1 : boolean;
  signal type_cast_916_inst_ack_1 : boolean;
  signal call_stmt_1754_call_req_1 : boolean;
  signal call_stmt_1761_call_req_1 : boolean;
  signal array_obj_ref_1648_index_offset_req_0 : boolean;
  signal if_stmt_1209_branch_req_0 : boolean;
  signal if_stmt_1476_branch_ack_0 : boolean;
  signal if_stmt_1209_branch_ack_1 : boolean;
  signal if_stmt_1209_branch_ack_0 : boolean;
  signal type_cast_1708_inst_ack_0 : boolean;
  signal type_cast_1230_inst_req_0 : boolean;
  signal type_cast_1230_inst_ack_0 : boolean;
  signal type_cast_1230_inst_req_1 : boolean;
  signal type_cast_1230_inst_ack_1 : boolean;
  signal call_stmt_1761_call_req_0 : boolean;
  signal call_stmt_1761_call_ack_1 : boolean;
  signal call_stmt_1659_call_ack_1 : boolean;
  signal call_stmt_1659_call_req_1 : boolean;
  signal type_cast_1717_inst_ack_1 : boolean;
  signal type_cast_1234_inst_req_0 : boolean;
  signal type_cast_1234_inst_ack_0 : boolean;
  signal type_cast_1717_inst_req_1 : boolean;
  signal type_cast_1234_inst_req_1 : boolean;
  signal type_cast_1234_inst_ack_1 : boolean;
  signal call_stmt_1754_call_ack_0 : boolean;
  signal call_stmt_1754_call_req_0 : boolean;
  signal type_cast_1243_inst_req_0 : boolean;
  signal type_cast_1243_inst_ack_0 : boolean;
  signal type_cast_1243_inst_req_1 : boolean;
  signal type_cast_1243_inst_ack_1 : boolean;
  signal if_stmt_1476_branch_ack_1 : boolean;
  signal type_cast_1252_inst_req_0 : boolean;
  signal type_cast_1252_inst_ack_0 : boolean;
  signal type_cast_1252_inst_req_1 : boolean;
  signal type_cast_1252_inst_ack_1 : boolean;
  signal call_stmt_1659_call_ack_0 : boolean;
  signal call_stmt_1659_call_req_0 : boolean;
  signal if_stmt_1609_branch_ack_0 : boolean;
  signal if_stmt_1609_branch_ack_1 : boolean;
  signal type_cast_1717_inst_ack_0 : boolean;
  signal type_cast_1261_inst_req_0 : boolean;
  signal type_cast_1261_inst_ack_0 : boolean;
  signal type_cast_1717_inst_req_0 : boolean;
  signal type_cast_1261_inst_req_1 : boolean;
  signal type_cast_1261_inst_ack_1 : boolean;
  signal type_cast_1542_inst_ack_1 : boolean;
  signal type_cast_1542_inst_req_1 : boolean;
  signal if_stmt_1609_branch_req_0 : boolean;
  signal type_cast_1266_inst_req_0 : boolean;
  signal type_cast_1266_inst_ack_0 : boolean;
  signal type_cast_1266_inst_req_1 : boolean;
  signal type_cast_1266_inst_ack_1 : boolean;
  signal type_cast_1708_inst_req_0 : boolean;
  signal type_cast_1602_inst_ack_1 : boolean;
  signal type_cast_1602_inst_req_1 : boolean;
  signal type_cast_1750_inst_ack_1 : boolean;
  signal type_cast_1602_inst_ack_0 : boolean;
  signal array_obj_ref_1301_index_offset_req_0 : boolean;
  signal array_obj_ref_1301_index_offset_ack_0 : boolean;
  signal type_cast_1542_inst_ack_0 : boolean;
  signal array_obj_ref_1301_index_offset_req_1 : boolean;
  signal array_obj_ref_1301_index_offset_ack_1 : boolean;
  signal type_cast_1750_inst_req_1 : boolean;
  signal type_cast_1602_inst_req_0 : boolean;
  signal type_cast_1542_inst_req_0 : boolean;
  signal addr_of_1302_final_reg_req_0 : boolean;
  signal addr_of_1302_final_reg_ack_0 : boolean;
  signal addr_of_1302_final_reg_req_1 : boolean;
  signal addr_of_1302_final_reg_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1305_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1305_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1305_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1305_inst_ack_1 : boolean;
  signal type_cast_1750_inst_ack_0 : boolean;
  signal type_cast_1750_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1674_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1674_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1307_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1307_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1307_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1307_inst_ack_1 : boolean;
  signal type_cast_1587_inst_ack_1 : boolean;
  signal type_cast_1587_inst_req_1 : boolean;
  signal type_cast_1312_inst_req_0 : boolean;
  signal type_cast_1312_inst_ack_0 : boolean;
  signal type_cast_1312_inst_req_1 : boolean;
  signal type_cast_1312_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1674_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1321_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1321_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1321_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1321_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1674_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1323_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1323_inst_ack_0 : boolean;
  signal if_stmt_1527_branch_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1323_inst_req_1 : boolean;
  signal addr_of_1649_final_reg_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1323_inst_ack_1 : boolean;
  signal call_stmt_1754_call_ack_1 : boolean;
  signal type_cast_1587_inst_ack_0 : boolean;
  signal type_cast_1587_inst_req_0 : boolean;
  signal type_cast_1708_inst_ack_1 : boolean;
  signal type_cast_1328_inst_req_0 : boolean;
  signal addr_of_1649_final_reg_req_1 : boolean;
  signal type_cast_1328_inst_ack_0 : boolean;
  signal type_cast_1708_inst_req_1 : boolean;
  signal type_cast_1328_inst_req_1 : boolean;
  signal type_cast_1328_inst_ack_1 : boolean;
  signal if_stmt_1527_branch_ack_1 : boolean;
  signal ptr_deref_1652_store_0_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1342_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1342_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1342_inst_req_1 : boolean;
  signal addr_of_1649_final_reg_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1342_inst_ack_1 : boolean;
  signal WPIPE_num_out_pipe_1671_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1344_inst_req_0 : boolean;
  signal addr_of_1649_final_reg_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1344_inst_ack_0 : boolean;
  signal type_cast_1746_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1344_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1344_inst_ack_1 : boolean;
  signal type_cast_1746_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1582_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1582_inst_req_1 : boolean;
  signal type_cast_1349_inst_req_0 : boolean;
  signal type_cast_1349_inst_ack_0 : boolean;
  signal type_cast_1349_inst_req_1 : boolean;
  signal type_cast_1349_inst_ack_1 : boolean;
  signal if_stmt_1527_branch_req_0 : boolean;
  signal ptr_deref_1652_store_0_req_1 : boolean;
  signal WPIPE_num_out_pipe_1671_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1363_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1363_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1363_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1363_inst_ack_1 : boolean;
  signal WPIPE_num_out_pipe_1671_inst_ack_0 : boolean;
  signal WPIPE_num_out_pipe_1671_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1365_inst_req_0 : boolean;
  signal array_obj_ref_1648_index_offset_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1365_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1365_inst_req_1 : boolean;
  signal array_obj_ref_1648_index_offset_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1365_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1582_inst_ack_0 : boolean;
  signal type_cast_1746_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1582_inst_req_0 : boolean;
  signal type_cast_1370_inst_req_0 : boolean;
  signal type_cast_1370_inst_ack_0 : boolean;
  signal if_stmt_1476_branch_req_0 : boolean;
  signal type_cast_1370_inst_req_1 : boolean;
  signal type_cast_1370_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1384_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1384_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1384_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1384_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1386_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1386_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1386_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1386_inst_ack_1 : boolean;
  signal type_cast_1391_inst_req_0 : boolean;
  signal type_cast_1391_inst_ack_0 : boolean;
  signal type_cast_1391_inst_req_1 : boolean;
  signal type_cast_1391_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1405_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1405_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1405_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1405_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1407_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1407_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1407_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1407_inst_ack_1 : boolean;
  signal type_cast_1412_inst_req_0 : boolean;
  signal type_cast_1412_inst_ack_0 : boolean;
  signal type_cast_1412_inst_req_1 : boolean;
  signal type_cast_1412_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1426_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1426_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1426_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1426_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1428_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1428_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1428_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1428_inst_ack_1 : boolean;
  signal type_cast_1433_inst_req_0 : boolean;
  signal type_cast_1433_inst_ack_0 : boolean;
  signal type_cast_1433_inst_req_1 : boolean;
  signal type_cast_1433_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1447_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1447_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1447_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1447_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1449_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1449_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1449_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1449_inst_ack_1 : boolean;
  signal type_cast_1454_inst_req_0 : boolean;
  signal type_cast_1454_inst_ack_0 : boolean;
  signal type_cast_1454_inst_req_1 : boolean;
  signal type_cast_1454_inst_ack_1 : boolean;
  signal ptr_deref_1462_store_0_req_0 : boolean;
  signal ptr_deref_1462_store_0_ack_0 : boolean;
  signal ptr_deref_1462_store_0_req_1 : boolean;
  signal ptr_deref_1462_store_0_ack_1 : boolean;
  signal if_stmt_1773_branch_req_0 : boolean;
  signal if_stmt_1773_branch_ack_1 : boolean;
  signal if_stmt_1773_branch_ack_0 : boolean;
  signal type_cast_1783_inst_req_0 : boolean;
  signal type_cast_1783_inst_ack_0 : boolean;
  signal type_cast_1783_inst_req_1 : boolean;
  signal type_cast_1783_inst_ack_1 : boolean;
  signal call_stmt_1787_call_req_0 : boolean;
  signal call_stmt_1787_call_ack_0 : boolean;
  signal call_stmt_1787_call_req_1 : boolean;
  signal call_stmt_1787_call_ack_1 : boolean;
  signal type_cast_1791_inst_req_0 : boolean;
  signal type_cast_1791_inst_ack_0 : boolean;
  signal type_cast_1791_inst_req_1 : boolean;
  signal type_cast_1791_inst_ack_1 : boolean;
  signal WPIPE_elapsed_time_pipe_1798_inst_req_0 : boolean;
  signal WPIPE_elapsed_time_pipe_1798_inst_ack_0 : boolean;
  signal WPIPE_elapsed_time_pipe_1798_inst_req_1 : boolean;
  signal WPIPE_elapsed_time_pipe_1798_inst_ack_1 : boolean;
  signal phi_stmt_793_req_0 : boolean;
  signal type_cast_799_inst_req_0 : boolean;
  signal type_cast_799_inst_ack_0 : boolean;
  signal type_cast_799_inst_req_1 : boolean;
  signal type_cast_799_inst_ack_1 : boolean;
  signal phi_stmt_793_req_1 : boolean;
  signal phi_stmt_793_ack_0 : boolean;
  signal phi_stmt_1011_req_1 : boolean;
  signal type_cast_1014_inst_req_0 : boolean;
  signal type_cast_1014_inst_ack_0 : boolean;
  signal type_cast_1014_inst_req_1 : boolean;
  signal type_cast_1014_inst_ack_1 : boolean;
  signal phi_stmt_1011_req_0 : boolean;
  signal phi_stmt_1011_ack_0 : boolean;
  signal phi_stmt_1052_req_0 : boolean;
  signal phi_stmt_1059_req_0 : boolean;
  signal type_cast_1058_inst_req_0 : boolean;
  signal type_cast_1058_inst_ack_0 : boolean;
  signal type_cast_1058_inst_req_1 : boolean;
  signal type_cast_1058_inst_ack_1 : boolean;
  signal phi_stmt_1052_req_1 : boolean;
  signal type_cast_1065_inst_req_0 : boolean;
  signal type_cast_1065_inst_ack_0 : boolean;
  signal type_cast_1065_inst_req_1 : boolean;
  signal type_cast_1065_inst_ack_1 : boolean;
  signal phi_stmt_1059_req_1 : boolean;
  signal phi_stmt_1052_ack_0 : boolean;
  signal phi_stmt_1059_ack_0 : boolean;
  signal type_cast_1119_inst_req_0 : boolean;
  signal type_cast_1119_inst_ack_0 : boolean;
  signal type_cast_1119_inst_req_1 : boolean;
  signal type_cast_1119_inst_ack_1 : boolean;
  signal phi_stmt_1116_req_0 : boolean;
  signal phi_stmt_1116_ack_0 : boolean;
  signal phi_stmt_1289_req_0 : boolean;
  signal type_cast_1295_inst_req_0 : boolean;
  signal type_cast_1295_inst_ack_0 : boolean;
  signal type_cast_1295_inst_req_1 : boolean;
  signal type_cast_1295_inst_ack_1 : boolean;
  signal phi_stmt_1289_req_1 : boolean;
  signal phi_stmt_1289_ack_0 : boolean;
  signal type_cast_1510_inst_req_0 : boolean;
  signal type_cast_1510_inst_ack_0 : boolean;
  signal type_cast_1510_inst_req_1 : boolean;
  signal type_cast_1510_inst_ack_1 : boolean;
  signal phi_stmt_1507_req_0 : boolean;
  signal phi_stmt_1507_req_1 : boolean;
  signal phi_stmt_1507_ack_0 : boolean;
  signal phi_stmt_1552_req_0 : boolean;
  signal phi_stmt_1559_req_0 : boolean;
  signal type_cast_1558_inst_req_0 : boolean;
  signal type_cast_1558_inst_ack_0 : boolean;
  signal type_cast_1558_inst_req_1 : boolean;
  signal type_cast_1558_inst_ack_1 : boolean;
  signal phi_stmt_1552_req_1 : boolean;
  signal type_cast_1565_inst_req_0 : boolean;
  signal type_cast_1565_inst_ack_0 : boolean;
  signal type_cast_1565_inst_req_1 : boolean;
  signal type_cast_1565_inst_ack_1 : boolean;
  signal phi_stmt_1559_req_1 : boolean;
  signal phi_stmt_1552_ack_0 : boolean;
  signal phi_stmt_1559_ack_0 : boolean;
  signal type_cast_1619_inst_req_0 : boolean;
  signal type_cast_1619_inst_ack_0 : boolean;
  signal type_cast_1619_inst_req_1 : boolean;
  signal type_cast_1619_inst_ack_1 : boolean;
  signal phi_stmt_1616_req_0 : boolean;
  signal phi_stmt_1616_ack_0 : boolean;
  signal phi_stmt_1726_req_1 : boolean;
  signal type_cast_1729_inst_req_0 : boolean;
  signal type_cast_1729_inst_ack_0 : boolean;
  signal type_cast_1729_inst_req_1 : boolean;
  signal type_cast_1729_inst_ack_1 : boolean;
  signal phi_stmt_1726_req_0 : boolean;
  signal phi_stmt_1726_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convolution3D_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convolution3D_CP_1120_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convolution3D_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convolution3D_CP_1120_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convolution3D_CP_1120_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convolution3D_CP_1120_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convolution3D_CP_1120: Block -- control-path 
    signal convolution3D_CP_1120_elements: BooleanArray(430 downto 0);
    -- 
  begin -- 
    convolution3D_CP_1120_elements(0) <= convolution3D_CP_1120_start;
    convolution3D_CP_1120_symbol <= convolution3D_CP_1120_elements(362);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	6 
    -- CP-element group 0: 	13 
    -- CP-element group 0: 	20 
    -- CP-element group 0: 	27 
    -- CP-element group 0: 	34 
    -- CP-element group 0: 	41 
    -- CP-element group 0: 	48 
    -- CP-element group 0: 	55 
    -- CP-element group 0: 	62 
    -- CP-element group 0: 	69 
    -- CP-element group 0: 	76 
    -- CP-element group 0: 	83 
    -- CP-element group 0: 	90 
    -- CP-element group 0: 	97 
    -- CP-element group 0: 	104 
    -- CP-element group 0: 	111 
    -- CP-element group 0: 	114 
    -- CP-element group 0: 	117 
    -- CP-element group 0: 	120 
    -- CP-element group 0:  members (65) 
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_569_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_492_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_523_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_554_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_492_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_600_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_600_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_585_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_538_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_600_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_569_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_554_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_616_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_569_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_538_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_554_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_492_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_616_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_507_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_538_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_523_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_585_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_631_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_616_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_631_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_631_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_507_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_523_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_507_Update/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_436/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/branch_block_stmt_436__entry__
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714__entry__
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_438_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_438_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_438_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_445_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_445_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_445_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_461_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_585_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_461_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_461_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_476_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_476_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_476_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_647_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_647_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_647_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_662_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_662_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_662_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_678_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_678_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_678_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_687_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_687_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_687_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_691_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_691_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_691_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_707_update_start_
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_707_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_707_Update/cr
      -- 
    cr_1395_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1395_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_492_inst_req_1); -- 
    cr_1689_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1689_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_600_inst_req_1); -- 
    cr_1563_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1563_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_554_inst_req_1); -- 
    cr_1605_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1605_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_569_inst_req_1); -- 
    cr_1521_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1521_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_538_inst_req_1); -- 
    cr_1731_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1731_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_616_inst_req_1); -- 
    cr_1773_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1773_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_631_inst_req_1); -- 
    cr_1437_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1437_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_507_inst_req_1); -- 
    cr_1479_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1479_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_523_inst_req_1); -- 
    rr_1236_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1236_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => RPIPE_maxpool_input_pipe_438_inst_req_0); -- 
    cr_1269_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1269_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_445_inst_req_1); -- 
    cr_1647_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1647_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_585_inst_req_1); -- 
    cr_1311_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1311_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_461_inst_req_1); -- 
    cr_1353_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1353_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_476_inst_req_1); -- 
    cr_1815_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1815_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_647_inst_req_1); -- 
    cr_1857_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1857_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_662_inst_req_1); -- 
    cr_1899_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1899_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_678_inst_req_1); -- 
    cr_1913_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1913_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_687_inst_req_1); -- 
    cr_1927_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1927_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_691_inst_req_1); -- 
    cr_1941_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1941_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(0), ack => type_cast_707_inst_req_1); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_438_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_438_update_start_
      -- CP-element group 1: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_438_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_438_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_438_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_438_Update/cr
      -- 
    ra_1237_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_438_inst_ack_0, ack => convolution3D_CP_1120_elements(1)); -- 
    cr_1241_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1241_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(1), ack => RPIPE_maxpool_input_pipe_438_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	5 
    -- CP-element group 2: 	7 
    -- CP-element group 2:  members (12) 
      -- CP-element group 2: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_438_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_438_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_438_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_440_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_440_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_440_Sample/req
      -- CP-element group 2: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_445_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_445_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_445_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_454_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_454_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_454_Sample/rr
      -- 
    ca_1242_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_438_inst_ack_1, ack => convolution3D_CP_1120_elements(2)); -- 
    req_1250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(2), ack => WPIPE_maxpool_output_pipe_440_inst_req_0); -- 
    rr_1264_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1264_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(2), ack => type_cast_445_inst_req_0); -- 
    rr_1278_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1278_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(2), ack => RPIPE_maxpool_input_pipe_454_inst_req_0); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_440_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_440_update_start_
      -- CP-element group 3: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_440_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_440_Sample/ack
      -- CP-element group 3: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_440_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_440_Update/req
      -- 
    ack_1251_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_440_inst_ack_0, ack => convolution3D_CP_1120_elements(3)); -- 
    req_1255_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1255_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(3), ack => WPIPE_maxpool_output_pipe_440_inst_req_1); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	9 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_440_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_440_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_440_Update/ack
      -- 
    ack_1256_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_440_inst_ack_1, ack => convolution3D_CP_1120_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_445_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_445_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_445_Sample/ra
      -- 
    ra_1265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_445_inst_ack_0, ack => convolution3D_CP_1120_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	0 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	118 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_445_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_445_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_445_Update/ca
      -- 
    ca_1270_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_445_inst_ack_1, ack => convolution3D_CP_1120_elements(6)); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	2 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_454_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_454_update_start_
      -- CP-element group 7: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_454_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_454_Sample/ra
      -- CP-element group 7: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_454_Update/$entry
      -- CP-element group 7: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_454_Update/cr
      -- 
    ra_1279_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_454_inst_ack_0, ack => convolution3D_CP_1120_elements(7)); -- 
    cr_1283_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1283_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(7), ack => RPIPE_maxpool_input_pipe_454_inst_req_1); -- 
    -- CP-element group 8:  fork  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8: 	12 
    -- CP-element group 8: 	14 
    -- CP-element group 8:  members (9) 
      -- CP-element group 8: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_454_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_454_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_454_Update/ca
      -- CP-element group 8: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_461_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_461_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_461_Sample/rr
      -- CP-element group 8: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_469_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_469_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_469_Sample/rr
      -- 
    ca_1284_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_454_inst_ack_1, ack => convolution3D_CP_1120_elements(8)); -- 
    rr_1306_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1306_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(8), ack => type_cast_461_inst_req_0); -- 
    rr_1320_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1320_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(8), ack => RPIPE_maxpool_input_pipe_469_inst_req_0); -- 
    -- CP-element group 9:  join  transition  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	4 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_456_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_456_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_456_Sample/req
      -- 
    req_1292_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1292_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(9), ack => WPIPE_maxpool_output_pipe_456_inst_req_0); -- 
    convolution3D_cp_element_group_9: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "convolution3D_cp_element_group_9"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(4) & convolution3D_CP_1120_elements(8);
      gj_convolution3D_cp_element_group_9 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(9), clk => clk, reset => reset); --
    end block;
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_456_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_456_update_start_
      -- CP-element group 10: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_456_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_456_Sample/ack
      -- CP-element group 10: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_456_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_456_Update/req
      -- 
    ack_1293_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_456_inst_ack_0, ack => convolution3D_CP_1120_elements(10)); -- 
    req_1297_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1297_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(10), ack => WPIPE_maxpool_output_pipe_456_inst_req_1); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	16 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_456_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_456_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_456_Update/ack
      -- 
    ack_1298_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_456_inst_ack_1, ack => convolution3D_CP_1120_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	8 
    -- CP-element group 12: successors 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_461_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_461_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_461_Sample/ra
      -- 
    ra_1307_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_461_inst_ack_0, ack => convolution3D_CP_1120_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	0 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	118 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_461_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_461_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_461_Update/ca
      -- 
    ca_1312_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_461_inst_ack_1, ack => convolution3D_CP_1120_elements(13)); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	8 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_469_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_469_update_start_
      -- CP-element group 14: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_469_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_469_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_469_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_469_Update/cr
      -- 
    ra_1321_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_469_inst_ack_0, ack => convolution3D_CP_1120_elements(14)); -- 
    cr_1325_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1325_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(14), ack => RPIPE_maxpool_input_pipe_469_inst_req_1); -- 
    -- CP-element group 15:  fork  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15: 	19 
    -- CP-element group 15: 	21 
    -- CP-element group 15:  members (9) 
      -- CP-element group 15: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_469_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_469_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_469_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_476_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_476_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_476_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_485_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_485_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_485_Sample/rr
      -- 
    ca_1326_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_469_inst_ack_1, ack => convolution3D_CP_1120_elements(15)); -- 
    rr_1348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(15), ack => type_cast_476_inst_req_0); -- 
    rr_1362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(15), ack => RPIPE_maxpool_input_pipe_485_inst_req_0); -- 
    -- CP-element group 16:  join  transition  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	11 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_471_sample_start_
      -- CP-element group 16: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_471_Sample/$entry
      -- CP-element group 16: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_471_Sample/req
      -- 
    req_1334_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1334_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(16), ack => WPIPE_maxpool_output_pipe_471_inst_req_0); -- 
    convolution3D_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(11) & convolution3D_CP_1120_elements(15);
      gj_convolution3D_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_471_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_471_update_start_
      -- CP-element group 17: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_471_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_471_Sample/ack
      -- CP-element group 17: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_471_Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_471_Update/req
      -- 
    ack_1335_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_471_inst_ack_0, ack => convolution3D_CP_1120_elements(17)); -- 
    req_1339_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1339_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(17), ack => WPIPE_maxpool_output_pipe_471_inst_req_1); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	23 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_471_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_471_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_471_Update/ack
      -- 
    ack_1340_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_471_inst_ack_1, ack => convolution3D_CP_1120_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	15 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_476_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_476_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_476_Sample/ra
      -- 
    ra_1349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_476_inst_ack_0, ack => convolution3D_CP_1120_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	0 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	112 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_476_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_476_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_476_Update/ca
      -- 
    ca_1354_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_476_inst_ack_1, ack => convolution3D_CP_1120_elements(20)); -- 
    -- CP-element group 21:  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	15 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (6) 
      -- CP-element group 21: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_485_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_485_update_start_
      -- CP-element group 21: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_485_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_485_Sample/ra
      -- CP-element group 21: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_485_Update/$entry
      -- CP-element group 21: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_485_Update/cr
      -- 
    ra_1363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_485_inst_ack_0, ack => convolution3D_CP_1120_elements(21)); -- 
    cr_1367_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1367_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(21), ack => RPIPE_maxpool_input_pipe_485_inst_req_1); -- 
    -- CP-element group 22:  fork  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22: 	26 
    -- CP-element group 22: 	28 
    -- CP-element group 22:  members (9) 
      -- CP-element group 22: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_492_Sample/rr
      -- CP-element group 22: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_500_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_492_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_492_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_500_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_500_Sample/rr
      -- CP-element group 22: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_485_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_485_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_485_Update/ca
      -- 
    ca_1368_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_485_inst_ack_1, ack => convolution3D_CP_1120_elements(22)); -- 
    rr_1390_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1390_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(22), ack => type_cast_492_inst_req_0); -- 
    rr_1404_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1404_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(22), ack => RPIPE_maxpool_input_pipe_500_inst_req_0); -- 
    -- CP-element group 23:  join  transition  output  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	18 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_487_sample_start_
      -- CP-element group 23: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_487_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_487_Sample/req
      -- 
    req_1376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(23), ack => WPIPE_maxpool_output_pipe_487_inst_req_0); -- 
    convolution3D_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(18) & convolution3D_CP_1120_elements(22);
      gj_convolution3D_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  transition  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (6) 
      -- CP-element group 24: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_487_Update/req
      -- CP-element group 24: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_487_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_487_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_487_update_start_
      -- CP-element group 24: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_487_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_487_Sample/ack
      -- 
    ack_1377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_487_inst_ack_0, ack => convolution3D_CP_1120_elements(24)); -- 
    req_1381_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1381_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(24), ack => WPIPE_maxpool_output_pipe_487_inst_req_1); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	30 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_487_Update/ack
      -- CP-element group 25: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_487_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_487_update_completed_
      -- 
    ack_1382_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_487_inst_ack_1, ack => convolution3D_CP_1120_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	22 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_492_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_492_Sample/ra
      -- CP-element group 26: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_492_sample_completed_
      -- 
    ra_1391_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_492_inst_ack_0, ack => convolution3D_CP_1120_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	0 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	112 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_492_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_492_Update/ca
      -- CP-element group 27: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_492_update_completed_
      -- 
    ca_1396_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_492_inst_ack_1, ack => convolution3D_CP_1120_elements(27)); -- 
    -- CP-element group 28:  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	22 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (6) 
      -- CP-element group 28: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_500_update_start_
      -- CP-element group 28: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_500_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_500_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_500_Sample/ra
      -- CP-element group 28: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_500_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_500_Update/cr
      -- 
    ra_1405_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_500_inst_ack_0, ack => convolution3D_CP_1120_elements(28)); -- 
    cr_1409_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1409_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(28), ack => RPIPE_maxpool_input_pipe_500_inst_req_1); -- 
    -- CP-element group 29:  fork  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29: 	33 
    -- CP-element group 29: 	35 
    -- CP-element group 29:  members (9) 
      -- CP-element group 29: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_507_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_507_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_516_Sample/rr
      -- CP-element group 29: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_516_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_500_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_516_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_500_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_500_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_507_Sample/rr
      -- 
    ca_1410_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_500_inst_ack_1, ack => convolution3D_CP_1120_elements(29)); -- 
    rr_1432_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1432_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(29), ack => type_cast_507_inst_req_0); -- 
    rr_1446_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1446_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(29), ack => RPIPE_maxpool_input_pipe_516_inst_req_0); -- 
    -- CP-element group 30:  join  transition  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	25 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_502_Sample/req
      -- CP-element group 30: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_502_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_502_sample_start_
      -- 
    req_1418_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1418_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(30), ack => WPIPE_maxpool_output_pipe_502_inst_req_0); -- 
    convolution3D_cp_element_group_30: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_30"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(25) & convolution3D_CP_1120_elements(29);
      gj_convolution3D_cp_element_group_30 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(30), clk => clk, reset => reset); --
    end block;
    -- CP-element group 31:  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (6) 
      -- CP-element group 31: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_502_Update/req
      -- CP-element group 31: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_502_Update/$entry
      -- CP-element group 31: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_502_Sample/ack
      -- CP-element group 31: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_502_Sample/$exit
      -- CP-element group 31: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_502_update_start_
      -- CP-element group 31: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_502_sample_completed_
      -- 
    ack_1419_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_502_inst_ack_0, ack => convolution3D_CP_1120_elements(31)); -- 
    req_1423_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1423_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(31), ack => WPIPE_maxpool_output_pipe_502_inst_req_1); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	37 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_502_Update/ack
      -- CP-element group 32: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_502_Update/$exit
      -- CP-element group 32: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_502_update_completed_
      -- 
    ack_1424_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_502_inst_ack_1, ack => convolution3D_CP_1120_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	29 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_507_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_507_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_507_Sample/ra
      -- 
    ra_1433_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_507_inst_ack_0, ack => convolution3D_CP_1120_elements(33)); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	0 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	115 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_507_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_507_Update/ca
      -- CP-element group 34: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_507_Update/$exit
      -- 
    ca_1438_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_507_inst_ack_1, ack => convolution3D_CP_1120_elements(34)); -- 
    -- CP-element group 35:  transition  input  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	29 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (6) 
      -- CP-element group 35: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_516_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_516_Update/$entry
      -- CP-element group 35: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_516_update_start_
      -- CP-element group 35: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_516_Update/cr
      -- CP-element group 35: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_516_Sample/ra
      -- CP-element group 35: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_516_Sample/$exit
      -- 
    ra_1447_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_516_inst_ack_0, ack => convolution3D_CP_1120_elements(35)); -- 
    cr_1451_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1451_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(35), ack => RPIPE_maxpool_input_pipe_516_inst_req_1); -- 
    -- CP-element group 36:  fork  transition  input  output  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	37 
    -- CP-element group 36: 	40 
    -- CP-element group 36: 	42 
    -- CP-element group 36:  members (9) 
      -- CP-element group 36: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_531_Sample/rr
      -- CP-element group 36: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_516_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_531_Sample/$entry
      -- CP-element group 36: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_516_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_516_Update/ca
      -- CP-element group 36: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_523_Sample/$entry
      -- CP-element group 36: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_523_Sample/rr
      -- CP-element group 36: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_531_sample_start_
      -- CP-element group 36: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_523_sample_start_
      -- 
    ca_1452_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_516_inst_ack_1, ack => convolution3D_CP_1120_elements(36)); -- 
    rr_1474_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1474_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(36), ack => type_cast_523_inst_req_0); -- 
    rr_1488_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1488_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(36), ack => RPIPE_maxpool_input_pipe_531_inst_req_0); -- 
    -- CP-element group 37:  join  transition  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	32 
    -- CP-element group 37: 	36 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_518_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_518_Sample/req
      -- CP-element group 37: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_518_Sample/$entry
      -- 
    req_1460_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1460_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(37), ack => WPIPE_maxpool_output_pipe_518_inst_req_0); -- 
    convolution3D_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(32) & convolution3D_CP_1120_elements(36);
      gj_convolution3D_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (6) 
      -- CP-element group 38: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_518_Sample/ack
      -- CP-element group 38: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_518_Update/$entry
      -- CP-element group 38: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_518_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_518_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_518_update_start_
      -- CP-element group 38: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_518_Update/req
      -- 
    ack_1461_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_518_inst_ack_0, ack => convolution3D_CP_1120_elements(38)); -- 
    req_1465_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1465_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(38), ack => WPIPE_maxpool_output_pipe_518_inst_req_1); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	44 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_518_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_518_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_518_Update/ack
      -- 
    ack_1466_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_518_inst_ack_1, ack => convolution3D_CP_1120_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	36 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_523_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_523_Sample/ra
      -- CP-element group 40: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_523_sample_completed_
      -- 
    ra_1475_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_523_inst_ack_0, ack => convolution3D_CP_1120_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	0 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	115 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_523_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_523_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_523_Update/ca
      -- 
    ca_1480_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_523_inst_ack_1, ack => convolution3D_CP_1120_elements(41)); -- 
    -- CP-element group 42:  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	36 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (6) 
      -- CP-element group 42: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_531_Update/$entry
      -- CP-element group 42: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_531_Update/cr
      -- CP-element group 42: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_531_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_531_Sample/ra
      -- CP-element group 42: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_531_update_start_
      -- CP-element group 42: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_531_sample_completed_
      -- 
    ra_1489_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_531_inst_ack_0, ack => convolution3D_CP_1120_elements(42)); -- 
    cr_1493_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1493_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(42), ack => RPIPE_maxpool_input_pipe_531_inst_req_1); -- 
    -- CP-element group 43:  fork  transition  input  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43: 	47 
    -- CP-element group 43: 	49 
    -- CP-element group 43:  members (9) 
      -- CP-element group 43: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_531_Update/ca
      -- CP-element group 43: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_547_Sample/rr
      -- CP-element group 43: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_538_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_531_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_538_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_538_Sample/rr
      -- CP-element group 43: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_531_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_547_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_547_Sample/$entry
      -- 
    ca_1494_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_531_inst_ack_1, ack => convolution3D_CP_1120_elements(43)); -- 
    rr_1516_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1516_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(43), ack => type_cast_538_inst_req_0); -- 
    rr_1530_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1530_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(43), ack => RPIPE_maxpool_input_pipe_547_inst_req_0); -- 
    -- CP-element group 44:  join  transition  output  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	39 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_533_Sample/req
      -- CP-element group 44: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_533_sample_start_
      -- CP-element group 44: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_533_Sample/$entry
      -- 
    req_1502_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1502_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(44), ack => WPIPE_maxpool_output_pipe_533_inst_req_0); -- 
    convolution3D_cp_element_group_44: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_44"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(39) & convolution3D_CP_1120_elements(43);
      gj_convolution3D_cp_element_group_44 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(44), clk => clk, reset => reset); --
    end block;
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	44 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (6) 
      -- CP-element group 45: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_533_update_start_
      -- CP-element group 45: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_533_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_533_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_533_Update/$entry
      -- CP-element group 45: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_533_Sample/ack
      -- CP-element group 45: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_533_Update/req
      -- 
    ack_1503_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_533_inst_ack_0, ack => convolution3D_CP_1120_elements(45)); -- 
    req_1507_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1507_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(45), ack => WPIPE_maxpool_output_pipe_533_inst_req_1); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	51 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_533_Update/ack
      -- CP-element group 46: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_533_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_533_Update/$exit
      -- 
    ack_1508_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_533_inst_ack_1, ack => convolution3D_CP_1120_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	43 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_538_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_538_Sample/ra
      -- CP-element group 47: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_538_sample_completed_
      -- 
    ra_1517_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_538_inst_ack_0, ack => convolution3D_CP_1120_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	0 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	121 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_538_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_538_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_538_Update/ca
      -- 
    ca_1522_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_538_inst_ack_1, ack => convolution3D_CP_1120_elements(48)); -- 
    -- CP-element group 49:  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	43 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (6) 
      -- CP-element group 49: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_547_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_547_update_start_
      -- CP-element group 49: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_547_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_547_Update/cr
      -- CP-element group 49: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_547_Update/$entry
      -- CP-element group 49: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_547_Sample/ra
      -- 
    ra_1531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_547_inst_ack_0, ack => convolution3D_CP_1120_elements(49)); -- 
    cr_1535_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1535_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(49), ack => RPIPE_maxpool_input_pipe_547_inst_req_1); -- 
    -- CP-element group 50:  fork  transition  input  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50: 	54 
    -- CP-element group 50: 	56 
    -- CP-element group 50:  members (9) 
      -- CP-element group 50: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_562_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_554_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_554_Sample/rr
      -- CP-element group 50: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_562_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_562_Sample/rr
      -- CP-element group 50: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_547_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_554_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_547_Update/ca
      -- CP-element group 50: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_547_Update/$exit
      -- 
    ca_1536_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_547_inst_ack_1, ack => convolution3D_CP_1120_elements(50)); -- 
    rr_1558_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1558_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(50), ack => type_cast_554_inst_req_0); -- 
    rr_1572_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1572_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(50), ack => RPIPE_maxpool_input_pipe_562_inst_req_0); -- 
    -- CP-element group 51:  join  transition  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	46 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_549_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_549_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_549_Sample/req
      -- 
    req_1544_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1544_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(51), ack => WPIPE_maxpool_output_pipe_549_inst_req_0); -- 
    convolution3D_cp_element_group_51: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_51"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(46) & convolution3D_CP_1120_elements(50);
      gj_convolution3D_cp_element_group_51 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(51), clk => clk, reset => reset); --
    end block;
    -- CP-element group 52:  transition  input  output  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	53 
    -- CP-element group 52:  members (6) 
      -- CP-element group 52: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_549_update_start_
      -- CP-element group 52: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_549_sample_completed_
      -- CP-element group 52: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_549_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_549_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_549_Sample/ack
      -- CP-element group 52: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_549_Update/req
      -- 
    ack_1545_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_549_inst_ack_0, ack => convolution3D_CP_1120_elements(52)); -- 
    req_1549_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1549_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(52), ack => WPIPE_maxpool_output_pipe_549_inst_req_1); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	52 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	58 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_549_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_549_Update/ack
      -- CP-element group 53: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_549_Update/$exit
      -- 
    ack_1550_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_549_inst_ack_1, ack => convolution3D_CP_1120_elements(53)); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	50 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_554_Sample/ra
      -- CP-element group 54: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_554_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_554_Sample/$exit
      -- 
    ra_1559_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_554_inst_ack_0, ack => convolution3D_CP_1120_elements(54)); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	0 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	121 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_554_Update/ca
      -- CP-element group 55: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_554_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_554_update_completed_
      -- 
    ca_1564_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_554_inst_ack_1, ack => convolution3D_CP_1120_elements(55)); -- 
    -- CP-element group 56:  transition  input  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	50 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (6) 
      -- CP-element group 56: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_562_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_562_Update/cr
      -- CP-element group 56: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_562_update_start_
      -- CP-element group 56: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_562_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_562_Sample/ra
      -- CP-element group 56: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_562_Update/$entry
      -- 
    ra_1573_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_562_inst_ack_0, ack => convolution3D_CP_1120_elements(56)); -- 
    cr_1577_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1577_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(56), ack => RPIPE_maxpool_input_pipe_562_inst_req_1); -- 
    -- CP-element group 57:  fork  transition  input  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57: 	61 
    -- CP-element group 57: 	63 
    -- CP-element group 57:  members (9) 
      -- CP-element group 57: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_569_Sample/rr
      -- CP-element group 57: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_569_Sample/$entry
      -- CP-element group 57: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_578_sample_start_
      -- CP-element group 57: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_562_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_562_Update/ca
      -- CP-element group 57: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_569_sample_start_
      -- CP-element group 57: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_562_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_578_Sample/$entry
      -- CP-element group 57: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_578_Sample/rr
      -- 
    ca_1578_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_562_inst_ack_1, ack => convolution3D_CP_1120_elements(57)); -- 
    rr_1600_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1600_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(57), ack => type_cast_569_inst_req_0); -- 
    rr_1614_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1614_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(57), ack => RPIPE_maxpool_input_pipe_578_inst_req_0); -- 
    -- CP-element group 58:  join  transition  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	53 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_564_Sample/req
      -- CP-element group 58: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_564_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_564_Sample/$entry
      -- 
    req_1586_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1586_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(58), ack => WPIPE_maxpool_output_pipe_564_inst_req_0); -- 
    convolution3D_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(53) & convolution3D_CP_1120_elements(57);
      gj_convolution3D_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  transition  input  output  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59:  members (6) 
      -- CP-element group 59: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_564_Update/$entry
      -- CP-element group 59: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_564_Update/req
      -- CP-element group 59: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_564_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_564_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_564_Sample/ack
      -- CP-element group 59: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_564_update_start_
      -- 
    ack_1587_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_564_inst_ack_0, ack => convolution3D_CP_1120_elements(59)); -- 
    req_1591_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1591_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(59), ack => WPIPE_maxpool_output_pipe_564_inst_req_1); -- 
    -- CP-element group 60:  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	65 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_564_Update/ack
      -- CP-element group 60: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_564_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_564_update_completed_
      -- 
    ack_1592_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_564_inst_ack_1, ack => convolution3D_CP_1120_elements(60)); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	57 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_569_Sample/ra
      -- CP-element group 61: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_569_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_569_sample_completed_
      -- 
    ra_1601_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_569_inst_ack_0, ack => convolution3D_CP_1120_elements(61)); -- 
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	0 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	121 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_569_Update/ca
      -- CP-element group 62: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_569_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_569_update_completed_
      -- 
    ca_1606_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_569_inst_ack_1, ack => convolution3D_CP_1120_elements(62)); -- 
    -- CP-element group 63:  transition  input  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	57 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (6) 
      -- CP-element group 63: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_578_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_578_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_578_update_start_
      -- CP-element group 63: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_578_Update/cr
      -- CP-element group 63: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_578_Update/$entry
      -- CP-element group 63: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_578_Sample/ra
      -- 
    ra_1615_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_578_inst_ack_0, ack => convolution3D_CP_1120_elements(63)); -- 
    cr_1619_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1619_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(63), ack => RPIPE_maxpool_input_pipe_578_inst_req_1); -- 
    -- CP-element group 64:  fork  transition  input  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64: 	68 
    -- CP-element group 64: 	70 
    -- CP-element group 64:  members (9) 
      -- CP-element group 64: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_593_Sample/rr
      -- CP-element group 64: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_593_Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_585_Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_578_Update/ca
      -- CP-element group 64: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_585_sample_start_
      -- CP-element group 64: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_585_Sample/rr
      -- CP-element group 64: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_578_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_578_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_593_sample_start_
      -- 
    ca_1620_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_578_inst_ack_1, ack => convolution3D_CP_1120_elements(64)); -- 
    rr_1642_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1642_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(64), ack => type_cast_585_inst_req_0); -- 
    rr_1656_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1656_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(64), ack => RPIPE_maxpool_input_pipe_593_inst_req_0); -- 
    -- CP-element group 65:  join  transition  output  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	60 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_580_Sample/req
      -- CP-element group 65: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_580_sample_start_
      -- CP-element group 65: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_580_Sample/$entry
      -- 
    req_1628_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1628_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(65), ack => WPIPE_maxpool_output_pipe_580_inst_req_0); -- 
    convolution3D_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(60) & convolution3D_CP_1120_elements(64);
      gj_convolution3D_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  transition  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	65 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (6) 
      -- CP-element group 66: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_580_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_580_update_start_
      -- CP-element group 66: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_580_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_580_Sample/ack
      -- CP-element group 66: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_580_Update/req
      -- CP-element group 66: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_580_Update/$entry
      -- 
    ack_1629_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_580_inst_ack_0, ack => convolution3D_CP_1120_elements(66)); -- 
    req_1633_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1633_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(66), ack => WPIPE_maxpool_output_pipe_580_inst_req_1); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	72 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_580_Update/ack
      -- CP-element group 67: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_580_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_580_Update/$exit
      -- 
    ack_1634_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_580_inst_ack_1, ack => convolution3D_CP_1120_elements(67)); -- 
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	64 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_585_sample_completed_
      -- CP-element group 68: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_585_Sample/$exit
      -- CP-element group 68: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_585_Sample/ra
      -- 
    ra_1643_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_585_inst_ack_0, ack => convolution3D_CP_1120_elements(68)); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	0 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	121 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_585_update_completed_
      -- CP-element group 69: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_585_Update/$exit
      -- CP-element group 69: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_585_Update/ca
      -- 
    ca_1648_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_585_inst_ack_1, ack => convolution3D_CP_1120_elements(69)); -- 
    -- CP-element group 70:  transition  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	64 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70:  members (6) 
      -- CP-element group 70: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_593_Update/cr
      -- CP-element group 70: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_593_Sample/$exit
      -- CP-element group 70: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_593_Sample/ra
      -- CP-element group 70: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_593_update_start_
      -- CP-element group 70: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_593_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_593_sample_completed_
      -- 
    ra_1657_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_593_inst_ack_0, ack => convolution3D_CP_1120_elements(70)); -- 
    cr_1661_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1661_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(70), ack => RPIPE_maxpool_input_pipe_593_inst_req_1); -- 
    -- CP-element group 71:  fork  transition  input  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	72 
    -- CP-element group 71: 	75 
    -- CP-element group 71: 	77 
    -- CP-element group 71:  members (9) 
      -- CP-element group 71: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_593_Update/ca
      -- CP-element group 71: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_600_Sample/rr
      -- CP-element group 71: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_593_update_completed_
      -- CP-element group 71: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_593_Update/$exit
      -- CP-element group 71: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_609_sample_start_
      -- CP-element group 71: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_609_Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_600_Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_600_sample_start_
      -- CP-element group 71: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_609_Sample/rr
      -- 
    ca_1662_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_593_inst_ack_1, ack => convolution3D_CP_1120_elements(71)); -- 
    rr_1684_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1684_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(71), ack => type_cast_600_inst_req_0); -- 
    rr_1698_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1698_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(71), ack => RPIPE_maxpool_input_pipe_609_inst_req_0); -- 
    -- CP-element group 72:  join  transition  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	67 
    -- CP-element group 72: 	71 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	73 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_595_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_595_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_595_Sample/req
      -- 
    req_1670_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1670_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(72), ack => WPIPE_maxpool_output_pipe_595_inst_req_0); -- 
    convolution3D_cp_element_group_72: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_72"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(67) & convolution3D_CP_1120_elements(71);
      gj_convolution3D_cp_element_group_72 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(72), clk => clk, reset => reset); --
    end block;
    -- CP-element group 73:  transition  input  output  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	72 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (6) 
      -- CP-element group 73: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_595_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_595_update_start_
      -- CP-element group 73: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_595_Update/req
      -- CP-element group 73: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_595_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_595_Sample/ack
      -- CP-element group 73: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_595_Sample/$exit
      -- 
    ack_1671_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_595_inst_ack_0, ack => convolution3D_CP_1120_elements(73)); -- 
    req_1675_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1675_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(73), ack => WPIPE_maxpool_output_pipe_595_inst_req_1); -- 
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	79 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_595_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_595_Update/ack
      -- CP-element group 74: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_595_Update/$exit
      -- 
    ack_1676_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_595_inst_ack_1, ack => convolution3D_CP_1120_elements(74)); -- 
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	71 
    -- CP-element group 75: successors 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_600_Sample/$exit
      -- CP-element group 75: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_600_Sample/ra
      -- CP-element group 75: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_600_sample_completed_
      -- 
    ra_1685_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_600_inst_ack_0, ack => convolution3D_CP_1120_elements(75)); -- 
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	0 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	121 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_600_update_completed_
      -- CP-element group 76: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_600_Update/$exit
      -- CP-element group 76: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_600_Update/ca
      -- 
    ca_1690_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_600_inst_ack_1, ack => convolution3D_CP_1120_elements(76)); -- 
    -- CP-element group 77:  transition  input  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	71 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (6) 
      -- CP-element group 77: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_609_update_start_
      -- CP-element group 77: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_609_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_609_sample_completed_
      -- CP-element group 77: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_609_Update/cr
      -- CP-element group 77: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_609_Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_609_Sample/ra
      -- 
    ra_1699_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_609_inst_ack_0, ack => convolution3D_CP_1120_elements(77)); -- 
    cr_1703_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1703_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(77), ack => RPIPE_maxpool_input_pipe_609_inst_req_1); -- 
    -- CP-element group 78:  fork  transition  input  output  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78: 	82 
    -- CP-element group 78: 	84 
    -- CP-element group 78:  members (9) 
      -- CP-element group 78: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_609_update_completed_
      -- CP-element group 78: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_609_Update/ca
      -- CP-element group 78: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_624_sample_start_
      -- CP-element group 78: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_616_Sample/$entry
      -- CP-element group 78: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_609_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_616_Sample/rr
      -- CP-element group 78: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_624_Sample/$entry
      -- CP-element group 78: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_616_sample_start_
      -- CP-element group 78: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_624_Sample/rr
      -- 
    ca_1704_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_609_inst_ack_1, ack => convolution3D_CP_1120_elements(78)); -- 
    rr_1726_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1726_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(78), ack => type_cast_616_inst_req_0); -- 
    rr_1740_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1740_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(78), ack => RPIPE_maxpool_input_pipe_624_inst_req_0); -- 
    -- CP-element group 79:  join  transition  output  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	74 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_611_Sample/req
      -- CP-element group 79: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_611_sample_start_
      -- CP-element group 79: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_611_Sample/$entry
      -- 
    req_1712_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1712_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(79), ack => WPIPE_maxpool_output_pipe_611_inst_req_0); -- 
    convolution3D_cp_element_group_79: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_79"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(74) & convolution3D_CP_1120_elements(78);
      gj_convolution3D_cp_element_group_79 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(79), clk => clk, reset => reset); --
    end block;
    -- CP-element group 80:  transition  input  output  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (6) 
      -- CP-element group 80: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_611_Update/req
      -- CP-element group 80: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_611_Update/$entry
      -- CP-element group 80: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_611_sample_completed_
      -- CP-element group 80: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_611_Sample/$exit
      -- CP-element group 80: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_611_update_start_
      -- CP-element group 80: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_611_Sample/ack
      -- 
    ack_1713_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_611_inst_ack_0, ack => convolution3D_CP_1120_elements(80)); -- 
    req_1717_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1717_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(80), ack => WPIPE_maxpool_output_pipe_611_inst_req_1); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	86 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_611_Update/$exit
      -- CP-element group 81: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_611_update_completed_
      -- CP-element group 81: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_611_Update/ack
      -- 
    ack_1718_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_611_inst_ack_1, ack => convolution3D_CP_1120_elements(81)); -- 
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	78 
    -- CP-element group 82: successors 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_616_Sample/ra
      -- CP-element group 82: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_616_Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_616_sample_completed_
      -- 
    ra_1727_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_616_inst_ack_0, ack => convolution3D_CP_1120_elements(82)); -- 
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	0 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	121 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_616_update_completed_
      -- CP-element group 83: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_616_Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_616_Update/ca
      -- 
    ca_1732_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_616_inst_ack_1, ack => convolution3D_CP_1120_elements(83)); -- 
    -- CP-element group 84:  transition  input  output  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	78 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84:  members (6) 
      -- CP-element group 84: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_624_Update/$entry
      -- CP-element group 84: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_624_sample_completed_
      -- CP-element group 84: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_624_update_start_
      -- CP-element group 84: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_624_Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_624_Update/cr
      -- CP-element group 84: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_624_Sample/ra
      -- 
    ra_1741_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_624_inst_ack_0, ack => convolution3D_CP_1120_elements(84)); -- 
    cr_1745_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1745_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(84), ack => RPIPE_maxpool_input_pipe_624_inst_req_1); -- 
    -- CP-element group 85:  fork  transition  input  output  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85: 	89 
    -- CP-element group 85: 	91 
    -- CP-element group 85:  members (9) 
      -- CP-element group 85: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_624_update_completed_
      -- CP-element group 85: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_631_sample_start_
      -- CP-element group 85: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_640_Sample/$entry
      -- CP-element group 85: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_640_Sample/rr
      -- CP-element group 85: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_624_Update/ca
      -- CP-element group 85: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_631_Sample/$entry
      -- CP-element group 85: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_631_Sample/rr
      -- CP-element group 85: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_624_Update/$exit
      -- CP-element group 85: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_640_sample_start_
      -- 
    ca_1746_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_624_inst_ack_1, ack => convolution3D_CP_1120_elements(85)); -- 
    rr_1768_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1768_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(85), ack => type_cast_631_inst_req_0); -- 
    rr_1782_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1782_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(85), ack => RPIPE_maxpool_input_pipe_640_inst_req_0); -- 
    -- CP-element group 86:  join  transition  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	81 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (3) 
      -- CP-element group 86: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_626_Sample/$entry
      -- CP-element group 86: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_626_Sample/req
      -- CP-element group 86: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_626_sample_start_
      -- 
    req_1754_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1754_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(86), ack => WPIPE_maxpool_output_pipe_626_inst_req_0); -- 
    convolution3D_cp_element_group_86: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_86"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(81) & convolution3D_CP_1120_elements(85);
      gj_convolution3D_cp_element_group_86 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(86), clk => clk, reset => reset); --
    end block;
    -- CP-element group 87:  transition  input  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (6) 
      -- CP-element group 87: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_626_Update/req
      -- CP-element group 87: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_626_Sample/$exit
      -- CP-element group 87: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_626_Sample/ack
      -- CP-element group 87: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_626_sample_completed_
      -- CP-element group 87: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_626_update_start_
      -- CP-element group 87: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_626_Update/$entry
      -- 
    ack_1755_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_626_inst_ack_0, ack => convolution3D_CP_1120_elements(87)); -- 
    req_1759_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1759_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(87), ack => WPIPE_maxpool_output_pipe_626_inst_req_1); -- 
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	93 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_626_Update/ack
      -- CP-element group 88: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_626_update_completed_
      -- CP-element group 88: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_626_Update/$exit
      -- 
    ack_1760_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_626_inst_ack_1, ack => convolution3D_CP_1120_elements(88)); -- 
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	85 
    -- CP-element group 89: successors 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_631_sample_completed_
      -- CP-element group 89: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_631_Sample/$exit
      -- CP-element group 89: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_631_Sample/ra
      -- 
    ra_1769_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_631_inst_ack_0, ack => convolution3D_CP_1120_elements(89)); -- 
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	0 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	121 
    -- CP-element group 90:  members (3) 
      -- CP-element group 90: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_631_update_completed_
      -- CP-element group 90: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_631_Update/ca
      -- CP-element group 90: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_631_Update/$exit
      -- 
    ca_1774_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_631_inst_ack_1, ack => convolution3D_CP_1120_elements(90)); -- 
    -- CP-element group 91:  transition  input  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	85 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (6) 
      -- CP-element group 91: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_640_Sample/$exit
      -- CP-element group 91: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_640_Sample/ra
      -- CP-element group 91: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_640_Update/$entry
      -- CP-element group 91: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_640_Update/cr
      -- CP-element group 91: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_640_sample_completed_
      -- CP-element group 91: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_640_update_start_
      -- 
    ra_1783_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_640_inst_ack_0, ack => convolution3D_CP_1120_elements(91)); -- 
    cr_1787_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1787_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(91), ack => RPIPE_maxpool_input_pipe_640_inst_req_1); -- 
    -- CP-element group 92:  fork  transition  input  output  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	93 
    -- CP-element group 92: 	96 
    -- CP-element group 92: 	98 
    -- CP-element group 92:  members (9) 
      -- CP-element group 92: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_640_update_completed_
      -- CP-element group 92: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_640_Update/$exit
      -- CP-element group 92: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_640_Update/ca
      -- CP-element group 92: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_647_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_647_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_647_Sample/rr
      -- CP-element group 92: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_655_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_655_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_655_Sample/rr
      -- 
    ca_1788_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_640_inst_ack_1, ack => convolution3D_CP_1120_elements(92)); -- 
    rr_1810_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1810_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(92), ack => type_cast_647_inst_req_0); -- 
    rr_1824_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1824_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(92), ack => RPIPE_maxpool_input_pipe_655_inst_req_0); -- 
    -- CP-element group 93:  join  transition  output  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	88 
    -- CP-element group 93: 	92 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_642_sample_start_
      -- CP-element group 93: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_642_Sample/$entry
      -- CP-element group 93: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_642_Sample/req
      -- 
    req_1796_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1796_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(93), ack => WPIPE_maxpool_output_pipe_642_inst_req_0); -- 
    convolution3D_cp_element_group_93: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_93"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(88) & convolution3D_CP_1120_elements(92);
      gj_convolution3D_cp_element_group_93 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(93), clk => clk, reset => reset); --
    end block;
    -- CP-element group 94:  transition  input  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94:  members (6) 
      -- CP-element group 94: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_642_sample_completed_
      -- CP-element group 94: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_642_update_start_
      -- CP-element group 94: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_642_Sample/$exit
      -- CP-element group 94: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_642_Sample/ack
      -- CP-element group 94: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_642_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_642_Update/req
      -- 
    ack_1797_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_642_inst_ack_0, ack => convolution3D_CP_1120_elements(94)); -- 
    req_1801_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1801_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(94), ack => WPIPE_maxpool_output_pipe_642_inst_req_1); -- 
    -- CP-element group 95:  transition  input  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	100 
    -- CP-element group 95:  members (3) 
      -- CP-element group 95: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_642_update_completed_
      -- CP-element group 95: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_642_Update/$exit
      -- CP-element group 95: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_642_Update/ack
      -- 
    ack_1802_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_642_inst_ack_1, ack => convolution3D_CP_1120_elements(95)); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	92 
    -- CP-element group 96: successors 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_647_sample_completed_
      -- CP-element group 96: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_647_Sample/$exit
      -- CP-element group 96: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_647_Sample/ra
      -- 
    ra_1811_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_647_inst_ack_0, ack => convolution3D_CP_1120_elements(96)); -- 
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	0 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	121 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_647_update_completed_
      -- CP-element group 97: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_647_Update/$exit
      -- CP-element group 97: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_647_Update/ca
      -- 
    ca_1816_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_647_inst_ack_1, ack => convolution3D_CP_1120_elements(97)); -- 
    -- CP-element group 98:  transition  input  output  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	92 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (6) 
      -- CP-element group 98: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_655_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_655_sample_completed_
      -- CP-element group 98: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_655_update_start_
      -- CP-element group 98: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_655_Sample/$exit
      -- CP-element group 98: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_655_Sample/ra
      -- CP-element group 98: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_655_Update/cr
      -- 
    ra_1825_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_655_inst_ack_0, ack => convolution3D_CP_1120_elements(98)); -- 
    cr_1829_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1829_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(98), ack => RPIPE_maxpool_input_pipe_655_inst_req_1); -- 
    -- CP-element group 99:  fork  transition  input  output  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99: 	103 
    -- CP-element group 99: 	105 
    -- CP-element group 99:  members (9) 
      -- CP-element group 99: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_655_Update/$exit
      -- CP-element group 99: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_655_update_completed_
      -- CP-element group 99: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_655_Update/ca
      -- CP-element group 99: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_662_sample_start_
      -- CP-element group 99: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_662_Sample/$entry
      -- CP-element group 99: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_662_Sample/rr
      -- CP-element group 99: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_671_sample_start_
      -- CP-element group 99: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_671_Sample/$entry
      -- CP-element group 99: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_671_Sample/rr
      -- 
    ca_1830_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_655_inst_ack_1, ack => convolution3D_CP_1120_elements(99)); -- 
    rr_1852_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1852_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(99), ack => type_cast_662_inst_req_0); -- 
    rr_1866_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1866_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(99), ack => RPIPE_maxpool_input_pipe_671_inst_req_0); -- 
    -- CP-element group 100:  join  transition  output  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	95 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	101 
    -- CP-element group 100:  members (3) 
      -- CP-element group 100: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_657_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_657_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_657_Sample/req
      -- 
    req_1838_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1838_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(100), ack => WPIPE_maxpool_output_pipe_657_inst_req_0); -- 
    convolution3D_cp_element_group_100: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_100"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(95) & convolution3D_CP_1120_elements(99);
      gj_convolution3D_cp_element_group_100 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(100), clk => clk, reset => reset); --
    end block;
    -- CP-element group 101:  transition  input  output  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	100 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	102 
    -- CP-element group 101:  members (6) 
      -- CP-element group 101: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_657_sample_completed_
      -- CP-element group 101: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_657_update_start_
      -- CP-element group 101: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_657_Sample/$exit
      -- CP-element group 101: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_657_Sample/ack
      -- CP-element group 101: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_657_Update/$entry
      -- CP-element group 101: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_657_Update/req
      -- 
    ack_1839_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_657_inst_ack_0, ack => convolution3D_CP_1120_elements(101)); -- 
    req_1843_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1843_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(101), ack => WPIPE_maxpool_output_pipe_657_inst_req_1); -- 
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	101 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	107 
    -- CP-element group 102:  members (3) 
      -- CP-element group 102: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_657_update_completed_
      -- CP-element group 102: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_657_Update/$exit
      -- CP-element group 102: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_657_Update/ack
      -- 
    ack_1844_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_657_inst_ack_1, ack => convolution3D_CP_1120_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	99 
    -- CP-element group 103: successors 
    -- CP-element group 103:  members (3) 
      -- CP-element group 103: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_662_sample_completed_
      -- CP-element group 103: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_662_Sample/$exit
      -- CP-element group 103: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_662_Sample/ra
      -- 
    ra_1853_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_662_inst_ack_0, ack => convolution3D_CP_1120_elements(103)); -- 
    -- CP-element group 104:  transition  input  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	0 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	121 
    -- CP-element group 104:  members (3) 
      -- CP-element group 104: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_662_update_completed_
      -- CP-element group 104: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_662_Update/$exit
      -- CP-element group 104: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_662_Update/ca
      -- 
    ca_1858_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_662_inst_ack_1, ack => convolution3D_CP_1120_elements(104)); -- 
    -- CP-element group 105:  transition  input  output  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	99 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	106 
    -- CP-element group 105:  members (6) 
      -- CP-element group 105: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_671_sample_completed_
      -- CP-element group 105: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_671_update_start_
      -- CP-element group 105: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_671_Sample/$exit
      -- CP-element group 105: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_671_Sample/ra
      -- CP-element group 105: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_671_Update/$entry
      -- CP-element group 105: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_671_Update/cr
      -- 
    ra_1867_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_671_inst_ack_0, ack => convolution3D_CP_1120_elements(105)); -- 
    cr_1871_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1871_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(105), ack => RPIPE_maxpool_input_pipe_671_inst_req_1); -- 
    -- CP-element group 106:  fork  transition  input  output  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	105 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106: 	110 
    -- CP-element group 106:  members (6) 
      -- CP-element group 106: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_671_update_completed_
      -- CP-element group 106: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_671_Update/$exit
      -- CP-element group 106: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/RPIPE_maxpool_input_pipe_671_Update/ca
      -- CP-element group 106: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_678_sample_start_
      -- CP-element group 106: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_678_Sample/$entry
      -- CP-element group 106: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_678_Sample/rr
      -- 
    ca_1872_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_671_inst_ack_1, ack => convolution3D_CP_1120_elements(106)); -- 
    rr_1894_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1894_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(106), ack => type_cast_678_inst_req_0); -- 
    -- CP-element group 107:  join  transition  output  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	102 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107:  members (3) 
      -- CP-element group 107: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_673_sample_start_
      -- CP-element group 107: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_673_Sample/$entry
      -- CP-element group 107: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_673_Sample/req
      -- 
    req_1880_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1880_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(107), ack => WPIPE_maxpool_output_pipe_673_inst_req_0); -- 
    convolution3D_cp_element_group_107: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_107"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(102) & convolution3D_CP_1120_elements(106);
      gj_convolution3D_cp_element_group_107 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(107), clk => clk, reset => reset); --
    end block;
    -- CP-element group 108:  transition  input  output  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	109 
    -- CP-element group 108:  members (6) 
      -- CP-element group 108: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_673_sample_completed_
      -- CP-element group 108: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_673_update_start_
      -- CP-element group 108: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_673_Sample/$exit
      -- CP-element group 108: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_673_Sample/ack
      -- CP-element group 108: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_673_Update/$entry
      -- CP-element group 108: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_673_Update/req
      -- 
    ack_1881_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_673_inst_ack_0, ack => convolution3D_CP_1120_elements(108)); -- 
    req_1885_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1885_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(108), ack => WPIPE_maxpool_output_pipe_673_inst_req_1); -- 
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	108 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	121 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_673_update_completed_
      -- CP-element group 109: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_673_Update/$exit
      -- CP-element group 109: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/WPIPE_maxpool_output_pipe_673_Update/ack
      -- 
    ack_1886_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_673_inst_ack_1, ack => convolution3D_CP_1120_elements(109)); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	106 
    -- CP-element group 110: successors 
    -- CP-element group 110:  members (3) 
      -- CP-element group 110: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_678_sample_completed_
      -- CP-element group 110: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_678_Sample/$exit
      -- CP-element group 110: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_678_Sample/ra
      -- 
    ra_1895_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_678_inst_ack_0, ack => convolution3D_CP_1120_elements(110)); -- 
    -- CP-element group 111:  transition  input  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	0 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	121 
    -- CP-element group 111:  members (3) 
      -- CP-element group 111: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_678_update_completed_
      -- CP-element group 111: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_678_Update/$exit
      -- CP-element group 111: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_678_Update/ca
      -- 
    ca_1900_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_678_inst_ack_1, ack => convolution3D_CP_1120_elements(111)); -- 
    -- CP-element group 112:  join  transition  output  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	20 
    -- CP-element group 112: 	27 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	113 
    -- CP-element group 112:  members (3) 
      -- CP-element group 112: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_687_sample_start_
      -- CP-element group 112: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_687_Sample/$entry
      -- CP-element group 112: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_687_Sample/rr
      -- 
    rr_1908_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1908_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(112), ack => type_cast_687_inst_req_0); -- 
    convolution3D_cp_element_group_112: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_112"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(20) & convolution3D_CP_1120_elements(27);
      gj_convolution3D_cp_element_group_112 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(112), clk => clk, reset => reset); --
    end block;
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	112 
    -- CP-element group 113: successors 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_687_sample_completed_
      -- CP-element group 113: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_687_Sample/$exit
      -- CP-element group 113: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_687_Sample/ra
      -- 
    ra_1909_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_687_inst_ack_0, ack => convolution3D_CP_1120_elements(113)); -- 
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	0 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	118 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_687_update_completed_
      -- CP-element group 114: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_687_Update/$exit
      -- CP-element group 114: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_687_Update/ca
      -- 
    ca_1914_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_687_inst_ack_1, ack => convolution3D_CP_1120_elements(114)); -- 
    -- CP-element group 115:  join  transition  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	34 
    -- CP-element group 115: 	41 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	116 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_691_sample_start_
      -- CP-element group 115: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_691_Sample/$entry
      -- CP-element group 115: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_691_Sample/rr
      -- 
    rr_1922_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1922_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(115), ack => type_cast_691_inst_req_0); -- 
    convolution3D_cp_element_group_115: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_115"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(34) & convolution3D_CP_1120_elements(41);
      gj_convolution3D_cp_element_group_115 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(115), clk => clk, reset => reset); --
    end block;
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	115 
    -- CP-element group 116: successors 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_691_sample_completed_
      -- CP-element group 116: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_691_Sample/$exit
      -- CP-element group 116: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_691_Sample/ra
      -- 
    ra_1923_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_691_inst_ack_0, ack => convolution3D_CP_1120_elements(116)); -- 
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	0 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_691_update_completed_
      -- CP-element group 117: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_691_Update/$exit
      -- CP-element group 117: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_691_Update/ca
      -- 
    ca_1928_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_691_inst_ack_1, ack => convolution3D_CP_1120_elements(117)); -- 
    -- CP-element group 118:  join  transition  output  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	6 
    -- CP-element group 118: 	13 
    -- CP-element group 118: 	114 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	119 
    -- CP-element group 118:  members (3) 
      -- CP-element group 118: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_707_sample_start_
      -- CP-element group 118: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_707_Sample/$entry
      -- CP-element group 118: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_707_Sample/rr
      -- 
    rr_1936_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1936_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(118), ack => type_cast_707_inst_req_0); -- 
    convolution3D_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(6) & convolution3D_CP_1120_elements(13) & convolution3D_CP_1120_elements(114) & convolution3D_CP_1120_elements(117);
      gj_convolution3D_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  transition  input  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	118 
    -- CP-element group 119: successors 
    -- CP-element group 119:  members (3) 
      -- CP-element group 119: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_707_sample_completed_
      -- CP-element group 119: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_707_Sample/$exit
      -- CP-element group 119: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_707_Sample/ra
      -- 
    ra_1937_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_707_inst_ack_0, ack => convolution3D_CP_1120_elements(119)); -- 
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	0 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120:  members (3) 
      -- CP-element group 120: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_707_update_completed_
      -- CP-element group 120: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_707_Update/$exit
      -- CP-element group 120: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/type_cast_707_Update/ca
      -- 
    ca_1942_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_707_inst_ack_1, ack => convolution3D_CP_1120_elements(120)); -- 
    -- CP-element group 121:  branch  join  transition  place  output  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	48 
    -- CP-element group 121: 	55 
    -- CP-element group 121: 	62 
    -- CP-element group 121: 	69 
    -- CP-element group 121: 	76 
    -- CP-element group 121: 	83 
    -- CP-element group 121: 	90 
    -- CP-element group 121: 	97 
    -- CP-element group 121: 	104 
    -- CP-element group 121: 	109 
    -- CP-element group 121: 	111 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121: 	123 
    -- CP-element group 121:  members (10) 
      -- CP-element group 121: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714__exit__
      -- CP-element group 121: 	 branch_block_stmt_436/if_stmt_715__entry__
      -- CP-element group 121: 	 branch_block_stmt_436/assign_stmt_439_to_assign_stmt_714/$exit
      -- CP-element group 121: 	 branch_block_stmt_436/if_stmt_715_dead_link/$entry
      -- CP-element group 121: 	 branch_block_stmt_436/if_stmt_715_eval_test/$entry
      -- CP-element group 121: 	 branch_block_stmt_436/if_stmt_715_eval_test/$exit
      -- CP-element group 121: 	 branch_block_stmt_436/if_stmt_715_eval_test/branch_req
      -- CP-element group 121: 	 branch_block_stmt_436/R_cmp447_716_place
      -- CP-element group 121: 	 branch_block_stmt_436/if_stmt_715_if_link/$entry
      -- CP-element group 121: 	 branch_block_stmt_436/if_stmt_715_else_link/$entry
      -- 
    branch_req_1950_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1950_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(121), ack => if_stmt_715_branch_req_0); -- 
    convolution3D_cp_element_group_121: block -- 
      constant place_capacities: IntegerArray(0 to 11) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1);
      constant place_markings: IntegerArray(0 to 11)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0);
      constant place_delays: IntegerArray(0 to 11) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_121"; 
      signal preds: BooleanArray(1 to 12); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(48) & convolution3D_CP_1120_elements(55) & convolution3D_CP_1120_elements(62) & convolution3D_CP_1120_elements(69) & convolution3D_CP_1120_elements(76) & convolution3D_CP_1120_elements(83) & convolution3D_CP_1120_elements(90) & convolution3D_CP_1120_elements(97) & convolution3D_CP_1120_elements(104) & convolution3D_CP_1120_elements(109) & convolution3D_CP_1120_elements(111) & convolution3D_CP_1120_elements(120);
      gj_convolution3D_cp_element_group_121 : generic_join generic map(name => joinName, number_of_predecessors => 12, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(121), clk => clk, reset => reset); --
    end block;
    -- CP-element group 122:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	124 
    -- CP-element group 122: 	125 
    -- CP-element group 122: 	126 
    -- CP-element group 122: 	127 
    -- CP-element group 122: 	128 
    -- CP-element group 122: 	129 
    -- CP-element group 122: 	132 
    -- CP-element group 122:  members (33) 
      -- CP-element group 122: 	 branch_block_stmt_436/merge_stmt_721__exit__
      -- CP-element group 122: 	 branch_block_stmt_436/assign_stmt_726_to_assign_stmt_790__entry__
      -- CP-element group 122: 	 branch_block_stmt_436/if_stmt_715_if_link/$exit
      -- CP-element group 122: 	 branch_block_stmt_436/if_stmt_715_if_link/if_choice_transition
      -- CP-element group 122: 	 branch_block_stmt_436/entry_bbx_xnph449
      -- CP-element group 122: 	 branch_block_stmt_436/assign_stmt_726_to_assign_stmt_790/$entry
      -- CP-element group 122: 	 branch_block_stmt_436/assign_stmt_726_to_assign_stmt_790/type_cast_735_sample_start_
      -- CP-element group 122: 	 branch_block_stmt_436/assign_stmt_726_to_assign_stmt_790/type_cast_735_update_start_
      -- CP-element group 122: 	 branch_block_stmt_436/assign_stmt_726_to_assign_stmt_790/type_cast_735_Sample/$entry
      -- CP-element group 122: 	 branch_block_stmt_436/assign_stmt_726_to_assign_stmt_790/type_cast_735_Sample/rr
      -- CP-element group 122: 	 branch_block_stmt_436/assign_stmt_726_to_assign_stmt_790/type_cast_735_Update/$entry
      -- CP-element group 122: 	 branch_block_stmt_436/assign_stmt_726_to_assign_stmt_790/type_cast_735_Update/cr
      -- CP-element group 122: 	 branch_block_stmt_436/assign_stmt_726_to_assign_stmt_790/type_cast_751_sample_start_
      -- CP-element group 122: 	 branch_block_stmt_436/assign_stmt_726_to_assign_stmt_790/type_cast_751_update_start_
      -- CP-element group 122: 	 branch_block_stmt_436/assign_stmt_726_to_assign_stmt_790/type_cast_751_Sample/$entry
      -- CP-element group 122: 	 branch_block_stmt_436/assign_stmt_726_to_assign_stmt_790/type_cast_751_Sample/rr
      -- CP-element group 122: 	 branch_block_stmt_436/assign_stmt_726_to_assign_stmt_790/type_cast_751_Update/$entry
      -- CP-element group 122: 	 branch_block_stmt_436/assign_stmt_726_to_assign_stmt_790/type_cast_751_Update/cr
      -- CP-element group 122: 	 branch_block_stmt_436/assign_stmt_726_to_assign_stmt_790/type_cast_760_sample_start_
      -- CP-element group 122: 	 branch_block_stmt_436/assign_stmt_726_to_assign_stmt_790/type_cast_760_update_start_
      -- CP-element group 122: 	 branch_block_stmt_436/assign_stmt_726_to_assign_stmt_790/type_cast_760_Sample/$entry
      -- CP-element group 122: 	 branch_block_stmt_436/assign_stmt_726_to_assign_stmt_790/type_cast_760_Sample/rr
      -- CP-element group 122: 	 branch_block_stmt_436/assign_stmt_726_to_assign_stmt_790/type_cast_760_Update/$entry
      -- CP-element group 122: 	 branch_block_stmt_436/assign_stmt_726_to_assign_stmt_790/type_cast_760_Update/cr
      -- CP-element group 122: 	 branch_block_stmt_436/assign_stmt_726_to_assign_stmt_790/type_cast_770_update_start_
      -- CP-element group 122: 	 branch_block_stmt_436/assign_stmt_726_to_assign_stmt_790/type_cast_770_Update/$entry
      -- CP-element group 122: 	 branch_block_stmt_436/assign_stmt_726_to_assign_stmt_790/type_cast_770_Update/cr
      -- CP-element group 122: 	 branch_block_stmt_436/entry_bbx_xnph449_PhiReq/$entry
      -- CP-element group 122: 	 branch_block_stmt_436/entry_bbx_xnph449_PhiReq/$exit
      -- CP-element group 122: 	 branch_block_stmt_436/merge_stmt_721_PhiReqMerge
      -- CP-element group 122: 	 branch_block_stmt_436/merge_stmt_721_PhiAck/$entry
      -- CP-element group 122: 	 branch_block_stmt_436/merge_stmt_721_PhiAck/$exit
      -- CP-element group 122: 	 branch_block_stmt_436/merge_stmt_721_PhiAck/dummy
      -- 
    if_choice_transition_1955_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_715_branch_ack_1, ack => convolution3D_CP_1120_elements(122)); -- 
    rr_1972_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1972_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(122), ack => type_cast_735_inst_req_0); -- 
    cr_1977_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1977_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(122), ack => type_cast_735_inst_req_1); -- 
    rr_1986_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1986_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(122), ack => type_cast_751_inst_req_0); -- 
    cr_1991_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1991_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(122), ack => type_cast_751_inst_req_1); -- 
    rr_2000_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2000_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(122), ack => type_cast_760_inst_req_0); -- 
    cr_2005_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2005_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(122), ack => type_cast_760_inst_req_1); -- 
    cr_2019_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2019_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(122), ack => type_cast_770_inst_req_1); -- 
    -- CP-element group 123:  transition  place  input  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	121 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	369 
    -- CP-element group 123:  members (6) 
      -- CP-element group 123: 	 branch_block_stmt_436/if_stmt_715_else_link/$exit
      -- CP-element group 123: 	 branch_block_stmt_436/if_stmt_715_else_link/else_choice_transition
      -- CP-element group 123: 	 branch_block_stmt_436/entry_forx_xend
      -- CP-element group 123: 	 branch_block_stmt_436/entry_forx_xend_PhiReq/$entry
      -- CP-element group 123: 	 branch_block_stmt_436/entry_forx_xend_PhiReq/phi_stmt_1011/$entry
      -- CP-element group 123: 	 branch_block_stmt_436/entry_forx_xend_PhiReq/phi_stmt_1011/phi_stmt_1011_sources/$entry
      -- 
    else_choice_transition_1959_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_715_branch_ack_0, ack => convolution3D_CP_1120_elements(123)); -- 
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	122 
    -- CP-element group 124: successors 
    -- CP-element group 124:  members (3) 
      -- CP-element group 124: 	 branch_block_stmt_436/assign_stmt_726_to_assign_stmt_790/type_cast_735_sample_completed_
      -- CP-element group 124: 	 branch_block_stmt_436/assign_stmt_726_to_assign_stmt_790/type_cast_735_Sample/$exit
      -- CP-element group 124: 	 branch_block_stmt_436/assign_stmt_726_to_assign_stmt_790/type_cast_735_Sample/ra
      -- 
    ra_1973_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_735_inst_ack_0, ack => convolution3D_CP_1120_elements(124)); -- 
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	122 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	133 
    -- CP-element group 125:  members (3) 
      -- CP-element group 125: 	 branch_block_stmt_436/assign_stmt_726_to_assign_stmt_790/type_cast_735_update_completed_
      -- CP-element group 125: 	 branch_block_stmt_436/assign_stmt_726_to_assign_stmt_790/type_cast_735_Update/$exit
      -- CP-element group 125: 	 branch_block_stmt_436/assign_stmt_726_to_assign_stmt_790/type_cast_735_Update/ca
      -- 
    ca_1978_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_735_inst_ack_1, ack => convolution3D_CP_1120_elements(125)); -- 
    -- CP-element group 126:  transition  input  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	122 
    -- CP-element group 126: successors 
    -- CP-element group 126:  members (3) 
      -- CP-element group 126: 	 branch_block_stmt_436/assign_stmt_726_to_assign_stmt_790/type_cast_751_sample_completed_
      -- CP-element group 126: 	 branch_block_stmt_436/assign_stmt_726_to_assign_stmt_790/type_cast_751_Sample/$exit
      -- CP-element group 126: 	 branch_block_stmt_436/assign_stmt_726_to_assign_stmt_790/type_cast_751_Sample/ra
      -- 
    ra_1987_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_751_inst_ack_0, ack => convolution3D_CP_1120_elements(126)); -- 
    -- CP-element group 127:  transition  input  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	122 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	130 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 branch_block_stmt_436/assign_stmt_726_to_assign_stmt_790/type_cast_751_update_completed_
      -- CP-element group 127: 	 branch_block_stmt_436/assign_stmt_726_to_assign_stmt_790/type_cast_751_Update/$exit
      -- CP-element group 127: 	 branch_block_stmt_436/assign_stmt_726_to_assign_stmt_790/type_cast_751_Update/ca
      -- 
    ca_1992_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_751_inst_ack_1, ack => convolution3D_CP_1120_elements(127)); -- 
    -- CP-element group 128:  transition  input  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	122 
    -- CP-element group 128: successors 
    -- CP-element group 128:  members (3) 
      -- CP-element group 128: 	 branch_block_stmt_436/assign_stmt_726_to_assign_stmt_790/type_cast_760_sample_completed_
      -- CP-element group 128: 	 branch_block_stmt_436/assign_stmt_726_to_assign_stmt_790/type_cast_760_Sample/$exit
      -- CP-element group 128: 	 branch_block_stmt_436/assign_stmt_726_to_assign_stmt_790/type_cast_760_Sample/ra
      -- 
    ra_2001_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_760_inst_ack_0, ack => convolution3D_CP_1120_elements(128)); -- 
    -- CP-element group 129:  transition  input  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	122 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	130 
    -- CP-element group 129:  members (3) 
      -- CP-element group 129: 	 branch_block_stmt_436/assign_stmt_726_to_assign_stmt_790/type_cast_760_update_completed_
      -- CP-element group 129: 	 branch_block_stmt_436/assign_stmt_726_to_assign_stmt_790/type_cast_760_Update/$exit
      -- CP-element group 129: 	 branch_block_stmt_436/assign_stmt_726_to_assign_stmt_790/type_cast_760_Update/ca
      -- 
    ca_2006_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_760_inst_ack_1, ack => convolution3D_CP_1120_elements(129)); -- 
    -- CP-element group 130:  join  transition  output  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	127 
    -- CP-element group 130: 	129 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	131 
    -- CP-element group 130:  members (3) 
      -- CP-element group 130: 	 branch_block_stmt_436/assign_stmt_726_to_assign_stmt_790/type_cast_770_sample_start_
      -- CP-element group 130: 	 branch_block_stmt_436/assign_stmt_726_to_assign_stmt_790/type_cast_770_Sample/$entry
      -- CP-element group 130: 	 branch_block_stmt_436/assign_stmt_726_to_assign_stmt_790/type_cast_770_Sample/rr
      -- 
    rr_2014_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2014_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(130), ack => type_cast_770_inst_req_0); -- 
    convolution3D_cp_element_group_130: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_130"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(127) & convolution3D_CP_1120_elements(129);
      gj_convolution3D_cp_element_group_130 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(130), clk => clk, reset => reset); --
    end block;
    -- CP-element group 131:  transition  input  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	130 
    -- CP-element group 131: successors 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 branch_block_stmt_436/assign_stmt_726_to_assign_stmt_790/type_cast_770_sample_completed_
      -- CP-element group 131: 	 branch_block_stmt_436/assign_stmt_726_to_assign_stmt_790/type_cast_770_Sample/$exit
      -- CP-element group 131: 	 branch_block_stmt_436/assign_stmt_726_to_assign_stmt_790/type_cast_770_Sample/ra
      -- 
    ra_2015_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_770_inst_ack_0, ack => convolution3D_CP_1120_elements(131)); -- 
    -- CP-element group 132:  transition  input  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	122 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	133 
    -- CP-element group 132:  members (3) 
      -- CP-element group 132: 	 branch_block_stmt_436/assign_stmt_726_to_assign_stmt_790/type_cast_770_update_completed_
      -- CP-element group 132: 	 branch_block_stmt_436/assign_stmt_726_to_assign_stmt_790/type_cast_770_Update/$exit
      -- CP-element group 132: 	 branch_block_stmt_436/assign_stmt_726_to_assign_stmt_790/type_cast_770_Update/ca
      -- 
    ca_2020_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_770_inst_ack_1, ack => convolution3D_CP_1120_elements(132)); -- 
    -- CP-element group 133:  join  transition  place  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	125 
    -- CP-element group 133: 	132 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	363 
    -- CP-element group 133:  members (6) 
      -- CP-element group 133: 	 branch_block_stmt_436/assign_stmt_726_to_assign_stmt_790__exit__
      -- CP-element group 133: 	 branch_block_stmt_436/bbx_xnph449_forx_xbody
      -- CP-element group 133: 	 branch_block_stmt_436/assign_stmt_726_to_assign_stmt_790/$exit
      -- CP-element group 133: 	 branch_block_stmt_436/bbx_xnph449_forx_xbody_PhiReq/$entry
      -- CP-element group 133: 	 branch_block_stmt_436/bbx_xnph449_forx_xbody_PhiReq/phi_stmt_793/$entry
      -- CP-element group 133: 	 branch_block_stmt_436/bbx_xnph449_forx_xbody_PhiReq/phi_stmt_793/phi_stmt_793_sources/$entry
      -- 
    convolution3D_cp_element_group_133: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_133"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(125) & convolution3D_CP_1120_elements(132);
      gj_convolution3D_cp_element_group_133 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(133), clk => clk, reset => reset); --
    end block;
    -- CP-element group 134:  transition  input  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	368 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	196 
    -- CP-element group 134:  members (3) 
      -- CP-element group 134: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/array_obj_ref_805_final_index_sum_regn_sample_complete
      -- CP-element group 134: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/array_obj_ref_805_final_index_sum_regn_Sample/$exit
      -- CP-element group 134: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/array_obj_ref_805_final_index_sum_regn_Sample/ack
      -- 
    ack_2049_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_805_index_offset_ack_0, ack => convolution3D_CP_1120_elements(134)); -- 
    -- CP-element group 135:  transition  input  output  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	368 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	136 
    -- CP-element group 135:  members (11) 
      -- CP-element group 135: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/addr_of_806_sample_start_
      -- CP-element group 135: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/array_obj_ref_805_root_address_calculated
      -- CP-element group 135: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/array_obj_ref_805_offset_calculated
      -- CP-element group 135: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/array_obj_ref_805_final_index_sum_regn_Update/$exit
      -- CP-element group 135: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/array_obj_ref_805_final_index_sum_regn_Update/ack
      -- CP-element group 135: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/array_obj_ref_805_base_plus_offset/$entry
      -- CP-element group 135: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/array_obj_ref_805_base_plus_offset/$exit
      -- CP-element group 135: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/array_obj_ref_805_base_plus_offset/sum_rename_req
      -- CP-element group 135: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/array_obj_ref_805_base_plus_offset/sum_rename_ack
      -- CP-element group 135: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/addr_of_806_request/$entry
      -- CP-element group 135: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/addr_of_806_request/req
      -- 
    ack_2054_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_805_index_offset_ack_1, ack => convolution3D_CP_1120_elements(135)); -- 
    req_2063_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2063_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(135), ack => addr_of_806_final_reg_req_0); -- 
    -- CP-element group 136:  transition  input  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	135 
    -- CP-element group 136: successors 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/addr_of_806_sample_completed_
      -- CP-element group 136: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/addr_of_806_request/$exit
      -- CP-element group 136: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/addr_of_806_request/ack
      -- 
    ack_2064_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_806_final_reg_ack_0, ack => convolution3D_CP_1120_elements(136)); -- 
    -- CP-element group 137:  fork  transition  input  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	368 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	193 
    -- CP-element group 137:  members (19) 
      -- CP-element group 137: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/ptr_deref_966_word_addrgen/root_register_ack
      -- CP-element group 137: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/ptr_deref_966_word_addrgen/root_register_req
      -- CP-element group 137: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/ptr_deref_966_word_addrgen/$exit
      -- CP-element group 137: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/ptr_deref_966_word_addrgen/$entry
      -- CP-element group 137: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/ptr_deref_966_base_plus_offset/sum_rename_ack
      -- CP-element group 137: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/ptr_deref_966_base_plus_offset/sum_rename_req
      -- CP-element group 137: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/ptr_deref_966_base_plus_offset/$exit
      -- CP-element group 137: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/ptr_deref_966_base_plus_offset/$entry
      -- CP-element group 137: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/ptr_deref_966_base_addr_resize/base_resize_ack
      -- CP-element group 137: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/ptr_deref_966_base_addr_resize/base_resize_req
      -- CP-element group 137: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/ptr_deref_966_base_addr_resize/$exit
      -- CP-element group 137: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/ptr_deref_966_base_addr_resize/$entry
      -- CP-element group 137: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/ptr_deref_966_base_address_resized
      -- CP-element group 137: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/ptr_deref_966_root_address_calculated
      -- CP-element group 137: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/ptr_deref_966_word_address_calculated
      -- CP-element group 137: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/ptr_deref_966_base_address_calculated
      -- CP-element group 137: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/addr_of_806_update_completed_
      -- CP-element group 137: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/addr_of_806_complete/$exit
      -- CP-element group 137: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/addr_of_806_complete/ack
      -- 
    ack_2069_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_806_final_reg_ack_1, ack => convolution3D_CP_1120_elements(137)); -- 
    -- CP-element group 138:  transition  input  output  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	368 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	139 
    -- CP-element group 138:  members (6) 
      -- CP-element group 138: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_809_sample_completed_
      -- CP-element group 138: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_809_update_start_
      -- CP-element group 138: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_809_Sample/$exit
      -- CP-element group 138: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_809_Sample/ra
      -- CP-element group 138: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_809_Update/$entry
      -- CP-element group 138: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_809_Update/cr
      -- 
    ra_2078_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_809_inst_ack_0, ack => convolution3D_CP_1120_elements(138)); -- 
    cr_2082_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2082_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(138), ack => RPIPE_maxpool_input_pipe_809_inst_req_1); -- 
    -- CP-element group 139:  fork  transition  input  output  bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	138 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	140 
    -- CP-element group 139: 	142 
    -- CP-element group 139: 	144 
    -- CP-element group 139:  members (12) 
      -- CP-element group 139: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_809_update_completed_
      -- CP-element group 139: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_809_Update/$exit
      -- CP-element group 139: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_809_Update/ca
      -- CP-element group 139: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_811_sample_start_
      -- CP-element group 139: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_811_Sample/$entry
      -- CP-element group 139: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_811_Sample/req
      -- CP-element group 139: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_816_sample_start_
      -- CP-element group 139: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_816_Sample/$entry
      -- CP-element group 139: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_816_Sample/rr
      -- CP-element group 139: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_825_sample_start_
      -- CP-element group 139: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_825_Sample/$entry
      -- CP-element group 139: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_825_Sample/rr
      -- 
    ca_2083_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_809_inst_ack_1, ack => convolution3D_CP_1120_elements(139)); -- 
    req_2091_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2091_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(139), ack => WPIPE_maxpool_output_pipe_811_inst_req_0); -- 
    rr_2105_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2105_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(139), ack => type_cast_816_inst_req_0); -- 
    rr_2119_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2119_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(139), ack => RPIPE_maxpool_input_pipe_825_inst_req_0); -- 
    -- CP-element group 140:  transition  input  output  bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	139 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	141 
    -- CP-element group 140:  members (6) 
      -- CP-element group 140: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_811_sample_completed_
      -- CP-element group 140: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_811_update_start_
      -- CP-element group 140: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_811_Sample/$exit
      -- CP-element group 140: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_811_Sample/ack
      -- CP-element group 140: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_811_Update/$entry
      -- CP-element group 140: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_811_Update/req
      -- 
    ack_2092_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_811_inst_ack_0, ack => convolution3D_CP_1120_elements(140)); -- 
    req_2096_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2096_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(140), ack => WPIPE_maxpool_output_pipe_811_inst_req_1); -- 
    -- CP-element group 141:  transition  input  bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	140 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	146 
    -- CP-element group 141:  members (3) 
      -- CP-element group 141: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_811_update_completed_
      -- CP-element group 141: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_811_Update/$exit
      -- CP-element group 141: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_811_Update/ack
      -- 
    ack_2097_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_811_inst_ack_1, ack => convolution3D_CP_1120_elements(141)); -- 
    -- CP-element group 142:  transition  input  bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	139 
    -- CP-element group 142: successors 
    -- CP-element group 142:  members (3) 
      -- CP-element group 142: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_816_sample_completed_
      -- CP-element group 142: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_816_Sample/$exit
      -- CP-element group 142: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_816_Sample/ra
      -- 
    ra_2106_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_816_inst_ack_0, ack => convolution3D_CP_1120_elements(142)); -- 
    -- CP-element group 143:  transition  input  bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	368 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	193 
    -- CP-element group 143:  members (3) 
      -- CP-element group 143: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_816_update_completed_
      -- CP-element group 143: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_816_Update/$exit
      -- CP-element group 143: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_816_Update/ca
      -- 
    ca_2111_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_816_inst_ack_1, ack => convolution3D_CP_1120_elements(143)); -- 
    -- CP-element group 144:  transition  input  output  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	139 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	145 
    -- CP-element group 144:  members (6) 
      -- CP-element group 144: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_825_sample_completed_
      -- CP-element group 144: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_825_update_start_
      -- CP-element group 144: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_825_Sample/$exit
      -- CP-element group 144: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_825_Sample/ra
      -- CP-element group 144: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_825_Update/$entry
      -- CP-element group 144: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_825_Update/cr
      -- 
    ra_2120_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_825_inst_ack_0, ack => convolution3D_CP_1120_elements(144)); -- 
    cr_2124_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2124_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(144), ack => RPIPE_maxpool_input_pipe_825_inst_req_1); -- 
    -- CP-element group 145:  fork  transition  input  output  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	144 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	146 
    -- CP-element group 145: 	149 
    -- CP-element group 145: 	151 
    -- CP-element group 145:  members (9) 
      -- CP-element group 145: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_825_update_completed_
      -- CP-element group 145: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_825_Update/$exit
      -- CP-element group 145: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_825_Update/ca
      -- CP-element group 145: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_832_sample_start_
      -- CP-element group 145: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_832_Sample/$entry
      -- CP-element group 145: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_832_Sample/rr
      -- CP-element group 145: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_846_sample_start_
      -- CP-element group 145: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_846_Sample/$entry
      -- CP-element group 145: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_846_Sample/rr
      -- 
    ca_2125_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_825_inst_ack_1, ack => convolution3D_CP_1120_elements(145)); -- 
    rr_2147_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2147_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(145), ack => type_cast_832_inst_req_0); -- 
    rr_2161_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2161_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(145), ack => RPIPE_maxpool_input_pipe_846_inst_req_0); -- 
    -- CP-element group 146:  join  transition  output  bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	141 
    -- CP-element group 146: 	145 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	147 
    -- CP-element group 146:  members (3) 
      -- CP-element group 146: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_827_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_827_Sample/$entry
      -- CP-element group 146: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_827_Sample/req
      -- 
    req_2133_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2133_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(146), ack => WPIPE_maxpool_output_pipe_827_inst_req_0); -- 
    convolution3D_cp_element_group_146: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_146"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(141) & convolution3D_CP_1120_elements(145);
      gj_convolution3D_cp_element_group_146 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(146), clk => clk, reset => reset); --
    end block;
    -- CP-element group 147:  transition  input  output  bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	146 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	148 
    -- CP-element group 147:  members (6) 
      -- CP-element group 147: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_827_sample_completed_
      -- CP-element group 147: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_827_update_start_
      -- CP-element group 147: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_827_Sample/$exit
      -- CP-element group 147: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_827_Sample/ack
      -- CP-element group 147: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_827_Update/$entry
      -- CP-element group 147: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_827_Update/req
      -- 
    ack_2134_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_827_inst_ack_0, ack => convolution3D_CP_1120_elements(147)); -- 
    req_2138_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2138_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(147), ack => WPIPE_maxpool_output_pipe_827_inst_req_1); -- 
    -- CP-element group 148:  transition  input  bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	147 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	153 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_827_update_completed_
      -- CP-element group 148: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_827_Update/$exit
      -- CP-element group 148: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_827_Update/ack
      -- 
    ack_2139_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_827_inst_ack_1, ack => convolution3D_CP_1120_elements(148)); -- 
    -- CP-element group 149:  transition  input  bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	145 
    -- CP-element group 149: successors 
    -- CP-element group 149:  members (3) 
      -- CP-element group 149: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_832_sample_completed_
      -- CP-element group 149: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_832_Sample/$exit
      -- CP-element group 149: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_832_Sample/ra
      -- 
    ra_2148_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_832_inst_ack_0, ack => convolution3D_CP_1120_elements(149)); -- 
    -- CP-element group 150:  transition  input  bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	368 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	193 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_832_update_completed_
      -- CP-element group 150: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_832_Update/$exit
      -- CP-element group 150: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_832_Update/ca
      -- 
    ca_2153_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_832_inst_ack_1, ack => convolution3D_CP_1120_elements(150)); -- 
    -- CP-element group 151:  transition  input  output  bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	145 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	152 
    -- CP-element group 151:  members (6) 
      -- CP-element group 151: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_846_sample_completed_
      -- CP-element group 151: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_846_update_start_
      -- CP-element group 151: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_846_Sample/$exit
      -- CP-element group 151: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_846_Sample/ra
      -- CP-element group 151: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_846_Update/$entry
      -- CP-element group 151: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_846_Update/cr
      -- 
    ra_2162_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_846_inst_ack_0, ack => convolution3D_CP_1120_elements(151)); -- 
    cr_2166_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2166_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(151), ack => RPIPE_maxpool_input_pipe_846_inst_req_1); -- 
    -- CP-element group 152:  fork  transition  input  output  bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	151 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	153 
    -- CP-element group 152: 	156 
    -- CP-element group 152: 	158 
    -- CP-element group 152:  members (9) 
      -- CP-element group 152: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_846_update_completed_
      -- CP-element group 152: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_846_Update/$exit
      -- CP-element group 152: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_846_Update/ca
      -- CP-element group 152: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_853_sample_start_
      -- CP-element group 152: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_853_Sample/$entry
      -- CP-element group 152: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_853_Sample/rr
      -- CP-element group 152: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_867_sample_start_
      -- CP-element group 152: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_867_Sample/$entry
      -- CP-element group 152: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_867_Sample/rr
      -- 
    ca_2167_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_846_inst_ack_1, ack => convolution3D_CP_1120_elements(152)); -- 
    rr_2189_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2189_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(152), ack => type_cast_853_inst_req_0); -- 
    rr_2203_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2203_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(152), ack => RPIPE_maxpool_input_pipe_867_inst_req_0); -- 
    -- CP-element group 153:  join  transition  output  bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	148 
    -- CP-element group 153: 	152 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	154 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_848_sample_start_
      -- CP-element group 153: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_848_Sample/$entry
      -- CP-element group 153: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_848_Sample/req
      -- 
    req_2175_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2175_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(153), ack => WPIPE_maxpool_output_pipe_848_inst_req_0); -- 
    convolution3D_cp_element_group_153: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_153"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(148) & convolution3D_CP_1120_elements(152);
      gj_convolution3D_cp_element_group_153 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(153), clk => clk, reset => reset); --
    end block;
    -- CP-element group 154:  transition  input  output  bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	153 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	155 
    -- CP-element group 154:  members (6) 
      -- CP-element group 154: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_848_sample_completed_
      -- CP-element group 154: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_848_update_start_
      -- CP-element group 154: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_848_Sample/$exit
      -- CP-element group 154: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_848_Sample/ack
      -- CP-element group 154: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_848_Update/$entry
      -- CP-element group 154: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_848_Update/req
      -- 
    ack_2176_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_848_inst_ack_0, ack => convolution3D_CP_1120_elements(154)); -- 
    req_2180_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2180_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(154), ack => WPIPE_maxpool_output_pipe_848_inst_req_1); -- 
    -- CP-element group 155:  transition  input  bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	154 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	160 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_848_update_completed_
      -- CP-element group 155: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_848_Update/$exit
      -- CP-element group 155: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_848_Update/ack
      -- 
    ack_2181_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_848_inst_ack_1, ack => convolution3D_CP_1120_elements(155)); -- 
    -- CP-element group 156:  transition  input  bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	152 
    -- CP-element group 156: successors 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_853_sample_completed_
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_853_Sample/$exit
      -- CP-element group 156: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_853_Sample/ra
      -- 
    ra_2190_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_853_inst_ack_0, ack => convolution3D_CP_1120_elements(156)); -- 
    -- CP-element group 157:  transition  input  bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	368 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	193 
    -- CP-element group 157:  members (3) 
      -- CP-element group 157: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_853_update_completed_
      -- CP-element group 157: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_853_Update/$exit
      -- CP-element group 157: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_853_Update/ca
      -- 
    ca_2195_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_853_inst_ack_1, ack => convolution3D_CP_1120_elements(157)); -- 
    -- CP-element group 158:  transition  input  output  bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	152 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	159 
    -- CP-element group 158:  members (6) 
      -- CP-element group 158: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_867_sample_completed_
      -- CP-element group 158: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_867_update_start_
      -- CP-element group 158: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_867_Sample/$exit
      -- CP-element group 158: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_867_Sample/ra
      -- CP-element group 158: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_867_Update/$entry
      -- CP-element group 158: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_867_Update/cr
      -- 
    ra_2204_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_867_inst_ack_0, ack => convolution3D_CP_1120_elements(158)); -- 
    cr_2208_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2208_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(158), ack => RPIPE_maxpool_input_pipe_867_inst_req_1); -- 
    -- CP-element group 159:  fork  transition  input  output  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	158 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	160 
    -- CP-element group 159: 	163 
    -- CP-element group 159: 	165 
    -- CP-element group 159:  members (9) 
      -- CP-element group 159: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_867_update_completed_
      -- CP-element group 159: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_867_Update/$exit
      -- CP-element group 159: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_867_Update/ca
      -- CP-element group 159: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_874_sample_start_
      -- CP-element group 159: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_874_Sample/$entry
      -- CP-element group 159: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_874_Sample/rr
      -- CP-element group 159: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_888_sample_start_
      -- CP-element group 159: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_888_Sample/$entry
      -- CP-element group 159: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_888_Sample/rr
      -- 
    ca_2209_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_867_inst_ack_1, ack => convolution3D_CP_1120_elements(159)); -- 
    rr_2231_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2231_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(159), ack => type_cast_874_inst_req_0); -- 
    rr_2245_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2245_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(159), ack => RPIPE_maxpool_input_pipe_888_inst_req_0); -- 
    -- CP-element group 160:  join  transition  output  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	155 
    -- CP-element group 160: 	159 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	161 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_869_sample_start_
      -- CP-element group 160: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_869_Sample/$entry
      -- CP-element group 160: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_869_Sample/req
      -- 
    req_2217_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2217_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(160), ack => WPIPE_maxpool_output_pipe_869_inst_req_0); -- 
    convolution3D_cp_element_group_160: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_160"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(155) & convolution3D_CP_1120_elements(159);
      gj_convolution3D_cp_element_group_160 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(160), clk => clk, reset => reset); --
    end block;
    -- CP-element group 161:  transition  input  output  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	160 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	162 
    -- CP-element group 161:  members (6) 
      -- CP-element group 161: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_869_sample_completed_
      -- CP-element group 161: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_869_update_start_
      -- CP-element group 161: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_869_Sample/$exit
      -- CP-element group 161: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_869_Sample/ack
      -- CP-element group 161: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_869_Update/$entry
      -- CP-element group 161: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_869_Update/req
      -- 
    ack_2218_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_869_inst_ack_0, ack => convolution3D_CP_1120_elements(161)); -- 
    req_2222_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2222_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(161), ack => WPIPE_maxpool_output_pipe_869_inst_req_1); -- 
    -- CP-element group 162:  transition  input  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	161 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	167 
    -- CP-element group 162:  members (3) 
      -- CP-element group 162: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_869_update_completed_
      -- CP-element group 162: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_869_Update/$exit
      -- CP-element group 162: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_869_Update/ack
      -- 
    ack_2223_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_869_inst_ack_1, ack => convolution3D_CP_1120_elements(162)); -- 
    -- CP-element group 163:  transition  input  bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	159 
    -- CP-element group 163: successors 
    -- CP-element group 163:  members (3) 
      -- CP-element group 163: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_874_sample_completed_
      -- CP-element group 163: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_874_Sample/$exit
      -- CP-element group 163: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_874_Sample/ra
      -- 
    ra_2232_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_874_inst_ack_0, ack => convolution3D_CP_1120_elements(163)); -- 
    -- CP-element group 164:  transition  input  bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	368 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	193 
    -- CP-element group 164:  members (3) 
      -- CP-element group 164: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_874_update_completed_
      -- CP-element group 164: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_874_Update/$exit
      -- CP-element group 164: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_874_Update/ca
      -- 
    ca_2237_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_874_inst_ack_1, ack => convolution3D_CP_1120_elements(164)); -- 
    -- CP-element group 165:  transition  input  output  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	159 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	166 
    -- CP-element group 165:  members (6) 
      -- CP-element group 165: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_888_sample_completed_
      -- CP-element group 165: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_888_update_start_
      -- CP-element group 165: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_888_Sample/$exit
      -- CP-element group 165: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_888_Sample/ra
      -- CP-element group 165: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_888_Update/$entry
      -- CP-element group 165: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_888_Update/cr
      -- 
    ra_2246_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_888_inst_ack_0, ack => convolution3D_CP_1120_elements(165)); -- 
    cr_2250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(165), ack => RPIPE_maxpool_input_pipe_888_inst_req_1); -- 
    -- CP-element group 166:  fork  transition  input  output  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	165 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	167 
    -- CP-element group 166: 	170 
    -- CP-element group 166: 	172 
    -- CP-element group 166:  members (9) 
      -- CP-element group 166: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_888_update_completed_
      -- CP-element group 166: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_888_Update/$exit
      -- CP-element group 166: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_888_Update/ca
      -- CP-element group 166: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_895_sample_start_
      -- CP-element group 166: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_895_Sample/$entry
      -- CP-element group 166: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_895_Sample/rr
      -- CP-element group 166: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_909_sample_start_
      -- CP-element group 166: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_909_Sample/$entry
      -- CP-element group 166: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_909_Sample/rr
      -- 
    ca_2251_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_888_inst_ack_1, ack => convolution3D_CP_1120_elements(166)); -- 
    rr_2273_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2273_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(166), ack => type_cast_895_inst_req_0); -- 
    rr_2287_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2287_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(166), ack => RPIPE_maxpool_input_pipe_909_inst_req_0); -- 
    -- CP-element group 167:  join  transition  output  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	162 
    -- CP-element group 167: 	166 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	168 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_890_sample_start_
      -- CP-element group 167: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_890_Sample/$entry
      -- CP-element group 167: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_890_Sample/req
      -- 
    req_2259_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2259_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(167), ack => WPIPE_maxpool_output_pipe_890_inst_req_0); -- 
    convolution3D_cp_element_group_167: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_167"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(162) & convolution3D_CP_1120_elements(166);
      gj_convolution3D_cp_element_group_167 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(167), clk => clk, reset => reset); --
    end block;
    -- CP-element group 168:  transition  input  output  bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	167 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	169 
    -- CP-element group 168:  members (6) 
      -- CP-element group 168: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_890_sample_completed_
      -- CP-element group 168: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_890_update_start_
      -- CP-element group 168: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_890_Sample/$exit
      -- CP-element group 168: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_890_Sample/ack
      -- CP-element group 168: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_890_Update/$entry
      -- CP-element group 168: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_890_Update/req
      -- 
    ack_2260_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_890_inst_ack_0, ack => convolution3D_CP_1120_elements(168)); -- 
    req_2264_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2264_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(168), ack => WPIPE_maxpool_output_pipe_890_inst_req_1); -- 
    -- CP-element group 169:  transition  input  bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	168 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	174 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_890_update_completed_
      -- CP-element group 169: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_890_Update/$exit
      -- CP-element group 169: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_890_Update/ack
      -- 
    ack_2265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_890_inst_ack_1, ack => convolution3D_CP_1120_elements(169)); -- 
    -- CP-element group 170:  transition  input  bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	166 
    -- CP-element group 170: successors 
    -- CP-element group 170:  members (3) 
      -- CP-element group 170: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_895_sample_completed_
      -- CP-element group 170: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_895_Sample/$exit
      -- CP-element group 170: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_895_Sample/ra
      -- 
    ra_2274_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_895_inst_ack_0, ack => convolution3D_CP_1120_elements(170)); -- 
    -- CP-element group 171:  transition  input  bypass 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	368 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	193 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_895_update_completed_
      -- CP-element group 171: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_895_Update/$exit
      -- CP-element group 171: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_895_Update/ca
      -- 
    ca_2279_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_895_inst_ack_1, ack => convolution3D_CP_1120_elements(171)); -- 
    -- CP-element group 172:  transition  input  output  bypass 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	166 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	173 
    -- CP-element group 172:  members (6) 
      -- CP-element group 172: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_909_sample_completed_
      -- CP-element group 172: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_909_update_start_
      -- CP-element group 172: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_909_Sample/$exit
      -- CP-element group 172: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_909_Sample/ra
      -- CP-element group 172: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_909_Update/$entry
      -- CP-element group 172: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_909_Update/cr
      -- 
    ra_2288_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_909_inst_ack_0, ack => convolution3D_CP_1120_elements(172)); -- 
    cr_2292_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2292_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(172), ack => RPIPE_maxpool_input_pipe_909_inst_req_1); -- 
    -- CP-element group 173:  fork  transition  input  output  bypass 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	172 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	174 
    -- CP-element group 173: 	177 
    -- CP-element group 173: 	179 
    -- CP-element group 173:  members (9) 
      -- CP-element group 173: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_930_Sample/rr
      -- CP-element group 173: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_930_Sample/$entry
      -- CP-element group 173: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_909_update_completed_
      -- CP-element group 173: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_909_Update/$exit
      -- CP-element group 173: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_909_Update/ca
      -- CP-element group 173: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_916_sample_start_
      -- CP-element group 173: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_916_Sample/$entry
      -- CP-element group 173: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_916_Sample/rr
      -- CP-element group 173: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_930_sample_start_
      -- 
    ca_2293_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_909_inst_ack_1, ack => convolution3D_CP_1120_elements(173)); -- 
    rr_2315_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2315_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(173), ack => type_cast_916_inst_req_0); -- 
    rr_2329_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2329_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(173), ack => RPIPE_maxpool_input_pipe_930_inst_req_0); -- 
    -- CP-element group 174:  join  transition  output  bypass 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	169 
    -- CP-element group 174: 	173 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	175 
    -- CP-element group 174:  members (3) 
      -- CP-element group 174: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_911_sample_start_
      -- CP-element group 174: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_911_Sample/$entry
      -- CP-element group 174: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_911_Sample/req
      -- 
    req_2301_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2301_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(174), ack => WPIPE_maxpool_output_pipe_911_inst_req_0); -- 
    convolution3D_cp_element_group_174: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_174"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(169) & convolution3D_CP_1120_elements(173);
      gj_convolution3D_cp_element_group_174 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(174), clk => clk, reset => reset); --
    end block;
    -- CP-element group 175:  transition  input  output  bypass 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	174 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	176 
    -- CP-element group 175:  members (6) 
      -- CP-element group 175: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_911_sample_completed_
      -- CP-element group 175: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_911_update_start_
      -- CP-element group 175: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_911_Sample/$exit
      -- CP-element group 175: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_911_Sample/ack
      -- CP-element group 175: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_911_Update/$entry
      -- CP-element group 175: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_911_Update/req
      -- 
    ack_2302_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_911_inst_ack_0, ack => convolution3D_CP_1120_elements(175)); -- 
    req_2306_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2306_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(175), ack => WPIPE_maxpool_output_pipe_911_inst_req_1); -- 
    -- CP-element group 176:  transition  input  bypass 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	175 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	181 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_911_update_completed_
      -- CP-element group 176: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_911_Update/$exit
      -- CP-element group 176: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_911_Update/ack
      -- 
    ack_2307_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_911_inst_ack_1, ack => convolution3D_CP_1120_elements(176)); -- 
    -- CP-element group 177:  transition  input  bypass 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	173 
    -- CP-element group 177: successors 
    -- CP-element group 177:  members (3) 
      -- CP-element group 177: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_916_sample_completed_
      -- CP-element group 177: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_916_Sample/$exit
      -- CP-element group 177: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_916_Sample/ra
      -- 
    ra_2316_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_916_inst_ack_0, ack => convolution3D_CP_1120_elements(177)); -- 
    -- CP-element group 178:  transition  input  bypass 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	368 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	193 
    -- CP-element group 178:  members (3) 
      -- CP-element group 178: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_916_update_completed_
      -- CP-element group 178: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_916_Update/$exit
      -- CP-element group 178: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_916_Update/ca
      -- 
    ca_2321_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_916_inst_ack_1, ack => convolution3D_CP_1120_elements(178)); -- 
    -- CP-element group 179:  transition  input  output  bypass 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	173 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	180 
    -- CP-element group 179:  members (6) 
      -- CP-element group 179: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_930_Update/cr
      -- CP-element group 179: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_930_Update/$entry
      -- CP-element group 179: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_930_Sample/ra
      -- CP-element group 179: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_930_Sample/$exit
      -- CP-element group 179: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_930_sample_completed_
      -- CP-element group 179: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_930_update_start_
      -- 
    ra_2330_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_930_inst_ack_0, ack => convolution3D_CP_1120_elements(179)); -- 
    cr_2334_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2334_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(179), ack => RPIPE_maxpool_input_pipe_930_inst_req_1); -- 
    -- CP-element group 180:  fork  transition  input  output  bypass 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	179 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	181 
    -- CP-element group 180: 	184 
    -- CP-element group 180: 	186 
    -- CP-element group 180:  members (9) 
      -- CP-element group 180: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_930_Update/ca
      -- CP-element group 180: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_930_Update/$exit
      -- CP-element group 180: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_951_Sample/rr
      -- CP-element group 180: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_951_Sample/$entry
      -- CP-element group 180: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_951_sample_start_
      -- CP-element group 180: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_937_Sample/rr
      -- CP-element group 180: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_937_Sample/$entry
      -- CP-element group 180: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_930_update_completed_
      -- CP-element group 180: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_937_sample_start_
      -- 
    ca_2335_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_930_inst_ack_1, ack => convolution3D_CP_1120_elements(180)); -- 
    rr_2357_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2357_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(180), ack => type_cast_937_inst_req_0); -- 
    rr_2371_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2371_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(180), ack => RPIPE_maxpool_input_pipe_951_inst_req_0); -- 
    -- CP-element group 181:  join  transition  output  bypass 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	176 
    -- CP-element group 181: 	180 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	182 
    -- CP-element group 181:  members (3) 
      -- CP-element group 181: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_932_Sample/$entry
      -- CP-element group 181: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_932_Sample/req
      -- CP-element group 181: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_932_sample_start_
      -- 
    req_2343_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2343_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(181), ack => WPIPE_maxpool_output_pipe_932_inst_req_0); -- 
    convolution3D_cp_element_group_181: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_181"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(176) & convolution3D_CP_1120_elements(180);
      gj_convolution3D_cp_element_group_181 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(181), clk => clk, reset => reset); --
    end block;
    -- CP-element group 182:  transition  input  output  bypass 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	181 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	183 
    -- CP-element group 182:  members (6) 
      -- CP-element group 182: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_932_update_start_
      -- CP-element group 182: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_932_Sample/$exit
      -- CP-element group 182: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_932_Sample/ack
      -- CP-element group 182: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_932_Update/$entry
      -- CP-element group 182: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_932_Update/req
      -- CP-element group 182: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_932_sample_completed_
      -- 
    ack_2344_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_932_inst_ack_0, ack => convolution3D_CP_1120_elements(182)); -- 
    req_2348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(182), ack => WPIPE_maxpool_output_pipe_932_inst_req_1); -- 
    -- CP-element group 183:  transition  input  bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	182 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	188 
    -- CP-element group 183:  members (3) 
      -- CP-element group 183: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_932_update_completed_
      -- CP-element group 183: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_932_Update/$exit
      -- CP-element group 183: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_932_Update/ack
      -- 
    ack_2349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_932_inst_ack_1, ack => convolution3D_CP_1120_elements(183)); -- 
    -- CP-element group 184:  transition  input  bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	180 
    -- CP-element group 184: successors 
    -- CP-element group 184:  members (3) 
      -- CP-element group 184: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_937_Sample/ra
      -- CP-element group 184: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_937_Sample/$exit
      -- CP-element group 184: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_937_sample_completed_
      -- 
    ra_2358_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_937_inst_ack_0, ack => convolution3D_CP_1120_elements(184)); -- 
    -- CP-element group 185:  transition  input  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	368 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	193 
    -- CP-element group 185:  members (3) 
      -- CP-element group 185: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_937_Update/ca
      -- CP-element group 185: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_937_Update/$exit
      -- CP-element group 185: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_937_update_completed_
      -- 
    ca_2363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_937_inst_ack_1, ack => convolution3D_CP_1120_elements(185)); -- 
    -- CP-element group 186:  transition  input  output  bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	180 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	187 
    -- CP-element group 186:  members (6) 
      -- CP-element group 186: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_951_Update/cr
      -- CP-element group 186: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_951_Sample/ra
      -- CP-element group 186: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_951_Update/$entry
      -- CP-element group 186: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_951_Sample/$exit
      -- CP-element group 186: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_951_update_start_
      -- CP-element group 186: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_951_sample_completed_
      -- 
    ra_2372_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_951_inst_ack_0, ack => convolution3D_CP_1120_elements(186)); -- 
    cr_2376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(186), ack => RPIPE_maxpool_input_pipe_951_inst_req_1); -- 
    -- CP-element group 187:  fork  transition  input  output  bypass 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	186 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	188 
    -- CP-element group 187: 	191 
    -- CP-element group 187:  members (6) 
      -- CP-element group 187: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_951_Update/$exit
      -- CP-element group 187: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_951_Update/ca
      -- CP-element group 187: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_951_update_completed_
      -- CP-element group 187: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_958_Sample/rr
      -- CP-element group 187: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_958_Sample/$entry
      -- CP-element group 187: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_958_sample_start_
      -- 
    ca_2377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_951_inst_ack_1, ack => convolution3D_CP_1120_elements(187)); -- 
    rr_2399_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2399_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(187), ack => type_cast_958_inst_req_0); -- 
    -- CP-element group 188:  join  transition  output  bypass 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	183 
    -- CP-element group 188: 	187 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	189 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_953_Sample/$entry
      -- CP-element group 188: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_953_Sample/req
      -- CP-element group 188: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_953_sample_start_
      -- 
    req_2385_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2385_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(188), ack => WPIPE_maxpool_output_pipe_953_inst_req_0); -- 
    convolution3D_cp_element_group_188: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_188"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(183) & convolution3D_CP_1120_elements(187);
      gj_convolution3D_cp_element_group_188 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(188), clk => clk, reset => reset); --
    end block;
    -- CP-element group 189:  transition  input  output  bypass 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	188 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	190 
    -- CP-element group 189:  members (6) 
      -- CP-element group 189: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_953_Sample/$exit
      -- CP-element group 189: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_953_Sample/ack
      -- CP-element group 189: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_953_update_start_
      -- CP-element group 189: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_953_sample_completed_
      -- CP-element group 189: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_953_Update/req
      -- CP-element group 189: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_953_Update/$entry
      -- 
    ack_2386_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_953_inst_ack_0, ack => convolution3D_CP_1120_elements(189)); -- 
    req_2390_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2390_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(189), ack => WPIPE_maxpool_output_pipe_953_inst_req_1); -- 
    -- CP-element group 190:  transition  input  bypass 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	189 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	196 
    -- CP-element group 190:  members (3) 
      -- CP-element group 190: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_953_update_completed_
      -- CP-element group 190: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_953_Update/ack
      -- CP-element group 190: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/WPIPE_maxpool_output_pipe_953_Update/$exit
      -- 
    ack_2391_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_953_inst_ack_1, ack => convolution3D_CP_1120_elements(190)); -- 
    -- CP-element group 191:  transition  input  bypass 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	187 
    -- CP-element group 191: successors 
    -- CP-element group 191:  members (3) 
      -- CP-element group 191: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_958_Sample/ra
      -- CP-element group 191: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_958_Sample/$exit
      -- CP-element group 191: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_958_sample_completed_
      -- 
    ra_2400_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_958_inst_ack_0, ack => convolution3D_CP_1120_elements(191)); -- 
    -- CP-element group 192:  transition  input  bypass 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	368 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	193 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_958_Update/ca
      -- CP-element group 192: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_958_Update/$exit
      -- CP-element group 192: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_958_update_completed_
      -- 
    ca_2405_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_958_inst_ack_1, ack => convolution3D_CP_1120_elements(192)); -- 
    -- CP-element group 193:  join  transition  output  bypass 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	137 
    -- CP-element group 193: 	143 
    -- CP-element group 193: 	150 
    -- CP-element group 193: 	157 
    -- CP-element group 193: 	164 
    -- CP-element group 193: 	171 
    -- CP-element group 193: 	178 
    -- CP-element group 193: 	185 
    -- CP-element group 193: 	192 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	194 
    -- CP-element group 193:  members (9) 
      -- CP-element group 193: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/ptr_deref_966_Sample/ptr_deref_966_Split/split_req
      -- CP-element group 193: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/ptr_deref_966_Sample/ptr_deref_966_Split/$entry
      -- CP-element group 193: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/ptr_deref_966_Sample/ptr_deref_966_Split/$exit
      -- CP-element group 193: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/ptr_deref_966_Sample/$entry
      -- CP-element group 193: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/ptr_deref_966_Sample/ptr_deref_966_Split/split_ack
      -- CP-element group 193: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/ptr_deref_966_Sample/word_access_start/$entry
      -- CP-element group 193: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/ptr_deref_966_Sample/word_access_start/word_0/$entry
      -- CP-element group 193: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/ptr_deref_966_Sample/word_access_start/word_0/rr
      -- CP-element group 193: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/ptr_deref_966_sample_start_
      -- 
    rr_2443_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2443_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(193), ack => ptr_deref_966_store_0_req_0); -- 
    convolution3D_cp_element_group_193: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_193"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(137) & convolution3D_CP_1120_elements(143) & convolution3D_CP_1120_elements(150) & convolution3D_CP_1120_elements(157) & convolution3D_CP_1120_elements(164) & convolution3D_CP_1120_elements(171) & convolution3D_CP_1120_elements(178) & convolution3D_CP_1120_elements(185) & convolution3D_CP_1120_elements(192);
      gj_convolution3D_cp_element_group_193 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(193), clk => clk, reset => reset); --
    end block;
    -- CP-element group 194:  transition  input  bypass 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	193 
    -- CP-element group 194: successors 
    -- CP-element group 194:  members (5) 
      -- CP-element group 194: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/ptr_deref_966_Sample/$exit
      -- CP-element group 194: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/ptr_deref_966_Sample/word_access_start/$exit
      -- CP-element group 194: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/ptr_deref_966_Sample/word_access_start/word_0/$exit
      -- CP-element group 194: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/ptr_deref_966_Sample/word_access_start/word_0/ra
      -- CP-element group 194: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/ptr_deref_966_sample_completed_
      -- 
    ra_2444_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_966_store_0_ack_0, ack => convolution3D_CP_1120_elements(194)); -- 
    -- CP-element group 195:  transition  input  bypass 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	368 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	196 
    -- CP-element group 195:  members (5) 
      -- CP-element group 195: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/ptr_deref_966_Update/$exit
      -- CP-element group 195: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/ptr_deref_966_Update/word_access_complete/$exit
      -- CP-element group 195: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/ptr_deref_966_Update/word_access_complete/word_0/ca
      -- CP-element group 195: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/ptr_deref_966_Update/word_access_complete/word_0/$exit
      -- CP-element group 195: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/ptr_deref_966_update_completed_
      -- 
    ca_2455_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_966_store_0_ack_1, ack => convolution3D_CP_1120_elements(195)); -- 
    -- CP-element group 196:  branch  join  transition  place  output  bypass 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	134 
    -- CP-element group 196: 	190 
    -- CP-element group 196: 	195 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	197 
    -- CP-element group 196: 	198 
    -- CP-element group 196:  members (10) 
      -- CP-element group 196: 	 branch_block_stmt_436/if_stmt_980_dead_link/$entry
      -- CP-element group 196: 	 branch_block_stmt_436/if_stmt_980_eval_test/$entry
      -- CP-element group 196: 	 branch_block_stmt_436/if_stmt_980_eval_test/$exit
      -- CP-element group 196: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979__exit__
      -- CP-element group 196: 	 branch_block_stmt_436/if_stmt_980__entry__
      -- CP-element group 196: 	 branch_block_stmt_436/R_exitcond32_981_place
      -- CP-element group 196: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/$exit
      -- CP-element group 196: 	 branch_block_stmt_436/if_stmt_980_else_link/$entry
      -- CP-element group 196: 	 branch_block_stmt_436/if_stmt_980_if_link/$entry
      -- CP-element group 196: 	 branch_block_stmt_436/if_stmt_980_eval_test/branch_req
      -- 
    branch_req_2463_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2463_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(196), ack => if_stmt_980_branch_req_0); -- 
    convolution3D_cp_element_group_196: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_196"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(134) & convolution3D_CP_1120_elements(190) & convolution3D_CP_1120_elements(195);
      gj_convolution3D_cp_element_group_196 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(196), clk => clk, reset => reset); --
    end block;
    -- CP-element group 197:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	196 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	370 
    -- CP-element group 197: 	371 
    -- CP-element group 197:  members (24) 
      -- CP-element group 197: 	 branch_block_stmt_436/merge_stmt_986__exit__
      -- CP-element group 197: 	 branch_block_stmt_436/assign_stmt_993_to_assign_stmt_1008__entry__
      -- CP-element group 197: 	 branch_block_stmt_436/assign_stmt_993_to_assign_stmt_1008__exit__
      -- CP-element group 197: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend
      -- CP-element group 197: 	 branch_block_stmt_436/forx_xbody_forx_xcondx_xforx_xend_crit_edge
      -- CP-element group 197: 	 branch_block_stmt_436/assign_stmt_993_to_assign_stmt_1008/$exit
      -- CP-element group 197: 	 branch_block_stmt_436/assign_stmt_993_to_assign_stmt_1008/$entry
      -- CP-element group 197: 	 branch_block_stmt_436/if_stmt_980_if_link/if_choice_transition
      -- CP-element group 197: 	 branch_block_stmt_436/if_stmt_980_if_link/$exit
      -- CP-element group 197: 	 branch_block_stmt_436/forx_xbody_forx_xcondx_xforx_xend_crit_edge_PhiReq/$entry
      -- CP-element group 197: 	 branch_block_stmt_436/forx_xbody_forx_xcondx_xforx_xend_crit_edge_PhiReq/$exit
      -- CP-element group 197: 	 branch_block_stmt_436/merge_stmt_986_PhiReqMerge
      -- CP-element group 197: 	 branch_block_stmt_436/merge_stmt_986_PhiAck/$entry
      -- CP-element group 197: 	 branch_block_stmt_436/merge_stmt_986_PhiAck/$exit
      -- CP-element group 197: 	 branch_block_stmt_436/merge_stmt_986_PhiAck/dummy
      -- CP-element group 197: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/$entry
      -- CP-element group 197: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1011/$entry
      -- CP-element group 197: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1011/phi_stmt_1011_sources/$entry
      -- CP-element group 197: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1011/phi_stmt_1011_sources/type_cast_1014/$entry
      -- CP-element group 197: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1011/phi_stmt_1011_sources/type_cast_1014/SplitProtocol/$entry
      -- CP-element group 197: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1011/phi_stmt_1011_sources/type_cast_1014/SplitProtocol/Sample/$entry
      -- CP-element group 197: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1011/phi_stmt_1011_sources/type_cast_1014/SplitProtocol/Sample/rr
      -- CP-element group 197: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1011/phi_stmt_1011_sources/type_cast_1014/SplitProtocol/Update/$entry
      -- CP-element group 197: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1011/phi_stmt_1011_sources/type_cast_1014/SplitProtocol/Update/cr
      -- 
    if_choice_transition_2468_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_980_branch_ack_1, ack => convolution3D_CP_1120_elements(197)); -- 
    rr_3843_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3843_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(197), ack => type_cast_1014_inst_req_0); -- 
    cr_3848_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3848_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(197), ack => type_cast_1014_inst_req_1); -- 
    -- CP-element group 198:  fork  transition  place  input  output  bypass 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	196 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	364 
    -- CP-element group 198: 	365 
    -- CP-element group 198:  members (12) 
      -- CP-element group 198: 	 branch_block_stmt_436/forx_xbody_forx_xbody
      -- CP-element group 198: 	 branch_block_stmt_436/if_stmt_980_else_link/else_choice_transition
      -- CP-element group 198: 	 branch_block_stmt_436/if_stmt_980_else_link/$exit
      -- CP-element group 198: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 198: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_793/$entry
      -- CP-element group 198: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_793/phi_stmt_793_sources/$entry
      -- CP-element group 198: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_793/phi_stmt_793_sources/type_cast_799/$entry
      -- CP-element group 198: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_793/phi_stmt_793_sources/type_cast_799/SplitProtocol/$entry
      -- CP-element group 198: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_793/phi_stmt_793_sources/type_cast_799/SplitProtocol/Sample/$entry
      -- CP-element group 198: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_793/phi_stmt_793_sources/type_cast_799/SplitProtocol/Sample/rr
      -- CP-element group 198: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_793/phi_stmt_793_sources/type_cast_799/SplitProtocol/Update/$entry
      -- CP-element group 198: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_793/phi_stmt_793_sources/type_cast_799/SplitProtocol/Update/cr
      -- 
    else_choice_transition_2472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_980_branch_ack_0, ack => convolution3D_CP_1120_elements(198)); -- 
    rr_3789_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3789_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(198), ack => type_cast_799_inst_req_0); -- 
    cr_3794_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3794_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(198), ack => type_cast_799_inst_req_1); -- 
    -- CP-element group 199:  transition  place  input  bypass 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	374 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	393 
    -- CP-element group 199:  members (5) 
      -- CP-element group 199: 	 branch_block_stmt_436/forx_xend_ifx_xend
      -- CP-element group 199: 	 branch_block_stmt_436/if_stmt_1031_if_link/if_choice_transition
      -- CP-element group 199: 	 branch_block_stmt_436/if_stmt_1031_if_link/$exit
      -- CP-element group 199: 	 branch_block_stmt_436/forx_xend_ifx_xend_PhiReq/$entry
      -- CP-element group 199: 	 branch_block_stmt_436/forx_xend_ifx_xend_PhiReq/$exit
      -- 
    if_choice_transition_2493_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1031_branch_ack_1, ack => convolution3D_CP_1120_elements(199)); -- 
    -- CP-element group 200:  merge  fork  transition  place  input  bypass 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	374 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	375 
    -- CP-element group 200: 	376 
    -- CP-element group 200:  members (20) 
      -- CP-element group 200: 	 branch_block_stmt_436/forx_xend_bbx_xnphx_xi
      -- CP-element group 200: 	 branch_block_stmt_436/merge_stmt_1037__exit__
      -- CP-element group 200: 	 branch_block_stmt_436/assign_stmt_1043_to_assign_stmt_1049__entry__
      -- CP-element group 200: 	 branch_block_stmt_436/assign_stmt_1043_to_assign_stmt_1049__exit__
      -- CP-element group 200: 	 branch_block_stmt_436/bbx_xnphx_xi_forx_xbodyx_xi
      -- CP-element group 200: 	 branch_block_stmt_436/assign_stmt_1043_to_assign_stmt_1049/$exit
      -- CP-element group 200: 	 branch_block_stmt_436/assign_stmt_1043_to_assign_stmt_1049/$entry
      -- CP-element group 200: 	 branch_block_stmt_436/if_stmt_1031_else_link/else_choice_transition
      -- CP-element group 200: 	 branch_block_stmt_436/if_stmt_1031_else_link/$exit
      -- CP-element group 200: 	 branch_block_stmt_436/forx_xend_bbx_xnphx_xi_PhiReq/$entry
      -- CP-element group 200: 	 branch_block_stmt_436/forx_xend_bbx_xnphx_xi_PhiReq/$exit
      -- CP-element group 200: 	 branch_block_stmt_436/merge_stmt_1037_PhiReqMerge
      -- CP-element group 200: 	 branch_block_stmt_436/merge_stmt_1037_PhiAck/$entry
      -- CP-element group 200: 	 branch_block_stmt_436/merge_stmt_1037_PhiAck/$exit
      -- CP-element group 200: 	 branch_block_stmt_436/merge_stmt_1037_PhiAck/dummy
      -- CP-element group 200: 	 branch_block_stmt_436/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/$entry
      -- CP-element group 200: 	 branch_block_stmt_436/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1052/$entry
      -- CP-element group 200: 	 branch_block_stmt_436/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1052/phi_stmt_1052_sources/$entry
      -- CP-element group 200: 	 branch_block_stmt_436/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1059/$entry
      -- CP-element group 200: 	 branch_block_stmt_436/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1059/phi_stmt_1059_sources/$entry
      -- 
    else_choice_transition_2497_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 200_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1031_branch_ack_0, ack => convolution3D_CP_1120_elements(200)); -- 
    -- CP-element group 201:  transition  input  output  bypass 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	388 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	202 
    -- CP-element group 201:  members (6) 
      -- CP-element group 201: 	 branch_block_stmt_436/assign_stmt_1072_to_assign_stmt_1108/RPIPE_maxpool_input_pipe_1080_Update/cr
      -- CP-element group 201: 	 branch_block_stmt_436/assign_stmt_1072_to_assign_stmt_1108/RPIPE_maxpool_input_pipe_1080_Update/$entry
      -- CP-element group 201: 	 branch_block_stmt_436/assign_stmt_1072_to_assign_stmt_1108/RPIPE_maxpool_input_pipe_1080_Sample/ra
      -- CP-element group 201: 	 branch_block_stmt_436/assign_stmt_1072_to_assign_stmt_1108/RPIPE_maxpool_input_pipe_1080_Sample/$exit
      -- CP-element group 201: 	 branch_block_stmt_436/assign_stmt_1072_to_assign_stmt_1108/RPIPE_maxpool_input_pipe_1080_update_start_
      -- CP-element group 201: 	 branch_block_stmt_436/assign_stmt_1072_to_assign_stmt_1108/RPIPE_maxpool_input_pipe_1080_sample_completed_
      -- 
    ra_2514_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1080_inst_ack_0, ack => convolution3D_CP_1120_elements(201)); -- 
    cr_2518_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2518_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(201), ack => RPIPE_maxpool_input_pipe_1080_inst_req_1); -- 
    -- CP-element group 202:  fork  transition  input  output  bypass 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	201 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	203 
    -- CP-element group 202: 	205 
    -- CP-element group 202:  members (9) 
      -- CP-element group 202: 	 branch_block_stmt_436/assign_stmt_1072_to_assign_stmt_1108/WPIPE_maxpool_output_pipe_1082_Sample/$entry
      -- CP-element group 202: 	 branch_block_stmt_436/assign_stmt_1072_to_assign_stmt_1108/WPIPE_maxpool_output_pipe_1082_sample_start_
      -- CP-element group 202: 	 branch_block_stmt_436/assign_stmt_1072_to_assign_stmt_1108/RPIPE_maxpool_input_pipe_1080_Update/ca
      -- CP-element group 202: 	 branch_block_stmt_436/assign_stmt_1072_to_assign_stmt_1108/RPIPE_maxpool_input_pipe_1080_Update/$exit
      -- CP-element group 202: 	 branch_block_stmt_436/assign_stmt_1072_to_assign_stmt_1108/RPIPE_maxpool_input_pipe_1080_update_completed_
      -- CP-element group 202: 	 branch_block_stmt_436/assign_stmt_1072_to_assign_stmt_1108/type_cast_1087_Sample/rr
      -- CP-element group 202: 	 branch_block_stmt_436/assign_stmt_1072_to_assign_stmt_1108/type_cast_1087_Sample/$entry
      -- CP-element group 202: 	 branch_block_stmt_436/assign_stmt_1072_to_assign_stmt_1108/type_cast_1087_sample_start_
      -- CP-element group 202: 	 branch_block_stmt_436/assign_stmt_1072_to_assign_stmt_1108/WPIPE_maxpool_output_pipe_1082_Sample/req
      -- 
    ca_2519_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1080_inst_ack_1, ack => convolution3D_CP_1120_elements(202)); -- 
    req_2527_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2527_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(202), ack => WPIPE_maxpool_output_pipe_1082_inst_req_0); -- 
    rr_2541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(202), ack => type_cast_1087_inst_req_0); -- 
    -- CP-element group 203:  transition  input  output  bypass 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	202 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	204 
    -- CP-element group 203:  members (6) 
      -- CP-element group 203: 	 branch_block_stmt_436/assign_stmt_1072_to_assign_stmt_1108/WPIPE_maxpool_output_pipe_1082_update_start_
      -- CP-element group 203: 	 branch_block_stmt_436/assign_stmt_1072_to_assign_stmt_1108/WPIPE_maxpool_output_pipe_1082_sample_completed_
      -- CP-element group 203: 	 branch_block_stmt_436/assign_stmt_1072_to_assign_stmt_1108/WPIPE_maxpool_output_pipe_1082_Update/req
      -- CP-element group 203: 	 branch_block_stmt_436/assign_stmt_1072_to_assign_stmt_1108/WPIPE_maxpool_output_pipe_1082_Update/$entry
      -- CP-element group 203: 	 branch_block_stmt_436/assign_stmt_1072_to_assign_stmt_1108/WPIPE_maxpool_output_pipe_1082_Sample/ack
      -- CP-element group 203: 	 branch_block_stmt_436/assign_stmt_1072_to_assign_stmt_1108/WPIPE_maxpool_output_pipe_1082_Sample/$exit
      -- 
    ack_2528_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 203_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1082_inst_ack_0, ack => convolution3D_CP_1120_elements(203)); -- 
    req_2532_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2532_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(203), ack => WPIPE_maxpool_output_pipe_1082_inst_req_1); -- 
    -- CP-element group 204:  transition  input  bypass 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	203 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	209 
    -- CP-element group 204:  members (3) 
      -- CP-element group 204: 	 branch_block_stmt_436/assign_stmt_1072_to_assign_stmt_1108/WPIPE_maxpool_output_pipe_1082_update_completed_
      -- CP-element group 204: 	 branch_block_stmt_436/assign_stmt_1072_to_assign_stmt_1108/WPIPE_maxpool_output_pipe_1082_Update/ack
      -- CP-element group 204: 	 branch_block_stmt_436/assign_stmt_1072_to_assign_stmt_1108/WPIPE_maxpool_output_pipe_1082_Update/$exit
      -- 
    ack_2533_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 204_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1082_inst_ack_1, ack => convolution3D_CP_1120_elements(204)); -- 
    -- CP-element group 205:  transition  input  bypass 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	202 
    -- CP-element group 205: successors 
    -- CP-element group 205:  members (3) 
      -- CP-element group 205: 	 branch_block_stmt_436/assign_stmt_1072_to_assign_stmt_1108/type_cast_1087_Sample/ra
      -- CP-element group 205: 	 branch_block_stmt_436/assign_stmt_1072_to_assign_stmt_1108/type_cast_1087_Sample/$exit
      -- CP-element group 205: 	 branch_block_stmt_436/assign_stmt_1072_to_assign_stmt_1108/type_cast_1087_sample_completed_
      -- 
    ra_2542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1087_inst_ack_0, ack => convolution3D_CP_1120_elements(205)); -- 
    -- CP-element group 206:  transition  input  bypass 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	388 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	209 
    -- CP-element group 206:  members (3) 
      -- CP-element group 206: 	 branch_block_stmt_436/assign_stmt_1072_to_assign_stmt_1108/type_cast_1087_Update/ca
      -- CP-element group 206: 	 branch_block_stmt_436/assign_stmt_1072_to_assign_stmt_1108/type_cast_1087_Update/$exit
      -- CP-element group 206: 	 branch_block_stmt_436/assign_stmt_1072_to_assign_stmt_1108/type_cast_1087_update_completed_
      -- 
    ca_2547_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 206_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1087_inst_ack_1, ack => convolution3D_CP_1120_elements(206)); -- 
    -- CP-element group 207:  transition  input  bypass 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	388 
    -- CP-element group 207: successors 
    -- CP-element group 207:  members (3) 
      -- CP-element group 207: 	 branch_block_stmt_436/assign_stmt_1072_to_assign_stmt_1108/type_cast_1102_Sample/ra
      -- CP-element group 207: 	 branch_block_stmt_436/assign_stmt_1072_to_assign_stmt_1108/type_cast_1102_Sample/$exit
      -- CP-element group 207: 	 branch_block_stmt_436/assign_stmt_1072_to_assign_stmt_1108/type_cast_1102_sample_completed_
      -- 
    ra_2556_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 207_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1102_inst_ack_0, ack => convolution3D_CP_1120_elements(207)); -- 
    -- CP-element group 208:  transition  input  bypass 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	388 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	209 
    -- CP-element group 208:  members (3) 
      -- CP-element group 208: 	 branch_block_stmt_436/assign_stmt_1072_to_assign_stmt_1108/type_cast_1102_Update/ca
      -- CP-element group 208: 	 branch_block_stmt_436/assign_stmt_1072_to_assign_stmt_1108/type_cast_1102_Update/$exit
      -- CP-element group 208: 	 branch_block_stmt_436/assign_stmt_1072_to_assign_stmt_1108/type_cast_1102_update_completed_
      -- 
    ca_2561_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 208_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1102_inst_ack_1, ack => convolution3D_CP_1120_elements(208)); -- 
    -- CP-element group 209:  branch  join  transition  place  output  bypass 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	204 
    -- CP-element group 209: 	206 
    -- CP-element group 209: 	208 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	210 
    -- CP-element group 209: 	211 
    -- CP-element group 209:  members (10) 
      -- CP-element group 209: 	 branch_block_stmt_436/R_cmpx_xi_1110_place
      -- CP-element group 209: 	 branch_block_stmt_436/if_stmt_1109_dead_link/$entry
      -- CP-element group 209: 	 branch_block_stmt_436/if_stmt_1109_eval_test/$exit
      -- CP-element group 209: 	 branch_block_stmt_436/assign_stmt_1072_to_assign_stmt_1108__exit__
      -- CP-element group 209: 	 branch_block_stmt_436/if_stmt_1109__entry__
      -- CP-element group 209: 	 branch_block_stmt_436/if_stmt_1109_eval_test/$entry
      -- CP-element group 209: 	 branch_block_stmt_436/if_stmt_1109_else_link/$entry
      -- CP-element group 209: 	 branch_block_stmt_436/if_stmt_1109_if_link/$entry
      -- CP-element group 209: 	 branch_block_stmt_436/assign_stmt_1072_to_assign_stmt_1108/$exit
      -- CP-element group 209: 	 branch_block_stmt_436/if_stmt_1109_eval_test/branch_req
      -- 
    branch_req_2569_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2569_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(209), ack => if_stmt_1109_branch_req_0); -- 
    convolution3D_cp_element_group_209: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_209"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(204) & convolution3D_CP_1120_elements(206) & convolution3D_CP_1120_elements(208);
      gj_convolution3D_cp_element_group_209 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(209), clk => clk, reset => reset); --
    end block;
    -- CP-element group 210:  fork  transition  place  input  output  bypass 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	209 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	378 
    -- CP-element group 210: 	379 
    -- CP-element group 210: 	381 
    -- CP-element group 210: 	382 
    -- CP-element group 210:  members (20) 
      -- CP-element group 210: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi
      -- CP-element group 210: 	 branch_block_stmt_436/if_stmt_1109_if_link/if_choice_transition
      -- CP-element group 210: 	 branch_block_stmt_436/if_stmt_1109_if_link/$exit
      -- CP-element group 210: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/$entry
      -- CP-element group 210: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1052/$entry
      -- CP-element group 210: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1052/phi_stmt_1052_sources/$entry
      -- CP-element group 210: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1052/phi_stmt_1052_sources/type_cast_1058/$entry
      -- CP-element group 210: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1052/phi_stmt_1052_sources/type_cast_1058/SplitProtocol/$entry
      -- CP-element group 210: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1052/phi_stmt_1052_sources/type_cast_1058/SplitProtocol/Sample/$entry
      -- CP-element group 210: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1052/phi_stmt_1052_sources/type_cast_1058/SplitProtocol/Sample/rr
      -- CP-element group 210: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1052/phi_stmt_1052_sources/type_cast_1058/SplitProtocol/Update/$entry
      -- CP-element group 210: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1052/phi_stmt_1052_sources/type_cast_1058/SplitProtocol/Update/cr
      -- CP-element group 210: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1059/$entry
      -- CP-element group 210: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1059/phi_stmt_1059_sources/$entry
      -- CP-element group 210: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1059/phi_stmt_1059_sources/type_cast_1065/$entry
      -- CP-element group 210: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1059/phi_stmt_1059_sources/type_cast_1065/SplitProtocol/$entry
      -- CP-element group 210: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1059/phi_stmt_1059_sources/type_cast_1065/SplitProtocol/Sample/$entry
      -- CP-element group 210: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1059/phi_stmt_1059_sources/type_cast_1065/SplitProtocol/Sample/rr
      -- CP-element group 210: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1059/phi_stmt_1059_sources/type_cast_1065/SplitProtocol/Update/$entry
      -- CP-element group 210: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1059/phi_stmt_1059_sources/type_cast_1065/SplitProtocol/Update/cr
      -- 
    if_choice_transition_2574_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 210_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1109_branch_ack_1, ack => convolution3D_CP_1120_elements(210)); -- 
    rr_3905_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3905_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(210), ack => type_cast_1058_inst_req_0); -- 
    cr_3910_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3910_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(210), ack => type_cast_1058_inst_req_1); -- 
    rr_3928_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3928_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(210), ack => type_cast_1065_inst_req_0); -- 
    cr_3933_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3933_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(210), ack => type_cast_1065_inst_req_1); -- 
    -- CP-element group 211:  fork  transition  place  input  output  bypass 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	209 
    -- CP-element group 211: successors 
    -- CP-element group 211: 	389 
    -- CP-element group 211: 	390 
    -- CP-element group 211:  members (12) 
      -- CP-element group 211: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit
      -- CP-element group 211: 	 branch_block_stmt_436/if_stmt_1109_else_link/else_choice_transition
      -- CP-element group 211: 	 branch_block_stmt_436/if_stmt_1109_else_link/$exit
      -- CP-element group 211: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/$entry
      -- CP-element group 211: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1116/$entry
      -- CP-element group 211: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1116/phi_stmt_1116_sources/$entry
      -- CP-element group 211: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1116/phi_stmt_1116_sources/type_cast_1119/$entry
      -- CP-element group 211: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1116/phi_stmt_1116_sources/type_cast_1119/SplitProtocol/$entry
      -- CP-element group 211: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1116/phi_stmt_1116_sources/type_cast_1119/SplitProtocol/Sample/$entry
      -- CP-element group 211: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1116/phi_stmt_1116_sources/type_cast_1119/SplitProtocol/Sample/rr
      -- CP-element group 211: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1116/phi_stmt_1116_sources/type_cast_1119/SplitProtocol/Update/$entry
      -- CP-element group 211: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1116/phi_stmt_1116_sources/type_cast_1119/SplitProtocol/Update/cr
      -- 
    else_choice_transition_2578_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 211_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1109_branch_ack_0, ack => convolution3D_CP_1120_elements(211)); -- 
    rr_3964_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3964_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(211), ack => type_cast_1119_inst_req_0); -- 
    cr_3969_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3969_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(211), ack => type_cast_1119_inst_req_1); -- 
    -- CP-element group 212:  transition  input  bypass 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	392 
    -- CP-element group 212: successors 
    -- CP-element group 212: 	218 
    -- CP-element group 212:  members (3) 
      -- CP-element group 212: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/array_obj_ref_1148_final_index_sum_regn_Sample/$exit
      -- CP-element group 212: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/array_obj_ref_1148_final_index_sum_regn_sample_complete
      -- CP-element group 212: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/array_obj_ref_1148_final_index_sum_regn_Sample/ack
      -- 
    ack_2609_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 212_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1148_index_offset_ack_0, ack => convolution3D_CP_1120_elements(212)); -- 
    -- CP-element group 213:  transition  input  output  bypass 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	392 
    -- CP-element group 213: successors 
    -- CP-element group 213: 	214 
    -- CP-element group 213:  members (11) 
      -- CP-element group 213: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/array_obj_ref_1148_base_plus_offset/sum_rename_req
      -- CP-element group 213: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/array_obj_ref_1148_base_plus_offset/$exit
      -- CP-element group 213: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/array_obj_ref_1148_base_plus_offset/$entry
      -- CP-element group 213: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/array_obj_ref_1148_offset_calculated
      -- CP-element group 213: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/array_obj_ref_1148_root_address_calculated
      -- CP-element group 213: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/array_obj_ref_1148_final_index_sum_regn_Update/ack
      -- CP-element group 213: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/addr_of_1149_sample_start_
      -- CP-element group 213: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/array_obj_ref_1148_final_index_sum_regn_Update/$exit
      -- CP-element group 213: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/addr_of_1149_request/req
      -- CP-element group 213: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/addr_of_1149_request/$entry
      -- CP-element group 213: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/array_obj_ref_1148_base_plus_offset/sum_rename_ack
      -- 
    ack_2614_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1148_index_offset_ack_1, ack => convolution3D_CP_1120_elements(213)); -- 
    req_2623_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2623_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(213), ack => addr_of_1149_final_reg_req_0); -- 
    -- CP-element group 214:  transition  input  bypass 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	213 
    -- CP-element group 214: successors 
    -- CP-element group 214:  members (3) 
      -- CP-element group 214: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/addr_of_1149_sample_completed_
      -- CP-element group 214: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/addr_of_1149_request/ack
      -- CP-element group 214: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/addr_of_1149_request/$exit
      -- 
    ack_2624_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 214_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1149_final_reg_ack_0, ack => convolution3D_CP_1120_elements(214)); -- 
    -- CP-element group 215:  join  fork  transition  input  output  bypass 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	392 
    -- CP-element group 215: successors 
    -- CP-element group 215: 	216 
    -- CP-element group 215:  members (28) 
      -- CP-element group 215: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/ptr_deref_1152_Sample/$entry
      -- CP-element group 215: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/ptr_deref_1152_word_addrgen/root_register_ack
      -- CP-element group 215: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/ptr_deref_1152_word_addrgen/root_register_req
      -- CP-element group 215: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/ptr_deref_1152_word_addrgen/$exit
      -- CP-element group 215: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/ptr_deref_1152_word_addrgen/$entry
      -- CP-element group 215: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/addr_of_1149_update_completed_
      -- CP-element group 215: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/ptr_deref_1152_base_plus_offset/sum_rename_ack
      -- CP-element group 215: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/ptr_deref_1152_base_plus_offset/sum_rename_req
      -- CP-element group 215: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/ptr_deref_1152_base_plus_offset/$exit
      -- CP-element group 215: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/ptr_deref_1152_base_plus_offset/$entry
      -- CP-element group 215: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/ptr_deref_1152_base_addr_resize/base_resize_ack
      -- CP-element group 215: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/ptr_deref_1152_base_addr_resize/base_resize_req
      -- CP-element group 215: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/ptr_deref_1152_base_addr_resize/$exit
      -- CP-element group 215: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/ptr_deref_1152_base_addr_resize/$entry
      -- CP-element group 215: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/ptr_deref_1152_base_address_resized
      -- CP-element group 215: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/ptr_deref_1152_root_address_calculated
      -- CP-element group 215: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/ptr_deref_1152_word_address_calculated
      -- CP-element group 215: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/ptr_deref_1152_base_address_calculated
      -- CP-element group 215: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/ptr_deref_1152_Sample/word_access_start/word_0/rr
      -- CP-element group 215: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/ptr_deref_1152_Sample/word_access_start/word_0/$entry
      -- CP-element group 215: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/ptr_deref_1152_sample_start_
      -- CP-element group 215: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/addr_of_1149_complete/ack
      -- CP-element group 215: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/addr_of_1149_complete/$exit
      -- CP-element group 215: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/ptr_deref_1152_Sample/word_access_start/$entry
      -- CP-element group 215: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/ptr_deref_1152_Sample/ptr_deref_1152_Split/split_ack
      -- CP-element group 215: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/ptr_deref_1152_Sample/ptr_deref_1152_Split/split_req
      -- CP-element group 215: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/ptr_deref_1152_Sample/ptr_deref_1152_Split/$exit
      -- CP-element group 215: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/ptr_deref_1152_Sample/ptr_deref_1152_Split/$entry
      -- 
    ack_2629_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 215_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1149_final_reg_ack_1, ack => convolution3D_CP_1120_elements(215)); -- 
    rr_2667_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2667_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(215), ack => ptr_deref_1152_store_0_req_0); -- 
    -- CP-element group 216:  transition  input  bypass 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	215 
    -- CP-element group 216: successors 
    -- CP-element group 216:  members (5) 
      -- CP-element group 216: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/ptr_deref_1152_Sample/$exit
      -- CP-element group 216: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/ptr_deref_1152_Sample/word_access_start/word_0/ra
      -- CP-element group 216: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/ptr_deref_1152_Sample/word_access_start/word_0/$exit
      -- CP-element group 216: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/ptr_deref_1152_Sample/word_access_start/$exit
      -- CP-element group 216: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/ptr_deref_1152_sample_completed_
      -- 
    ra_2668_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1152_store_0_ack_0, ack => convolution3D_CP_1120_elements(216)); -- 
    -- CP-element group 217:  transition  input  bypass 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	392 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	218 
    -- CP-element group 217:  members (5) 
      -- CP-element group 217: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/ptr_deref_1152_Update/word_access_complete/word_0/ca
      -- CP-element group 217: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/ptr_deref_1152_update_completed_
      -- CP-element group 217: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/ptr_deref_1152_Update/word_access_complete/word_0/$exit
      -- CP-element group 217: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/ptr_deref_1152_Update/word_access_complete/$exit
      -- CP-element group 217: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/ptr_deref_1152_Update/$exit
      -- 
    ca_2679_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 217_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1152_store_0_ack_1, ack => convolution3D_CP_1120_elements(217)); -- 
    -- CP-element group 218:  join  transition  place  bypass 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	212 
    -- CP-element group 218: 	217 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	393 
    -- CP-element group 218:  members (5) 
      -- CP-element group 218: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154__exit__
      -- CP-element group 218: 	 branch_block_stmt_436/getRemainingElementsx_xexit_ifx_xend
      -- CP-element group 218: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/$exit
      -- CP-element group 218: 	 branch_block_stmt_436/getRemainingElementsx_xexit_ifx_xend_PhiReq/$entry
      -- CP-element group 218: 	 branch_block_stmt_436/getRemainingElementsx_xexit_ifx_xend_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_218: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_218"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(212) & convolution3D_CP_1120_elements(217);
      gj_convolution3D_cp_element_group_218 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(218), clk => clk, reset => reset); --
    end block;
    -- CP-element group 219:  transition  input  bypass 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	393 
    -- CP-element group 219: successors 
    -- CP-element group 219:  members (3) 
      -- CP-element group 219: 	 branch_block_stmt_436/assign_stmt_1160_to_assign_stmt_1208/type_cast_1159_Sample/ra
      -- CP-element group 219: 	 branch_block_stmt_436/assign_stmt_1160_to_assign_stmt_1208/type_cast_1159_Sample/$exit
      -- CP-element group 219: 	 branch_block_stmt_436/assign_stmt_1160_to_assign_stmt_1208/type_cast_1159_sample_completed_
      -- 
    ra_2691_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 219_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1159_inst_ack_0, ack => convolution3D_CP_1120_elements(219)); -- 
    -- CP-element group 220:  transition  input  bypass 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	393 
    -- CP-element group 220: successors 
    -- CP-element group 220: 	227 
    -- CP-element group 220:  members (3) 
      -- CP-element group 220: 	 branch_block_stmt_436/assign_stmt_1160_to_assign_stmt_1208/type_cast_1159_Update/$exit
      -- CP-element group 220: 	 branch_block_stmt_436/assign_stmt_1160_to_assign_stmt_1208/type_cast_1159_Update/ca
      -- CP-element group 220: 	 branch_block_stmt_436/assign_stmt_1160_to_assign_stmt_1208/type_cast_1159_update_completed_
      -- 
    ca_2696_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1159_inst_ack_1, ack => convolution3D_CP_1120_elements(220)); -- 
    -- CP-element group 221:  transition  input  bypass 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	393 
    -- CP-element group 221: successors 
    -- CP-element group 221:  members (3) 
      -- CP-element group 221: 	 branch_block_stmt_436/assign_stmt_1160_to_assign_stmt_1208/type_cast_1163_sample_completed_
      -- CP-element group 221: 	 branch_block_stmt_436/assign_stmt_1160_to_assign_stmt_1208/type_cast_1163_Sample/ra
      -- CP-element group 221: 	 branch_block_stmt_436/assign_stmt_1160_to_assign_stmt_1208/type_cast_1163_Sample/$exit
      -- 
    ra_2705_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1163_inst_ack_0, ack => convolution3D_CP_1120_elements(221)); -- 
    -- CP-element group 222:  transition  input  bypass 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	393 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	227 
    -- CP-element group 222:  members (3) 
      -- CP-element group 222: 	 branch_block_stmt_436/assign_stmt_1160_to_assign_stmt_1208/type_cast_1163_Update/ca
      -- CP-element group 222: 	 branch_block_stmt_436/assign_stmt_1160_to_assign_stmt_1208/type_cast_1163_Update/$exit
      -- CP-element group 222: 	 branch_block_stmt_436/assign_stmt_1160_to_assign_stmt_1208/type_cast_1163_update_completed_
      -- 
    ca_2710_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 222_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1163_inst_ack_1, ack => convolution3D_CP_1120_elements(222)); -- 
    -- CP-element group 223:  transition  input  bypass 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	393 
    -- CP-element group 223: successors 
    -- CP-element group 223:  members (3) 
      -- CP-element group 223: 	 branch_block_stmt_436/assign_stmt_1160_to_assign_stmt_1208/type_cast_1167_sample_completed_
      -- CP-element group 223: 	 branch_block_stmt_436/assign_stmt_1160_to_assign_stmt_1208/type_cast_1167_Sample/$exit
      -- CP-element group 223: 	 branch_block_stmt_436/assign_stmt_1160_to_assign_stmt_1208/type_cast_1167_Sample/ra
      -- 
    ra_2719_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 223_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1167_inst_ack_0, ack => convolution3D_CP_1120_elements(223)); -- 
    -- CP-element group 224:  transition  input  bypass 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	393 
    -- CP-element group 224: successors 
    -- CP-element group 224: 	227 
    -- CP-element group 224:  members (3) 
      -- CP-element group 224: 	 branch_block_stmt_436/assign_stmt_1160_to_assign_stmt_1208/type_cast_1167_update_completed_
      -- CP-element group 224: 	 branch_block_stmt_436/assign_stmt_1160_to_assign_stmt_1208/type_cast_1167_Update/ca
      -- CP-element group 224: 	 branch_block_stmt_436/assign_stmt_1160_to_assign_stmt_1208/type_cast_1167_Update/$exit
      -- 
    ca_2724_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1167_inst_ack_1, ack => convolution3D_CP_1120_elements(224)); -- 
    -- CP-element group 225:  transition  input  bypass 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	393 
    -- CP-element group 225: successors 
    -- CP-element group 225:  members (3) 
      -- CP-element group 225: 	 branch_block_stmt_436/assign_stmt_1160_to_assign_stmt_1208/type_cast_1171_Sample/$exit
      -- CP-element group 225: 	 branch_block_stmt_436/assign_stmt_1160_to_assign_stmt_1208/type_cast_1171_sample_completed_
      -- CP-element group 225: 	 branch_block_stmt_436/assign_stmt_1160_to_assign_stmt_1208/type_cast_1171_Sample/ra
      -- 
    ra_2733_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 225_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1171_inst_ack_0, ack => convolution3D_CP_1120_elements(225)); -- 
    -- CP-element group 226:  transition  input  bypass 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	393 
    -- CP-element group 226: successors 
    -- CP-element group 226: 	227 
    -- CP-element group 226:  members (3) 
      -- CP-element group 226: 	 branch_block_stmt_436/assign_stmt_1160_to_assign_stmt_1208/type_cast_1171_update_completed_
      -- CP-element group 226: 	 branch_block_stmt_436/assign_stmt_1160_to_assign_stmt_1208/type_cast_1171_Update/$exit
      -- CP-element group 226: 	 branch_block_stmt_436/assign_stmt_1160_to_assign_stmt_1208/type_cast_1171_Update/ca
      -- 
    ca_2738_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 226_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1171_inst_ack_1, ack => convolution3D_CP_1120_elements(226)); -- 
    -- CP-element group 227:  branch  join  transition  place  output  bypass 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	220 
    -- CP-element group 227: 	222 
    -- CP-element group 227: 	224 
    -- CP-element group 227: 	226 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	228 
    -- CP-element group 227: 	229 
    -- CP-element group 227:  members (10) 
      -- CP-element group 227: 	 branch_block_stmt_436/assign_stmt_1160_to_assign_stmt_1208__exit__
      -- CP-element group 227: 	 branch_block_stmt_436/if_stmt_1209__entry__
      -- CP-element group 227: 	 branch_block_stmt_436/assign_stmt_1160_to_assign_stmt_1208/$exit
      -- CP-element group 227: 	 branch_block_stmt_436/if_stmt_1209_dead_link/$entry
      -- CP-element group 227: 	 branch_block_stmt_436/if_stmt_1209_eval_test/$entry
      -- CP-element group 227: 	 branch_block_stmt_436/if_stmt_1209_eval_test/$exit
      -- CP-element group 227: 	 branch_block_stmt_436/if_stmt_1209_eval_test/branch_req
      -- CP-element group 227: 	 branch_block_stmt_436/R_cmp255443_1210_place
      -- CP-element group 227: 	 branch_block_stmt_436/if_stmt_1209_if_link/$entry
      -- CP-element group 227: 	 branch_block_stmt_436/if_stmt_1209_else_link/$entry
      -- 
    branch_req_2746_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2746_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(227), ack => if_stmt_1209_branch_req_0); -- 
    convolution3D_cp_element_group_227: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_227"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(220) & convolution3D_CP_1120_elements(222) & convolution3D_CP_1120_elements(224) & convolution3D_CP_1120_elements(226);
      gj_convolution3D_cp_element_group_227 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(227), clk => clk, reset => reset); --
    end block;
    -- CP-element group 228:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	227 
    -- CP-element group 228: successors 
    -- CP-element group 228: 	230 
    -- CP-element group 228: 	231 
    -- CP-element group 228: 	232 
    -- CP-element group 228: 	233 
    -- CP-element group 228: 	234 
    -- CP-element group 228: 	235 
    -- CP-element group 228: 	236 
    -- CP-element group 228: 	237 
    -- CP-element group 228: 	240 
    -- CP-element group 228: 	242 
    -- CP-element group 228:  members (42) 
      -- CP-element group 228: 	 branch_block_stmt_436/merge_stmt_1215__exit__
      -- CP-element group 228: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286__entry__
      -- CP-element group 228: 	 branch_block_stmt_436/if_stmt_1209_if_link/$exit
      -- CP-element group 228: 	 branch_block_stmt_436/if_stmt_1209_if_link/if_choice_transition
      -- CP-element group 228: 	 branch_block_stmt_436/ifx_xend_bbx_xnph
      -- CP-element group 228: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/$entry
      -- CP-element group 228: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1230_sample_start_
      -- CP-element group 228: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1230_update_start_
      -- CP-element group 228: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1230_Sample/$entry
      -- CP-element group 228: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1230_Sample/rr
      -- CP-element group 228: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1230_Update/$entry
      -- CP-element group 228: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1230_Update/cr
      -- CP-element group 228: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1234_sample_start_
      -- CP-element group 228: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1234_update_start_
      -- CP-element group 228: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1234_Sample/$entry
      -- CP-element group 228: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1234_Sample/rr
      -- CP-element group 228: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1234_Update/$entry
      -- CP-element group 228: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1234_Update/cr
      -- CP-element group 228: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1243_sample_start_
      -- CP-element group 228: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1243_update_start_
      -- CP-element group 228: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1243_Sample/$entry
      -- CP-element group 228: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1243_Sample/rr
      -- CP-element group 228: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1243_Update/$entry
      -- CP-element group 228: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1243_Update/cr
      -- CP-element group 228: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1252_sample_start_
      -- CP-element group 228: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1252_update_start_
      -- CP-element group 228: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1252_Sample/$entry
      -- CP-element group 228: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1252_Sample/rr
      -- CP-element group 228: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1252_Update/$entry
      -- CP-element group 228: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1252_Update/cr
      -- CP-element group 228: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1261_update_start_
      -- CP-element group 228: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1261_Update/$entry
      -- CP-element group 228: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1261_Update/cr
      -- CP-element group 228: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1266_update_start_
      -- CP-element group 228: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1266_Update/$entry
      -- CP-element group 228: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1266_Update/cr
      -- CP-element group 228: 	 branch_block_stmt_436/ifx_xend_bbx_xnph_PhiReq/$entry
      -- CP-element group 228: 	 branch_block_stmt_436/ifx_xend_bbx_xnph_PhiReq/$exit
      -- CP-element group 228: 	 branch_block_stmt_436/merge_stmt_1215_PhiReqMerge
      -- CP-element group 228: 	 branch_block_stmt_436/merge_stmt_1215_PhiAck/$entry
      -- CP-element group 228: 	 branch_block_stmt_436/merge_stmt_1215_PhiAck/$exit
      -- CP-element group 228: 	 branch_block_stmt_436/merge_stmt_1215_PhiAck/dummy
      -- 
    if_choice_transition_2751_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 228_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1209_branch_ack_1, ack => convolution3D_CP_1120_elements(228)); -- 
    rr_2768_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2768_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(228), ack => type_cast_1230_inst_req_0); -- 
    cr_2773_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2773_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(228), ack => type_cast_1230_inst_req_1); -- 
    rr_2782_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2782_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(228), ack => type_cast_1234_inst_req_0); -- 
    cr_2787_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2787_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(228), ack => type_cast_1234_inst_req_1); -- 
    rr_2796_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2796_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(228), ack => type_cast_1243_inst_req_0); -- 
    cr_2801_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2801_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(228), ack => type_cast_1243_inst_req_1); -- 
    rr_2810_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2810_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(228), ack => type_cast_1252_inst_req_0); -- 
    cr_2815_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2815_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(228), ack => type_cast_1252_inst_req_1); -- 
    cr_2829_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2829_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(228), ack => type_cast_1261_inst_req_1); -- 
    cr_2843_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2843_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(228), ack => type_cast_1266_inst_req_1); -- 
    -- CP-element group 229:  transition  place  input  bypass 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	227 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	403 
    -- CP-element group 229:  members (6) 
      -- CP-element group 229: 	 branch_block_stmt_436/if_stmt_1209_else_link/$exit
      -- CP-element group 229: 	 branch_block_stmt_436/if_stmt_1209_else_link/else_choice_transition
      -- CP-element group 229: 	 branch_block_stmt_436/ifx_xend_forx_xend341
      -- CP-element group 229: 	 branch_block_stmt_436/ifx_xend_forx_xend341_PhiReq/$entry
      -- CP-element group 229: 	 branch_block_stmt_436/ifx_xend_forx_xend341_PhiReq/phi_stmt_1507/$entry
      -- CP-element group 229: 	 branch_block_stmt_436/ifx_xend_forx_xend341_PhiReq/phi_stmt_1507/phi_stmt_1507_sources/$entry
      -- 
    else_choice_transition_2755_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 229_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1209_branch_ack_0, ack => convolution3D_CP_1120_elements(229)); -- 
    -- CP-element group 230:  transition  input  bypass 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	228 
    -- CP-element group 230: successors 
    -- CP-element group 230:  members (3) 
      -- CP-element group 230: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1230_sample_completed_
      -- CP-element group 230: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1230_Sample/$exit
      -- CP-element group 230: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1230_Sample/ra
      -- 
    ra_2769_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 230_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1230_inst_ack_0, ack => convolution3D_CP_1120_elements(230)); -- 
    -- CP-element group 231:  transition  input  bypass 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	228 
    -- CP-element group 231: successors 
    -- CP-element group 231: 	238 
    -- CP-element group 231:  members (3) 
      -- CP-element group 231: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1230_update_completed_
      -- CP-element group 231: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1230_Update/$exit
      -- CP-element group 231: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1230_Update/ca
      -- 
    ca_2774_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 231_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1230_inst_ack_1, ack => convolution3D_CP_1120_elements(231)); -- 
    -- CP-element group 232:  transition  input  bypass 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	228 
    -- CP-element group 232: successors 
    -- CP-element group 232:  members (3) 
      -- CP-element group 232: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1234_sample_completed_
      -- CP-element group 232: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1234_Sample/$exit
      -- CP-element group 232: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1234_Sample/ra
      -- 
    ra_2783_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 232_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1234_inst_ack_0, ack => convolution3D_CP_1120_elements(232)); -- 
    -- CP-element group 233:  transition  input  bypass 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	228 
    -- CP-element group 233: successors 
    -- CP-element group 233: 	238 
    -- CP-element group 233:  members (3) 
      -- CP-element group 233: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1234_update_completed_
      -- CP-element group 233: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1234_Update/$exit
      -- CP-element group 233: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1234_Update/ca
      -- 
    ca_2788_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 233_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1234_inst_ack_1, ack => convolution3D_CP_1120_elements(233)); -- 
    -- CP-element group 234:  transition  input  bypass 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	228 
    -- CP-element group 234: successors 
    -- CP-element group 234:  members (3) 
      -- CP-element group 234: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1243_sample_completed_
      -- CP-element group 234: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1243_Sample/$exit
      -- CP-element group 234: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1243_Sample/ra
      -- 
    ra_2797_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 234_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1243_inst_ack_0, ack => convolution3D_CP_1120_elements(234)); -- 
    -- CP-element group 235:  transition  input  bypass 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	228 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	238 
    -- CP-element group 235:  members (3) 
      -- CP-element group 235: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1243_update_completed_
      -- CP-element group 235: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1243_Update/$exit
      -- CP-element group 235: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1243_Update/ca
      -- 
    ca_2802_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 235_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1243_inst_ack_1, ack => convolution3D_CP_1120_elements(235)); -- 
    -- CP-element group 236:  transition  input  bypass 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	228 
    -- CP-element group 236: successors 
    -- CP-element group 236:  members (3) 
      -- CP-element group 236: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1252_sample_completed_
      -- CP-element group 236: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1252_Sample/$exit
      -- CP-element group 236: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1252_Sample/ra
      -- 
    ra_2811_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 236_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1252_inst_ack_0, ack => convolution3D_CP_1120_elements(236)); -- 
    -- CP-element group 237:  transition  input  bypass 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	228 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	238 
    -- CP-element group 237:  members (3) 
      -- CP-element group 237: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1252_update_completed_
      -- CP-element group 237: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1252_Update/$exit
      -- CP-element group 237: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1252_Update/ca
      -- 
    ca_2816_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 237_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1252_inst_ack_1, ack => convolution3D_CP_1120_elements(237)); -- 
    -- CP-element group 238:  join  transition  output  bypass 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	231 
    -- CP-element group 238: 	233 
    -- CP-element group 238: 	235 
    -- CP-element group 238: 	237 
    -- CP-element group 238: successors 
    -- CP-element group 238: 	239 
    -- CP-element group 238:  members (3) 
      -- CP-element group 238: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1261_sample_start_
      -- CP-element group 238: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1261_Sample/$entry
      -- CP-element group 238: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1261_Sample/rr
      -- 
    rr_2824_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2824_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(238), ack => type_cast_1261_inst_req_0); -- 
    convolution3D_cp_element_group_238: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_238"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(231) & convolution3D_CP_1120_elements(233) & convolution3D_CP_1120_elements(235) & convolution3D_CP_1120_elements(237);
      gj_convolution3D_cp_element_group_238 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(238), clk => clk, reset => reset); --
    end block;
    -- CP-element group 239:  transition  input  bypass 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	238 
    -- CP-element group 239: successors 
    -- CP-element group 239:  members (3) 
      -- CP-element group 239: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1261_sample_completed_
      -- CP-element group 239: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1261_Sample/$exit
      -- CP-element group 239: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1261_Sample/ra
      -- 
    ra_2825_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 239_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1261_inst_ack_0, ack => convolution3D_CP_1120_elements(239)); -- 
    -- CP-element group 240:  transition  input  output  bypass 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	228 
    -- CP-element group 240: successors 
    -- CP-element group 240: 	241 
    -- CP-element group 240:  members (6) 
      -- CP-element group 240: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1261_update_completed_
      -- CP-element group 240: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1261_Update/$exit
      -- CP-element group 240: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1261_Update/ca
      -- CP-element group 240: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1266_sample_start_
      -- CP-element group 240: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1266_Sample/$entry
      -- CP-element group 240: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1266_Sample/rr
      -- 
    ca_2830_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 240_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1261_inst_ack_1, ack => convolution3D_CP_1120_elements(240)); -- 
    rr_2838_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2838_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(240), ack => type_cast_1266_inst_req_0); -- 
    -- CP-element group 241:  transition  input  bypass 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	240 
    -- CP-element group 241: successors 
    -- CP-element group 241:  members (3) 
      -- CP-element group 241: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1266_sample_completed_
      -- CP-element group 241: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1266_Sample/$exit
      -- CP-element group 241: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1266_Sample/ra
      -- 
    ra_2839_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 241_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1266_inst_ack_0, ack => convolution3D_CP_1120_elements(241)); -- 
    -- CP-element group 242:  transition  place  input  bypass 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	228 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	394 
    -- CP-element group 242:  members (9) 
      -- CP-element group 242: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286__exit__
      -- CP-element group 242: 	 branch_block_stmt_436/bbx_xnph_forx_xbody257
      -- CP-element group 242: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/$exit
      -- CP-element group 242: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1266_update_completed_
      -- CP-element group 242: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1266_Update/$exit
      -- CP-element group 242: 	 branch_block_stmt_436/assign_stmt_1221_to_assign_stmt_1286/type_cast_1266_Update/ca
      -- CP-element group 242: 	 branch_block_stmt_436/bbx_xnph_forx_xbody257_PhiReq/$entry
      -- CP-element group 242: 	 branch_block_stmt_436/bbx_xnph_forx_xbody257_PhiReq/phi_stmt_1289/$entry
      -- CP-element group 242: 	 branch_block_stmt_436/bbx_xnph_forx_xbody257_PhiReq/phi_stmt_1289/phi_stmt_1289_sources/$entry
      -- 
    ca_2844_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 242_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1266_inst_ack_1, ack => convolution3D_CP_1120_elements(242)); -- 
    -- CP-element group 243:  transition  input  bypass 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	399 
    -- CP-element group 243: successors 
    -- CP-element group 243: 	305 
    -- CP-element group 243:  members (3) 
      -- CP-element group 243: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/array_obj_ref_1301_final_index_sum_regn_sample_complete
      -- CP-element group 243: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/array_obj_ref_1301_final_index_sum_regn_Sample/$exit
      -- CP-element group 243: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/array_obj_ref_1301_final_index_sum_regn_Sample/ack
      -- 
    ack_2873_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 243_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1301_index_offset_ack_0, ack => convolution3D_CP_1120_elements(243)); -- 
    -- CP-element group 244:  transition  input  output  bypass 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	399 
    -- CP-element group 244: successors 
    -- CP-element group 244: 	245 
    -- CP-element group 244:  members (11) 
      -- CP-element group 244: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/addr_of_1302_sample_start_
      -- CP-element group 244: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/array_obj_ref_1301_root_address_calculated
      -- CP-element group 244: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/array_obj_ref_1301_offset_calculated
      -- CP-element group 244: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/array_obj_ref_1301_final_index_sum_regn_Update/$exit
      -- CP-element group 244: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/array_obj_ref_1301_final_index_sum_regn_Update/ack
      -- CP-element group 244: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/array_obj_ref_1301_base_plus_offset/$entry
      -- CP-element group 244: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/array_obj_ref_1301_base_plus_offset/$exit
      -- CP-element group 244: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/array_obj_ref_1301_base_plus_offset/sum_rename_req
      -- CP-element group 244: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/array_obj_ref_1301_base_plus_offset/sum_rename_ack
      -- CP-element group 244: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/addr_of_1302_request/$entry
      -- CP-element group 244: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/addr_of_1302_request/req
      -- 
    ack_2878_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 244_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1301_index_offset_ack_1, ack => convolution3D_CP_1120_elements(244)); -- 
    req_2887_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2887_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(244), ack => addr_of_1302_final_reg_req_0); -- 
    -- CP-element group 245:  transition  input  bypass 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	244 
    -- CP-element group 245: successors 
    -- CP-element group 245:  members (3) 
      -- CP-element group 245: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/addr_of_1302_sample_completed_
      -- CP-element group 245: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/addr_of_1302_request/$exit
      -- CP-element group 245: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/addr_of_1302_request/ack
      -- 
    ack_2888_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 245_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1302_final_reg_ack_0, ack => convolution3D_CP_1120_elements(245)); -- 
    -- CP-element group 246:  fork  transition  input  bypass 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	399 
    -- CP-element group 246: successors 
    -- CP-element group 246: 	302 
    -- CP-element group 246:  members (19) 
      -- CP-element group 246: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/addr_of_1302_update_completed_
      -- CP-element group 246: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/addr_of_1302_complete/$exit
      -- CP-element group 246: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/addr_of_1302_complete/ack
      -- CP-element group 246: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/ptr_deref_1462_base_address_calculated
      -- CP-element group 246: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/ptr_deref_1462_word_address_calculated
      -- CP-element group 246: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/ptr_deref_1462_root_address_calculated
      -- CP-element group 246: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/ptr_deref_1462_base_address_resized
      -- CP-element group 246: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/ptr_deref_1462_base_addr_resize/$entry
      -- CP-element group 246: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/ptr_deref_1462_base_addr_resize/$exit
      -- CP-element group 246: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/ptr_deref_1462_base_addr_resize/base_resize_req
      -- CP-element group 246: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/ptr_deref_1462_base_addr_resize/base_resize_ack
      -- CP-element group 246: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/ptr_deref_1462_base_plus_offset/$entry
      -- CP-element group 246: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/ptr_deref_1462_base_plus_offset/$exit
      -- CP-element group 246: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/ptr_deref_1462_base_plus_offset/sum_rename_req
      -- CP-element group 246: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/ptr_deref_1462_base_plus_offset/sum_rename_ack
      -- CP-element group 246: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/ptr_deref_1462_word_addrgen/$entry
      -- CP-element group 246: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/ptr_deref_1462_word_addrgen/$exit
      -- CP-element group 246: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/ptr_deref_1462_word_addrgen/root_register_req
      -- CP-element group 246: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/ptr_deref_1462_word_addrgen/root_register_ack
      -- 
    ack_2893_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 246_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1302_final_reg_ack_1, ack => convolution3D_CP_1120_elements(246)); -- 
    -- CP-element group 247:  transition  input  output  bypass 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	399 
    -- CP-element group 247: successors 
    -- CP-element group 247: 	248 
    -- CP-element group 247:  members (6) 
      -- CP-element group 247: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1305_sample_completed_
      -- CP-element group 247: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1305_update_start_
      -- CP-element group 247: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1305_Sample/$exit
      -- CP-element group 247: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1305_Sample/ra
      -- CP-element group 247: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1305_Update/$entry
      -- CP-element group 247: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1305_Update/cr
      -- 
    ra_2902_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 247_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1305_inst_ack_0, ack => convolution3D_CP_1120_elements(247)); -- 
    cr_2906_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2906_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(247), ack => RPIPE_maxpool_input_pipe_1305_inst_req_1); -- 
    -- CP-element group 248:  fork  transition  input  output  bypass 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	247 
    -- CP-element group 248: successors 
    -- CP-element group 248: 	249 
    -- CP-element group 248: 	251 
    -- CP-element group 248: 	253 
    -- CP-element group 248:  members (12) 
      -- CP-element group 248: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1305_update_completed_
      -- CP-element group 248: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1305_Update/$exit
      -- CP-element group 248: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1305_Update/ca
      -- CP-element group 248: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1307_sample_start_
      -- CP-element group 248: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1307_Sample/$entry
      -- CP-element group 248: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1307_Sample/req
      -- CP-element group 248: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1312_sample_start_
      -- CP-element group 248: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1312_Sample/$entry
      -- CP-element group 248: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1312_Sample/rr
      -- CP-element group 248: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1321_sample_start_
      -- CP-element group 248: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1321_Sample/$entry
      -- CP-element group 248: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1321_Sample/rr
      -- 
    ca_2907_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 248_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1305_inst_ack_1, ack => convolution3D_CP_1120_elements(248)); -- 
    req_2915_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2915_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(248), ack => WPIPE_maxpool_output_pipe_1307_inst_req_0); -- 
    rr_2929_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2929_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(248), ack => type_cast_1312_inst_req_0); -- 
    rr_2943_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2943_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(248), ack => RPIPE_maxpool_input_pipe_1321_inst_req_0); -- 
    -- CP-element group 249:  transition  input  output  bypass 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	248 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	250 
    -- CP-element group 249:  members (6) 
      -- CP-element group 249: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1307_sample_completed_
      -- CP-element group 249: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1307_update_start_
      -- CP-element group 249: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1307_Sample/$exit
      -- CP-element group 249: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1307_Sample/ack
      -- CP-element group 249: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1307_Update/$entry
      -- CP-element group 249: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1307_Update/req
      -- 
    ack_2916_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 249_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1307_inst_ack_0, ack => convolution3D_CP_1120_elements(249)); -- 
    req_2920_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2920_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(249), ack => WPIPE_maxpool_output_pipe_1307_inst_req_1); -- 
    -- CP-element group 250:  transition  input  bypass 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	249 
    -- CP-element group 250: successors 
    -- CP-element group 250: 	255 
    -- CP-element group 250:  members (3) 
      -- CP-element group 250: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1307_update_completed_
      -- CP-element group 250: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1307_Update/$exit
      -- CP-element group 250: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1307_Update/ack
      -- 
    ack_2921_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 250_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1307_inst_ack_1, ack => convolution3D_CP_1120_elements(250)); -- 
    -- CP-element group 251:  transition  input  bypass 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	248 
    -- CP-element group 251: successors 
    -- CP-element group 251:  members (3) 
      -- CP-element group 251: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1312_sample_completed_
      -- CP-element group 251: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1312_Sample/$exit
      -- CP-element group 251: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1312_Sample/ra
      -- 
    ra_2930_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 251_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1312_inst_ack_0, ack => convolution3D_CP_1120_elements(251)); -- 
    -- CP-element group 252:  transition  input  bypass 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	399 
    -- CP-element group 252: successors 
    -- CP-element group 252: 	302 
    -- CP-element group 252:  members (3) 
      -- CP-element group 252: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1312_update_completed_
      -- CP-element group 252: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1312_Update/$exit
      -- CP-element group 252: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1312_Update/ca
      -- 
    ca_2935_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 252_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1312_inst_ack_1, ack => convolution3D_CP_1120_elements(252)); -- 
    -- CP-element group 253:  transition  input  output  bypass 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	248 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	254 
    -- CP-element group 253:  members (6) 
      -- CP-element group 253: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1321_sample_completed_
      -- CP-element group 253: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1321_update_start_
      -- CP-element group 253: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1321_Sample/$exit
      -- CP-element group 253: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1321_Sample/ra
      -- CP-element group 253: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1321_Update/$entry
      -- CP-element group 253: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1321_Update/cr
      -- 
    ra_2944_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 253_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1321_inst_ack_0, ack => convolution3D_CP_1120_elements(253)); -- 
    cr_2948_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2948_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(253), ack => RPIPE_maxpool_input_pipe_1321_inst_req_1); -- 
    -- CP-element group 254:  fork  transition  input  output  bypass 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	253 
    -- CP-element group 254: successors 
    -- CP-element group 254: 	255 
    -- CP-element group 254: 	258 
    -- CP-element group 254: 	260 
    -- CP-element group 254:  members (9) 
      -- CP-element group 254: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1321_update_completed_
      -- CP-element group 254: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1321_Update/$exit
      -- CP-element group 254: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1321_Update/ca
      -- CP-element group 254: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1328_sample_start_
      -- CP-element group 254: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1328_Sample/$entry
      -- CP-element group 254: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1328_Sample/rr
      -- CP-element group 254: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1342_sample_start_
      -- CP-element group 254: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1342_Sample/$entry
      -- CP-element group 254: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1342_Sample/rr
      -- 
    ca_2949_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 254_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1321_inst_ack_1, ack => convolution3D_CP_1120_elements(254)); -- 
    rr_2971_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2971_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(254), ack => type_cast_1328_inst_req_0); -- 
    rr_2985_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2985_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(254), ack => RPIPE_maxpool_input_pipe_1342_inst_req_0); -- 
    -- CP-element group 255:  join  transition  output  bypass 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	250 
    -- CP-element group 255: 	254 
    -- CP-element group 255: successors 
    -- CP-element group 255: 	256 
    -- CP-element group 255:  members (3) 
      -- CP-element group 255: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1323_sample_start_
      -- CP-element group 255: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1323_Sample/$entry
      -- CP-element group 255: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1323_Sample/req
      -- 
    req_2957_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2957_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(255), ack => WPIPE_maxpool_output_pipe_1323_inst_req_0); -- 
    convolution3D_cp_element_group_255: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_255"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(250) & convolution3D_CP_1120_elements(254);
      gj_convolution3D_cp_element_group_255 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(255), clk => clk, reset => reset); --
    end block;
    -- CP-element group 256:  transition  input  output  bypass 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	255 
    -- CP-element group 256: successors 
    -- CP-element group 256: 	257 
    -- CP-element group 256:  members (6) 
      -- CP-element group 256: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1323_sample_completed_
      -- CP-element group 256: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1323_update_start_
      -- CP-element group 256: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1323_Sample/$exit
      -- CP-element group 256: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1323_Sample/ack
      -- CP-element group 256: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1323_Update/$entry
      -- CP-element group 256: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1323_Update/req
      -- 
    ack_2958_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 256_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1323_inst_ack_0, ack => convolution3D_CP_1120_elements(256)); -- 
    req_2962_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2962_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(256), ack => WPIPE_maxpool_output_pipe_1323_inst_req_1); -- 
    -- CP-element group 257:  transition  input  bypass 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	256 
    -- CP-element group 257: successors 
    -- CP-element group 257: 	262 
    -- CP-element group 257:  members (3) 
      -- CP-element group 257: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1323_update_completed_
      -- CP-element group 257: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1323_Update/$exit
      -- CP-element group 257: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1323_Update/ack
      -- 
    ack_2963_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 257_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1323_inst_ack_1, ack => convolution3D_CP_1120_elements(257)); -- 
    -- CP-element group 258:  transition  input  bypass 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	254 
    -- CP-element group 258: successors 
    -- CP-element group 258:  members (3) 
      -- CP-element group 258: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1328_sample_completed_
      -- CP-element group 258: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1328_Sample/$exit
      -- CP-element group 258: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1328_Sample/ra
      -- 
    ra_2972_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 258_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1328_inst_ack_0, ack => convolution3D_CP_1120_elements(258)); -- 
    -- CP-element group 259:  transition  input  bypass 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	399 
    -- CP-element group 259: successors 
    -- CP-element group 259: 	302 
    -- CP-element group 259:  members (3) 
      -- CP-element group 259: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1328_update_completed_
      -- CP-element group 259: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1328_Update/$exit
      -- CP-element group 259: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1328_Update/ca
      -- 
    ca_2977_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 259_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1328_inst_ack_1, ack => convolution3D_CP_1120_elements(259)); -- 
    -- CP-element group 260:  transition  input  output  bypass 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	254 
    -- CP-element group 260: successors 
    -- CP-element group 260: 	261 
    -- CP-element group 260:  members (6) 
      -- CP-element group 260: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1342_sample_completed_
      -- CP-element group 260: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1342_update_start_
      -- CP-element group 260: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1342_Sample/$exit
      -- CP-element group 260: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1342_Sample/ra
      -- CP-element group 260: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1342_Update/$entry
      -- CP-element group 260: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1342_Update/cr
      -- 
    ra_2986_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 260_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1342_inst_ack_0, ack => convolution3D_CP_1120_elements(260)); -- 
    cr_2990_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2990_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(260), ack => RPIPE_maxpool_input_pipe_1342_inst_req_1); -- 
    -- CP-element group 261:  fork  transition  input  output  bypass 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	260 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	262 
    -- CP-element group 261: 	265 
    -- CP-element group 261: 	267 
    -- CP-element group 261:  members (9) 
      -- CP-element group 261: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1342_update_completed_
      -- CP-element group 261: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1342_Update/$exit
      -- CP-element group 261: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1342_Update/ca
      -- CP-element group 261: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1349_sample_start_
      -- CP-element group 261: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1349_Sample/$entry
      -- CP-element group 261: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1349_Sample/rr
      -- CP-element group 261: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1363_sample_start_
      -- CP-element group 261: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1363_Sample/$entry
      -- CP-element group 261: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1363_Sample/rr
      -- 
    ca_2991_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 261_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1342_inst_ack_1, ack => convolution3D_CP_1120_elements(261)); -- 
    rr_3013_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3013_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(261), ack => type_cast_1349_inst_req_0); -- 
    rr_3027_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3027_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(261), ack => RPIPE_maxpool_input_pipe_1363_inst_req_0); -- 
    -- CP-element group 262:  join  transition  output  bypass 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	257 
    -- CP-element group 262: 	261 
    -- CP-element group 262: successors 
    -- CP-element group 262: 	263 
    -- CP-element group 262:  members (3) 
      -- CP-element group 262: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1344_sample_start_
      -- CP-element group 262: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1344_Sample/$entry
      -- CP-element group 262: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1344_Sample/req
      -- 
    req_2999_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2999_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(262), ack => WPIPE_maxpool_output_pipe_1344_inst_req_0); -- 
    convolution3D_cp_element_group_262: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_262"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(257) & convolution3D_CP_1120_elements(261);
      gj_convolution3D_cp_element_group_262 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(262), clk => clk, reset => reset); --
    end block;
    -- CP-element group 263:  transition  input  output  bypass 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	262 
    -- CP-element group 263: successors 
    -- CP-element group 263: 	264 
    -- CP-element group 263:  members (6) 
      -- CP-element group 263: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1344_sample_completed_
      -- CP-element group 263: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1344_update_start_
      -- CP-element group 263: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1344_Sample/$exit
      -- CP-element group 263: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1344_Sample/ack
      -- CP-element group 263: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1344_Update/$entry
      -- CP-element group 263: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1344_Update/req
      -- 
    ack_3000_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 263_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1344_inst_ack_0, ack => convolution3D_CP_1120_elements(263)); -- 
    req_3004_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3004_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(263), ack => WPIPE_maxpool_output_pipe_1344_inst_req_1); -- 
    -- CP-element group 264:  transition  input  bypass 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	263 
    -- CP-element group 264: successors 
    -- CP-element group 264: 	269 
    -- CP-element group 264:  members (3) 
      -- CP-element group 264: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1344_update_completed_
      -- CP-element group 264: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1344_Update/$exit
      -- CP-element group 264: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1344_Update/ack
      -- 
    ack_3005_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 264_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1344_inst_ack_1, ack => convolution3D_CP_1120_elements(264)); -- 
    -- CP-element group 265:  transition  input  bypass 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	261 
    -- CP-element group 265: successors 
    -- CP-element group 265:  members (3) 
      -- CP-element group 265: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1349_sample_completed_
      -- CP-element group 265: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1349_Sample/$exit
      -- CP-element group 265: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1349_Sample/ra
      -- 
    ra_3014_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 265_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1349_inst_ack_0, ack => convolution3D_CP_1120_elements(265)); -- 
    -- CP-element group 266:  transition  input  bypass 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	399 
    -- CP-element group 266: successors 
    -- CP-element group 266: 	302 
    -- CP-element group 266:  members (3) 
      -- CP-element group 266: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1349_update_completed_
      -- CP-element group 266: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1349_Update/$exit
      -- CP-element group 266: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1349_Update/ca
      -- 
    ca_3019_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 266_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1349_inst_ack_1, ack => convolution3D_CP_1120_elements(266)); -- 
    -- CP-element group 267:  transition  input  output  bypass 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	261 
    -- CP-element group 267: successors 
    -- CP-element group 267: 	268 
    -- CP-element group 267:  members (6) 
      -- CP-element group 267: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1363_sample_completed_
      -- CP-element group 267: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1363_update_start_
      -- CP-element group 267: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1363_Sample/$exit
      -- CP-element group 267: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1363_Sample/ra
      -- CP-element group 267: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1363_Update/$entry
      -- CP-element group 267: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1363_Update/cr
      -- 
    ra_3028_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 267_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1363_inst_ack_0, ack => convolution3D_CP_1120_elements(267)); -- 
    cr_3032_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3032_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(267), ack => RPIPE_maxpool_input_pipe_1363_inst_req_1); -- 
    -- CP-element group 268:  fork  transition  input  output  bypass 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	267 
    -- CP-element group 268: successors 
    -- CP-element group 268: 	269 
    -- CP-element group 268: 	272 
    -- CP-element group 268: 	274 
    -- CP-element group 268:  members (9) 
      -- CP-element group 268: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1363_update_completed_
      -- CP-element group 268: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1363_Update/$exit
      -- CP-element group 268: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1363_Update/ca
      -- CP-element group 268: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1370_sample_start_
      -- CP-element group 268: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1370_Sample/$entry
      -- CP-element group 268: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1370_Sample/rr
      -- CP-element group 268: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1384_sample_start_
      -- CP-element group 268: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1384_Sample/$entry
      -- CP-element group 268: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1384_Sample/rr
      -- 
    ca_3033_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 268_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1363_inst_ack_1, ack => convolution3D_CP_1120_elements(268)); -- 
    rr_3055_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3055_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(268), ack => type_cast_1370_inst_req_0); -- 
    rr_3069_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3069_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(268), ack => RPIPE_maxpool_input_pipe_1384_inst_req_0); -- 
    -- CP-element group 269:  join  transition  output  bypass 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: 	264 
    -- CP-element group 269: 	268 
    -- CP-element group 269: successors 
    -- CP-element group 269: 	270 
    -- CP-element group 269:  members (3) 
      -- CP-element group 269: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1365_sample_start_
      -- CP-element group 269: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1365_Sample/$entry
      -- CP-element group 269: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1365_Sample/req
      -- 
    req_3041_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3041_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(269), ack => WPIPE_maxpool_output_pipe_1365_inst_req_0); -- 
    convolution3D_cp_element_group_269: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_269"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(264) & convolution3D_CP_1120_elements(268);
      gj_convolution3D_cp_element_group_269 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(269), clk => clk, reset => reset); --
    end block;
    -- CP-element group 270:  transition  input  output  bypass 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	269 
    -- CP-element group 270: successors 
    -- CP-element group 270: 	271 
    -- CP-element group 270:  members (6) 
      -- CP-element group 270: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1365_sample_completed_
      -- CP-element group 270: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1365_update_start_
      -- CP-element group 270: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1365_Sample/$exit
      -- CP-element group 270: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1365_Sample/ack
      -- CP-element group 270: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1365_Update/$entry
      -- CP-element group 270: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1365_Update/req
      -- 
    ack_3042_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 270_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1365_inst_ack_0, ack => convolution3D_CP_1120_elements(270)); -- 
    req_3046_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3046_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(270), ack => WPIPE_maxpool_output_pipe_1365_inst_req_1); -- 
    -- CP-element group 271:  transition  input  bypass 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	270 
    -- CP-element group 271: successors 
    -- CP-element group 271: 	276 
    -- CP-element group 271:  members (3) 
      -- CP-element group 271: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1365_update_completed_
      -- CP-element group 271: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1365_Update/$exit
      -- CP-element group 271: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1365_Update/ack
      -- 
    ack_3047_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 271_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1365_inst_ack_1, ack => convolution3D_CP_1120_elements(271)); -- 
    -- CP-element group 272:  transition  input  bypass 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	268 
    -- CP-element group 272: successors 
    -- CP-element group 272:  members (3) 
      -- CP-element group 272: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1370_sample_completed_
      -- CP-element group 272: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1370_Sample/$exit
      -- CP-element group 272: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1370_Sample/ra
      -- 
    ra_3056_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 272_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1370_inst_ack_0, ack => convolution3D_CP_1120_elements(272)); -- 
    -- CP-element group 273:  transition  input  bypass 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: 	399 
    -- CP-element group 273: successors 
    -- CP-element group 273: 	302 
    -- CP-element group 273:  members (3) 
      -- CP-element group 273: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1370_update_completed_
      -- CP-element group 273: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1370_Update/$exit
      -- CP-element group 273: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1370_Update/ca
      -- 
    ca_3061_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 273_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1370_inst_ack_1, ack => convolution3D_CP_1120_elements(273)); -- 
    -- CP-element group 274:  transition  input  output  bypass 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	268 
    -- CP-element group 274: successors 
    -- CP-element group 274: 	275 
    -- CP-element group 274:  members (6) 
      -- CP-element group 274: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1384_sample_completed_
      -- CP-element group 274: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1384_update_start_
      -- CP-element group 274: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1384_Sample/$exit
      -- CP-element group 274: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1384_Sample/ra
      -- CP-element group 274: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1384_Update/$entry
      -- CP-element group 274: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1384_Update/cr
      -- 
    ra_3070_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 274_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1384_inst_ack_0, ack => convolution3D_CP_1120_elements(274)); -- 
    cr_3074_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3074_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(274), ack => RPIPE_maxpool_input_pipe_1384_inst_req_1); -- 
    -- CP-element group 275:  fork  transition  input  output  bypass 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	274 
    -- CP-element group 275: successors 
    -- CP-element group 275: 	276 
    -- CP-element group 275: 	279 
    -- CP-element group 275: 	281 
    -- CP-element group 275:  members (9) 
      -- CP-element group 275: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1384_update_completed_
      -- CP-element group 275: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1384_Update/$exit
      -- CP-element group 275: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1384_Update/ca
      -- CP-element group 275: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1391_sample_start_
      -- CP-element group 275: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1391_Sample/$entry
      -- CP-element group 275: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1391_Sample/rr
      -- CP-element group 275: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1405_sample_start_
      -- CP-element group 275: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1405_Sample/$entry
      -- CP-element group 275: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1405_Sample/rr
      -- 
    ca_3075_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 275_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1384_inst_ack_1, ack => convolution3D_CP_1120_elements(275)); -- 
    rr_3097_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3097_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(275), ack => type_cast_1391_inst_req_0); -- 
    rr_3111_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3111_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(275), ack => RPIPE_maxpool_input_pipe_1405_inst_req_0); -- 
    -- CP-element group 276:  join  transition  output  bypass 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	271 
    -- CP-element group 276: 	275 
    -- CP-element group 276: successors 
    -- CP-element group 276: 	277 
    -- CP-element group 276:  members (3) 
      -- CP-element group 276: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1386_sample_start_
      -- CP-element group 276: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1386_Sample/$entry
      -- CP-element group 276: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1386_Sample/req
      -- 
    req_3083_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3083_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(276), ack => WPIPE_maxpool_output_pipe_1386_inst_req_0); -- 
    convolution3D_cp_element_group_276: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_276"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(271) & convolution3D_CP_1120_elements(275);
      gj_convolution3D_cp_element_group_276 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(276), clk => clk, reset => reset); --
    end block;
    -- CP-element group 277:  transition  input  output  bypass 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	276 
    -- CP-element group 277: successors 
    -- CP-element group 277: 	278 
    -- CP-element group 277:  members (6) 
      -- CP-element group 277: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1386_sample_completed_
      -- CP-element group 277: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1386_update_start_
      -- CP-element group 277: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1386_Sample/$exit
      -- CP-element group 277: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1386_Sample/ack
      -- CP-element group 277: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1386_Update/$entry
      -- CP-element group 277: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1386_Update/req
      -- 
    ack_3084_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 277_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1386_inst_ack_0, ack => convolution3D_CP_1120_elements(277)); -- 
    req_3088_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3088_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(277), ack => WPIPE_maxpool_output_pipe_1386_inst_req_1); -- 
    -- CP-element group 278:  transition  input  bypass 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	277 
    -- CP-element group 278: successors 
    -- CP-element group 278: 	283 
    -- CP-element group 278:  members (3) 
      -- CP-element group 278: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1386_update_completed_
      -- CP-element group 278: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1386_Update/$exit
      -- CP-element group 278: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1386_Update/ack
      -- 
    ack_3089_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 278_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1386_inst_ack_1, ack => convolution3D_CP_1120_elements(278)); -- 
    -- CP-element group 279:  transition  input  bypass 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	275 
    -- CP-element group 279: successors 
    -- CP-element group 279:  members (3) 
      -- CP-element group 279: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1391_sample_completed_
      -- CP-element group 279: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1391_Sample/$exit
      -- CP-element group 279: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1391_Sample/ra
      -- 
    ra_3098_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 279_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1391_inst_ack_0, ack => convolution3D_CP_1120_elements(279)); -- 
    -- CP-element group 280:  transition  input  bypass 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	399 
    -- CP-element group 280: successors 
    -- CP-element group 280: 	302 
    -- CP-element group 280:  members (3) 
      -- CP-element group 280: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1391_update_completed_
      -- CP-element group 280: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1391_Update/$exit
      -- CP-element group 280: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1391_Update/ca
      -- 
    ca_3103_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 280_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1391_inst_ack_1, ack => convolution3D_CP_1120_elements(280)); -- 
    -- CP-element group 281:  transition  input  output  bypass 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	275 
    -- CP-element group 281: successors 
    -- CP-element group 281: 	282 
    -- CP-element group 281:  members (6) 
      -- CP-element group 281: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1405_sample_completed_
      -- CP-element group 281: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1405_update_start_
      -- CP-element group 281: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1405_Sample/$exit
      -- CP-element group 281: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1405_Sample/ra
      -- CP-element group 281: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1405_Update/$entry
      -- CP-element group 281: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1405_Update/cr
      -- 
    ra_3112_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 281_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1405_inst_ack_0, ack => convolution3D_CP_1120_elements(281)); -- 
    cr_3116_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3116_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(281), ack => RPIPE_maxpool_input_pipe_1405_inst_req_1); -- 
    -- CP-element group 282:  fork  transition  input  output  bypass 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	281 
    -- CP-element group 282: successors 
    -- CP-element group 282: 	283 
    -- CP-element group 282: 	286 
    -- CP-element group 282: 	288 
    -- CP-element group 282:  members (9) 
      -- CP-element group 282: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1405_update_completed_
      -- CP-element group 282: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1405_Update/$exit
      -- CP-element group 282: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1405_Update/ca
      -- CP-element group 282: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1412_sample_start_
      -- CP-element group 282: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1412_Sample/$entry
      -- CP-element group 282: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1412_Sample/rr
      -- CP-element group 282: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1426_sample_start_
      -- CP-element group 282: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1426_Sample/$entry
      -- CP-element group 282: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1426_Sample/rr
      -- 
    ca_3117_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 282_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1405_inst_ack_1, ack => convolution3D_CP_1120_elements(282)); -- 
    rr_3139_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3139_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(282), ack => type_cast_1412_inst_req_0); -- 
    rr_3153_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3153_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(282), ack => RPIPE_maxpool_input_pipe_1426_inst_req_0); -- 
    -- CP-element group 283:  join  transition  output  bypass 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: 	278 
    -- CP-element group 283: 	282 
    -- CP-element group 283: successors 
    -- CP-element group 283: 	284 
    -- CP-element group 283:  members (3) 
      -- CP-element group 283: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1407_sample_start_
      -- CP-element group 283: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1407_Sample/$entry
      -- CP-element group 283: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1407_Sample/req
      -- 
    req_3125_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3125_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(283), ack => WPIPE_maxpool_output_pipe_1407_inst_req_0); -- 
    convolution3D_cp_element_group_283: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_283"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(278) & convolution3D_CP_1120_elements(282);
      gj_convolution3D_cp_element_group_283 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(283), clk => clk, reset => reset); --
    end block;
    -- CP-element group 284:  transition  input  output  bypass 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	283 
    -- CP-element group 284: successors 
    -- CP-element group 284: 	285 
    -- CP-element group 284:  members (6) 
      -- CP-element group 284: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1407_sample_completed_
      -- CP-element group 284: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1407_update_start_
      -- CP-element group 284: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1407_Sample/$exit
      -- CP-element group 284: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1407_Sample/ack
      -- CP-element group 284: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1407_Update/$entry
      -- CP-element group 284: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1407_Update/req
      -- 
    ack_3126_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 284_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1407_inst_ack_0, ack => convolution3D_CP_1120_elements(284)); -- 
    req_3130_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3130_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(284), ack => WPIPE_maxpool_output_pipe_1407_inst_req_1); -- 
    -- CP-element group 285:  transition  input  bypass 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: 	284 
    -- CP-element group 285: successors 
    -- CP-element group 285: 	290 
    -- CP-element group 285:  members (3) 
      -- CP-element group 285: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1407_update_completed_
      -- CP-element group 285: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1407_Update/$exit
      -- CP-element group 285: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1407_Update/ack
      -- 
    ack_3131_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 285_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1407_inst_ack_1, ack => convolution3D_CP_1120_elements(285)); -- 
    -- CP-element group 286:  transition  input  bypass 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	282 
    -- CP-element group 286: successors 
    -- CP-element group 286:  members (3) 
      -- CP-element group 286: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1412_sample_completed_
      -- CP-element group 286: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1412_Sample/$exit
      -- CP-element group 286: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1412_Sample/ra
      -- 
    ra_3140_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 286_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1412_inst_ack_0, ack => convolution3D_CP_1120_elements(286)); -- 
    -- CP-element group 287:  transition  input  bypass 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	399 
    -- CP-element group 287: successors 
    -- CP-element group 287: 	302 
    -- CP-element group 287:  members (3) 
      -- CP-element group 287: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1412_update_completed_
      -- CP-element group 287: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1412_Update/$exit
      -- CP-element group 287: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1412_Update/ca
      -- 
    ca_3145_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 287_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1412_inst_ack_1, ack => convolution3D_CP_1120_elements(287)); -- 
    -- CP-element group 288:  transition  input  output  bypass 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	282 
    -- CP-element group 288: successors 
    -- CP-element group 288: 	289 
    -- CP-element group 288:  members (6) 
      -- CP-element group 288: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1426_sample_completed_
      -- CP-element group 288: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1426_update_start_
      -- CP-element group 288: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1426_Sample/$exit
      -- CP-element group 288: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1426_Sample/ra
      -- CP-element group 288: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1426_Update/$entry
      -- CP-element group 288: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1426_Update/cr
      -- 
    ra_3154_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 288_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1426_inst_ack_0, ack => convolution3D_CP_1120_elements(288)); -- 
    cr_3158_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3158_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(288), ack => RPIPE_maxpool_input_pipe_1426_inst_req_1); -- 
    -- CP-element group 289:  fork  transition  input  output  bypass 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: 	288 
    -- CP-element group 289: successors 
    -- CP-element group 289: 	290 
    -- CP-element group 289: 	293 
    -- CP-element group 289: 	295 
    -- CP-element group 289:  members (9) 
      -- CP-element group 289: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1426_update_completed_
      -- CP-element group 289: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1426_Update/$exit
      -- CP-element group 289: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1426_Update/ca
      -- CP-element group 289: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1433_sample_start_
      -- CP-element group 289: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1433_Sample/$entry
      -- CP-element group 289: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1433_Sample/rr
      -- CP-element group 289: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1447_sample_start_
      -- CP-element group 289: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1447_Sample/$entry
      -- CP-element group 289: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1447_Sample/rr
      -- 
    ca_3159_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 289_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1426_inst_ack_1, ack => convolution3D_CP_1120_elements(289)); -- 
    rr_3181_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3181_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(289), ack => type_cast_1433_inst_req_0); -- 
    rr_3195_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3195_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(289), ack => RPIPE_maxpool_input_pipe_1447_inst_req_0); -- 
    -- CP-element group 290:  join  transition  output  bypass 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: 	285 
    -- CP-element group 290: 	289 
    -- CP-element group 290: successors 
    -- CP-element group 290: 	291 
    -- CP-element group 290:  members (3) 
      -- CP-element group 290: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1428_sample_start_
      -- CP-element group 290: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1428_Sample/$entry
      -- CP-element group 290: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1428_Sample/req
      -- 
    req_3167_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3167_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(290), ack => WPIPE_maxpool_output_pipe_1428_inst_req_0); -- 
    convolution3D_cp_element_group_290: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_290"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(285) & convolution3D_CP_1120_elements(289);
      gj_convolution3D_cp_element_group_290 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(290), clk => clk, reset => reset); --
    end block;
    -- CP-element group 291:  transition  input  output  bypass 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	290 
    -- CP-element group 291: successors 
    -- CP-element group 291: 	292 
    -- CP-element group 291:  members (6) 
      -- CP-element group 291: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1428_sample_completed_
      -- CP-element group 291: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1428_update_start_
      -- CP-element group 291: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1428_Sample/$exit
      -- CP-element group 291: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1428_Sample/ack
      -- CP-element group 291: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1428_Update/$entry
      -- CP-element group 291: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1428_Update/req
      -- 
    ack_3168_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 291_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1428_inst_ack_0, ack => convolution3D_CP_1120_elements(291)); -- 
    req_3172_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3172_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(291), ack => WPIPE_maxpool_output_pipe_1428_inst_req_1); -- 
    -- CP-element group 292:  transition  input  bypass 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	291 
    -- CP-element group 292: successors 
    -- CP-element group 292: 	297 
    -- CP-element group 292:  members (3) 
      -- CP-element group 292: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1428_update_completed_
      -- CP-element group 292: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1428_Update/$exit
      -- CP-element group 292: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1428_Update/ack
      -- 
    ack_3173_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 292_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1428_inst_ack_1, ack => convolution3D_CP_1120_elements(292)); -- 
    -- CP-element group 293:  transition  input  bypass 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: 	289 
    -- CP-element group 293: successors 
    -- CP-element group 293:  members (3) 
      -- CP-element group 293: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1433_sample_completed_
      -- CP-element group 293: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1433_Sample/$exit
      -- CP-element group 293: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1433_Sample/ra
      -- 
    ra_3182_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 293_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1433_inst_ack_0, ack => convolution3D_CP_1120_elements(293)); -- 
    -- CP-element group 294:  transition  input  bypass 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: 	399 
    -- CP-element group 294: successors 
    -- CP-element group 294: 	302 
    -- CP-element group 294:  members (3) 
      -- CP-element group 294: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1433_update_completed_
      -- CP-element group 294: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1433_Update/$exit
      -- CP-element group 294: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1433_Update/ca
      -- 
    ca_3187_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 294_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1433_inst_ack_1, ack => convolution3D_CP_1120_elements(294)); -- 
    -- CP-element group 295:  transition  input  output  bypass 
    -- CP-element group 295: predecessors 
    -- CP-element group 295: 	289 
    -- CP-element group 295: successors 
    -- CP-element group 295: 	296 
    -- CP-element group 295:  members (6) 
      -- CP-element group 295: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1447_sample_completed_
      -- CP-element group 295: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1447_update_start_
      -- CP-element group 295: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1447_Sample/$exit
      -- CP-element group 295: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1447_Sample/ra
      -- CP-element group 295: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1447_Update/$entry
      -- CP-element group 295: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1447_Update/cr
      -- 
    ra_3196_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 295_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1447_inst_ack_0, ack => convolution3D_CP_1120_elements(295)); -- 
    cr_3200_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3200_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(295), ack => RPIPE_maxpool_input_pipe_1447_inst_req_1); -- 
    -- CP-element group 296:  fork  transition  input  output  bypass 
    -- CP-element group 296: predecessors 
    -- CP-element group 296: 	295 
    -- CP-element group 296: successors 
    -- CP-element group 296: 	297 
    -- CP-element group 296: 	300 
    -- CP-element group 296:  members (6) 
      -- CP-element group 296: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1447_update_completed_
      -- CP-element group 296: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1447_Update/$exit
      -- CP-element group 296: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1447_Update/ca
      -- CP-element group 296: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1454_sample_start_
      -- CP-element group 296: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1454_Sample/$entry
      -- CP-element group 296: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1454_Sample/rr
      -- 
    ca_3201_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 296_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1447_inst_ack_1, ack => convolution3D_CP_1120_elements(296)); -- 
    rr_3223_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3223_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(296), ack => type_cast_1454_inst_req_0); -- 
    -- CP-element group 297:  join  transition  output  bypass 
    -- CP-element group 297: predecessors 
    -- CP-element group 297: 	292 
    -- CP-element group 297: 	296 
    -- CP-element group 297: successors 
    -- CP-element group 297: 	298 
    -- CP-element group 297:  members (3) 
      -- CP-element group 297: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1449_sample_start_
      -- CP-element group 297: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1449_Sample/$entry
      -- CP-element group 297: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1449_Sample/req
      -- 
    req_3209_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3209_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(297), ack => WPIPE_maxpool_output_pipe_1449_inst_req_0); -- 
    convolution3D_cp_element_group_297: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_297"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(292) & convolution3D_CP_1120_elements(296);
      gj_convolution3D_cp_element_group_297 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(297), clk => clk, reset => reset); --
    end block;
    -- CP-element group 298:  transition  input  output  bypass 
    -- CP-element group 298: predecessors 
    -- CP-element group 298: 	297 
    -- CP-element group 298: successors 
    -- CP-element group 298: 	299 
    -- CP-element group 298:  members (6) 
      -- CP-element group 298: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1449_sample_completed_
      -- CP-element group 298: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1449_update_start_
      -- CP-element group 298: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1449_Sample/$exit
      -- CP-element group 298: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1449_Sample/ack
      -- CP-element group 298: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1449_Update/$entry
      -- CP-element group 298: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1449_Update/req
      -- 
    ack_3210_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 298_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1449_inst_ack_0, ack => convolution3D_CP_1120_elements(298)); -- 
    req_3214_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3214_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(298), ack => WPIPE_maxpool_output_pipe_1449_inst_req_1); -- 
    -- CP-element group 299:  transition  input  bypass 
    -- CP-element group 299: predecessors 
    -- CP-element group 299: 	298 
    -- CP-element group 299: successors 
    -- CP-element group 299: 	305 
    -- CP-element group 299:  members (3) 
      -- CP-element group 299: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1449_update_completed_
      -- CP-element group 299: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1449_Update/$exit
      -- CP-element group 299: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/WPIPE_maxpool_output_pipe_1449_Update/ack
      -- 
    ack_3215_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 299_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1449_inst_ack_1, ack => convolution3D_CP_1120_elements(299)); -- 
    -- CP-element group 300:  transition  input  bypass 
    -- CP-element group 300: predecessors 
    -- CP-element group 300: 	296 
    -- CP-element group 300: successors 
    -- CP-element group 300:  members (3) 
      -- CP-element group 300: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1454_sample_completed_
      -- CP-element group 300: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1454_Sample/$exit
      -- CP-element group 300: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1454_Sample/ra
      -- 
    ra_3224_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 300_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1454_inst_ack_0, ack => convolution3D_CP_1120_elements(300)); -- 
    -- CP-element group 301:  transition  input  bypass 
    -- CP-element group 301: predecessors 
    -- CP-element group 301: 	399 
    -- CP-element group 301: successors 
    -- CP-element group 301: 	302 
    -- CP-element group 301:  members (3) 
      -- CP-element group 301: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1454_update_completed_
      -- CP-element group 301: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1454_Update/$exit
      -- CP-element group 301: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1454_Update/ca
      -- 
    ca_3229_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 301_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1454_inst_ack_1, ack => convolution3D_CP_1120_elements(301)); -- 
    -- CP-element group 302:  join  transition  output  bypass 
    -- CP-element group 302: predecessors 
    -- CP-element group 302: 	246 
    -- CP-element group 302: 	252 
    -- CP-element group 302: 	259 
    -- CP-element group 302: 	266 
    -- CP-element group 302: 	273 
    -- CP-element group 302: 	280 
    -- CP-element group 302: 	287 
    -- CP-element group 302: 	294 
    -- CP-element group 302: 	301 
    -- CP-element group 302: successors 
    -- CP-element group 302: 	303 
    -- CP-element group 302:  members (9) 
      -- CP-element group 302: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/ptr_deref_1462_sample_start_
      -- CP-element group 302: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/ptr_deref_1462_Sample/$entry
      -- CP-element group 302: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/ptr_deref_1462_Sample/ptr_deref_1462_Split/$entry
      -- CP-element group 302: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/ptr_deref_1462_Sample/ptr_deref_1462_Split/$exit
      -- CP-element group 302: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/ptr_deref_1462_Sample/ptr_deref_1462_Split/split_req
      -- CP-element group 302: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/ptr_deref_1462_Sample/ptr_deref_1462_Split/split_ack
      -- CP-element group 302: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/ptr_deref_1462_Sample/word_access_start/$entry
      -- CP-element group 302: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/ptr_deref_1462_Sample/word_access_start/word_0/$entry
      -- CP-element group 302: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/ptr_deref_1462_Sample/word_access_start/word_0/rr
      -- 
    rr_3267_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3267_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(302), ack => ptr_deref_1462_store_0_req_0); -- 
    convolution3D_cp_element_group_302: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_302"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(246) & convolution3D_CP_1120_elements(252) & convolution3D_CP_1120_elements(259) & convolution3D_CP_1120_elements(266) & convolution3D_CP_1120_elements(273) & convolution3D_CP_1120_elements(280) & convolution3D_CP_1120_elements(287) & convolution3D_CP_1120_elements(294) & convolution3D_CP_1120_elements(301);
      gj_convolution3D_cp_element_group_302 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(302), clk => clk, reset => reset); --
    end block;
    -- CP-element group 303:  transition  input  bypass 
    -- CP-element group 303: predecessors 
    -- CP-element group 303: 	302 
    -- CP-element group 303: successors 
    -- CP-element group 303:  members (5) 
      -- CP-element group 303: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/ptr_deref_1462_sample_completed_
      -- CP-element group 303: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/ptr_deref_1462_Sample/$exit
      -- CP-element group 303: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/ptr_deref_1462_Sample/word_access_start/$exit
      -- CP-element group 303: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/ptr_deref_1462_Sample/word_access_start/word_0/$exit
      -- CP-element group 303: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/ptr_deref_1462_Sample/word_access_start/word_0/ra
      -- 
    ra_3268_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 303_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1462_store_0_ack_0, ack => convolution3D_CP_1120_elements(303)); -- 
    -- CP-element group 304:  transition  input  bypass 
    -- CP-element group 304: predecessors 
    -- CP-element group 304: 	399 
    -- CP-element group 304: successors 
    -- CP-element group 304: 	305 
    -- CP-element group 304:  members (5) 
      -- CP-element group 304: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/ptr_deref_1462_update_completed_
      -- CP-element group 304: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/ptr_deref_1462_Update/$exit
      -- CP-element group 304: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/ptr_deref_1462_Update/word_access_complete/$exit
      -- CP-element group 304: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/ptr_deref_1462_Update/word_access_complete/word_0/$exit
      -- CP-element group 304: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/ptr_deref_1462_Update/word_access_complete/word_0/ca
      -- 
    ca_3279_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 304_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1462_store_0_ack_1, ack => convolution3D_CP_1120_elements(304)); -- 
    -- CP-element group 305:  branch  join  transition  place  output  bypass 
    -- CP-element group 305: predecessors 
    -- CP-element group 305: 	243 
    -- CP-element group 305: 	299 
    -- CP-element group 305: 	304 
    -- CP-element group 305: successors 
    -- CP-element group 305: 	306 
    -- CP-element group 305: 	307 
    -- CP-element group 305:  members (10) 
      -- CP-element group 305: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475__exit__
      -- CP-element group 305: 	 branch_block_stmt_436/if_stmt_1476__entry__
      -- CP-element group 305: 	 branch_block_stmt_436/if_stmt_1476_eval_test/$exit
      -- CP-element group 305: 	 branch_block_stmt_436/if_stmt_1476_else_link/$entry
      -- CP-element group 305: 	 branch_block_stmt_436/if_stmt_1476_eval_test/$entry
      -- CP-element group 305: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/$exit
      -- CP-element group 305: 	 branch_block_stmt_436/if_stmt_1476_dead_link/$entry
      -- CP-element group 305: 	 branch_block_stmt_436/R_exitcond_1477_place
      -- CP-element group 305: 	 branch_block_stmt_436/if_stmt_1476_if_link/$entry
      -- CP-element group 305: 	 branch_block_stmt_436/if_stmt_1476_eval_test/branch_req
      -- 
    branch_req_3287_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3287_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(305), ack => if_stmt_1476_branch_req_0); -- 
    convolution3D_cp_element_group_305: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_305"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(243) & convolution3D_CP_1120_elements(299) & convolution3D_CP_1120_elements(304);
      gj_convolution3D_cp_element_group_305 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(305), clk => clk, reset => reset); --
    end block;
    -- CP-element group 306:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 306: predecessors 
    -- CP-element group 306: 	305 
    -- CP-element group 306: successors 
    -- CP-element group 306: 	400 
    -- CP-element group 306: 	401 
    -- CP-element group 306:  members (24) 
      -- CP-element group 306: 	 branch_block_stmt_436/merge_stmt_1482__exit__
      -- CP-element group 306: 	 branch_block_stmt_436/assign_stmt_1489_to_assign_stmt_1504__entry__
      -- CP-element group 306: 	 branch_block_stmt_436/assign_stmt_1489_to_assign_stmt_1504__exit__
      -- CP-element group 306: 	 branch_block_stmt_436/forx_xcond250x_xforx_xend341_crit_edge_forx_xend341
      -- CP-element group 306: 	 branch_block_stmt_436/assign_stmt_1489_to_assign_stmt_1504/$exit
      -- CP-element group 306: 	 branch_block_stmt_436/assign_stmt_1489_to_assign_stmt_1504/$entry
      -- CP-element group 306: 	 branch_block_stmt_436/if_stmt_1476_if_link/if_choice_transition
      -- CP-element group 306: 	 branch_block_stmt_436/if_stmt_1476_if_link/$exit
      -- CP-element group 306: 	 branch_block_stmt_436/forx_xbody257_forx_xcond250x_xforx_xend341_crit_edge
      -- CP-element group 306: 	 branch_block_stmt_436/forx_xbody257_forx_xcond250x_xforx_xend341_crit_edge_PhiReq/$entry
      -- CP-element group 306: 	 branch_block_stmt_436/forx_xbody257_forx_xcond250x_xforx_xend341_crit_edge_PhiReq/$exit
      -- CP-element group 306: 	 branch_block_stmt_436/merge_stmt_1482_PhiReqMerge
      -- CP-element group 306: 	 branch_block_stmt_436/merge_stmt_1482_PhiAck/$entry
      -- CP-element group 306: 	 branch_block_stmt_436/merge_stmt_1482_PhiAck/$exit
      -- CP-element group 306: 	 branch_block_stmt_436/merge_stmt_1482_PhiAck/dummy
      -- CP-element group 306: 	 branch_block_stmt_436/forx_xcond250x_xforx_xend341_crit_edge_forx_xend341_PhiReq/$entry
      -- CP-element group 306: 	 branch_block_stmt_436/forx_xcond250x_xforx_xend341_crit_edge_forx_xend341_PhiReq/phi_stmt_1507/$entry
      -- CP-element group 306: 	 branch_block_stmt_436/forx_xcond250x_xforx_xend341_crit_edge_forx_xend341_PhiReq/phi_stmt_1507/phi_stmt_1507_sources/$entry
      -- CP-element group 306: 	 branch_block_stmt_436/forx_xcond250x_xforx_xend341_crit_edge_forx_xend341_PhiReq/phi_stmt_1507/phi_stmt_1507_sources/type_cast_1510/$entry
      -- CP-element group 306: 	 branch_block_stmt_436/forx_xcond250x_xforx_xend341_crit_edge_forx_xend341_PhiReq/phi_stmt_1507/phi_stmt_1507_sources/type_cast_1510/SplitProtocol/$entry
      -- CP-element group 306: 	 branch_block_stmt_436/forx_xcond250x_xforx_xend341_crit_edge_forx_xend341_PhiReq/phi_stmt_1507/phi_stmt_1507_sources/type_cast_1510/SplitProtocol/Sample/$entry
      -- CP-element group 306: 	 branch_block_stmt_436/forx_xcond250x_xforx_xend341_crit_edge_forx_xend341_PhiReq/phi_stmt_1507/phi_stmt_1507_sources/type_cast_1510/SplitProtocol/Sample/rr
      -- CP-element group 306: 	 branch_block_stmt_436/forx_xcond250x_xforx_xend341_crit_edge_forx_xend341_PhiReq/phi_stmt_1507/phi_stmt_1507_sources/type_cast_1510/SplitProtocol/Update/$entry
      -- CP-element group 306: 	 branch_block_stmt_436/forx_xcond250x_xforx_xend341_crit_edge_forx_xend341_PhiReq/phi_stmt_1507/phi_stmt_1507_sources/type_cast_1510/SplitProtocol/Update/cr
      -- 
    if_choice_transition_3292_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 306_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1476_branch_ack_1, ack => convolution3D_CP_1120_elements(306)); -- 
    rr_4072_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4072_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(306), ack => type_cast_1510_inst_req_0); -- 
    cr_4077_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4077_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(306), ack => type_cast_1510_inst_req_1); -- 
    -- CP-element group 307:  fork  transition  place  input  output  bypass 
    -- CP-element group 307: predecessors 
    -- CP-element group 307: 	305 
    -- CP-element group 307: successors 
    -- CP-element group 307: 	395 
    -- CP-element group 307: 	396 
    -- CP-element group 307:  members (12) 
      -- CP-element group 307: 	 branch_block_stmt_436/if_stmt_1476_else_link/else_choice_transition
      -- CP-element group 307: 	 branch_block_stmt_436/if_stmt_1476_else_link/$exit
      -- CP-element group 307: 	 branch_block_stmt_436/forx_xbody257_forx_xbody257
      -- CP-element group 307: 	 branch_block_stmt_436/forx_xbody257_forx_xbody257_PhiReq/$entry
      -- CP-element group 307: 	 branch_block_stmt_436/forx_xbody257_forx_xbody257_PhiReq/phi_stmt_1289/$entry
      -- CP-element group 307: 	 branch_block_stmt_436/forx_xbody257_forx_xbody257_PhiReq/phi_stmt_1289/phi_stmt_1289_sources/$entry
      -- CP-element group 307: 	 branch_block_stmt_436/forx_xbody257_forx_xbody257_PhiReq/phi_stmt_1289/phi_stmt_1289_sources/type_cast_1295/$entry
      -- CP-element group 307: 	 branch_block_stmt_436/forx_xbody257_forx_xbody257_PhiReq/phi_stmt_1289/phi_stmt_1289_sources/type_cast_1295/SplitProtocol/$entry
      -- CP-element group 307: 	 branch_block_stmt_436/forx_xbody257_forx_xbody257_PhiReq/phi_stmt_1289/phi_stmt_1289_sources/type_cast_1295/SplitProtocol/Sample/$entry
      -- CP-element group 307: 	 branch_block_stmt_436/forx_xbody257_forx_xbody257_PhiReq/phi_stmt_1289/phi_stmt_1289_sources/type_cast_1295/SplitProtocol/Sample/rr
      -- CP-element group 307: 	 branch_block_stmt_436/forx_xbody257_forx_xbody257_PhiReq/phi_stmt_1289/phi_stmt_1289_sources/type_cast_1295/SplitProtocol/Update/$entry
      -- CP-element group 307: 	 branch_block_stmt_436/forx_xbody257_forx_xbody257_PhiReq/phi_stmt_1289/phi_stmt_1289_sources/type_cast_1295/SplitProtocol/Update/cr
      -- 
    else_choice_transition_3296_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 307_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1476_branch_ack_0, ack => convolution3D_CP_1120_elements(307)); -- 
    rr_4029_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4029_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(307), ack => type_cast_1295_inst_req_0); -- 
    cr_4034_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4034_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(307), ack => type_cast_1295_inst_req_1); -- 
    -- CP-element group 308:  transition  place  input  bypass 
    -- CP-element group 308: predecessors 
    -- CP-element group 308: 	405 
    -- CP-element group 308: successors 
    -- CP-element group 308: 	424 
    -- CP-element group 308:  members (5) 
      -- CP-element group 308: 	 branch_block_stmt_436/forx_xend341_ifx_xend353
      -- CP-element group 308: 	 branch_block_stmt_436/if_stmt_1527_if_link/if_choice_transition
      -- CP-element group 308: 	 branch_block_stmt_436/if_stmt_1527_if_link/$exit
      -- CP-element group 308: 	 branch_block_stmt_436/forx_xend341_ifx_xend353_PhiReq/$entry
      -- CP-element group 308: 	 branch_block_stmt_436/forx_xend341_ifx_xend353_PhiReq/$exit
      -- 
    if_choice_transition_3317_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 308_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1527_branch_ack_1, ack => convolution3D_CP_1120_elements(308)); -- 
    -- CP-element group 309:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 309: predecessors 
    -- CP-element group 309: 	405 
    -- CP-element group 309: successors 
    -- CP-element group 309: 	310 
    -- CP-element group 309: 	311 
    -- CP-element group 309:  members (18) 
      -- CP-element group 309: 	 branch_block_stmt_436/merge_stmt_1533__exit__
      -- CP-element group 309: 	 branch_block_stmt_436/assign_stmt_1539_to_assign_stmt_1549__entry__
      -- CP-element group 309: 	 branch_block_stmt_436/forx_xend341_bbx_xnphx_xi420
      -- CP-element group 309: 	 branch_block_stmt_436/assign_stmt_1539_to_assign_stmt_1549/type_cast_1542_Update/cr
      -- CP-element group 309: 	 branch_block_stmt_436/assign_stmt_1539_to_assign_stmt_1549/type_cast_1542_Update/$entry
      -- CP-element group 309: 	 branch_block_stmt_436/assign_stmt_1539_to_assign_stmt_1549/type_cast_1542_Sample/rr
      -- CP-element group 309: 	 branch_block_stmt_436/assign_stmt_1539_to_assign_stmt_1549/type_cast_1542_Sample/$entry
      -- CP-element group 309: 	 branch_block_stmt_436/assign_stmt_1539_to_assign_stmt_1549/type_cast_1542_update_start_
      -- CP-element group 309: 	 branch_block_stmt_436/assign_stmt_1539_to_assign_stmt_1549/type_cast_1542_sample_start_
      -- CP-element group 309: 	 branch_block_stmt_436/assign_stmt_1539_to_assign_stmt_1549/$entry
      -- CP-element group 309: 	 branch_block_stmt_436/if_stmt_1527_else_link/else_choice_transition
      -- CP-element group 309: 	 branch_block_stmt_436/if_stmt_1527_else_link/$exit
      -- CP-element group 309: 	 branch_block_stmt_436/forx_xend341_bbx_xnphx_xi420_PhiReq/$entry
      -- CP-element group 309: 	 branch_block_stmt_436/forx_xend341_bbx_xnphx_xi420_PhiReq/$exit
      -- CP-element group 309: 	 branch_block_stmt_436/merge_stmt_1533_PhiReqMerge
      -- CP-element group 309: 	 branch_block_stmt_436/merge_stmt_1533_PhiAck/$entry
      -- CP-element group 309: 	 branch_block_stmt_436/merge_stmt_1533_PhiAck/$exit
      -- CP-element group 309: 	 branch_block_stmt_436/merge_stmt_1533_PhiAck/dummy
      -- 
    else_choice_transition_3321_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 309_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1527_branch_ack_0, ack => convolution3D_CP_1120_elements(309)); -- 
    cr_3339_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3339_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(309), ack => type_cast_1542_inst_req_1); -- 
    rr_3334_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3334_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(309), ack => type_cast_1542_inst_req_0); -- 
    -- CP-element group 310:  transition  input  bypass 
    -- CP-element group 310: predecessors 
    -- CP-element group 310: 	309 
    -- CP-element group 310: successors 
    -- CP-element group 310:  members (3) 
      -- CP-element group 310: 	 branch_block_stmt_436/assign_stmt_1539_to_assign_stmt_1549/type_cast_1542_Sample/ra
      -- CP-element group 310: 	 branch_block_stmt_436/assign_stmt_1539_to_assign_stmt_1549/type_cast_1542_Sample/$exit
      -- CP-element group 310: 	 branch_block_stmt_436/assign_stmt_1539_to_assign_stmt_1549/type_cast_1542_sample_completed_
      -- 
    ra_3335_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 310_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1542_inst_ack_0, ack => convolution3D_CP_1120_elements(310)); -- 
    -- CP-element group 311:  fork  transition  place  input  bypass 
    -- CP-element group 311: predecessors 
    -- CP-element group 311: 	309 
    -- CP-element group 311: successors 
    -- CP-element group 311: 	406 
    -- CP-element group 311: 	407 
    -- CP-element group 311:  members (11) 
      -- CP-element group 311: 	 branch_block_stmt_436/assign_stmt_1539_to_assign_stmt_1549__exit__
      -- CP-element group 311: 	 branch_block_stmt_436/bbx_xnphx_xi420_forx_xbodyx_xi429
      -- CP-element group 311: 	 branch_block_stmt_436/assign_stmt_1539_to_assign_stmt_1549/type_cast_1542_Update/ca
      -- CP-element group 311: 	 branch_block_stmt_436/assign_stmt_1539_to_assign_stmt_1549/type_cast_1542_Update/$exit
      -- CP-element group 311: 	 branch_block_stmt_436/assign_stmt_1539_to_assign_stmt_1549/type_cast_1542_update_completed_
      -- CP-element group 311: 	 branch_block_stmt_436/assign_stmt_1539_to_assign_stmt_1549/$exit
      -- CP-element group 311: 	 branch_block_stmt_436/bbx_xnphx_xi420_forx_xbodyx_xi429_PhiReq/$entry
      -- CP-element group 311: 	 branch_block_stmt_436/bbx_xnphx_xi420_forx_xbodyx_xi429_PhiReq/phi_stmt_1552/$entry
      -- CP-element group 311: 	 branch_block_stmt_436/bbx_xnphx_xi420_forx_xbodyx_xi429_PhiReq/phi_stmt_1552/phi_stmt_1552_sources/$entry
      -- CP-element group 311: 	 branch_block_stmt_436/bbx_xnphx_xi420_forx_xbodyx_xi429_PhiReq/phi_stmt_1559/$entry
      -- CP-element group 311: 	 branch_block_stmt_436/bbx_xnphx_xi420_forx_xbodyx_xi429_PhiReq/phi_stmt_1559/phi_stmt_1559_sources/$entry
      -- 
    ca_3340_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 311_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1542_inst_ack_1, ack => convolution3D_CP_1120_elements(311)); -- 
    -- CP-element group 312:  transition  input  output  bypass 
    -- CP-element group 312: predecessors 
    -- CP-element group 312: 	419 
    -- CP-element group 312: successors 
    -- CP-element group 312: 	313 
    -- CP-element group 312:  members (6) 
      -- CP-element group 312: 	 branch_block_stmt_436/assign_stmt_1572_to_assign_stmt_1608/RPIPE_maxpool_input_pipe_1580_sample_completed_
      -- CP-element group 312: 	 branch_block_stmt_436/assign_stmt_1572_to_assign_stmt_1608/RPIPE_maxpool_input_pipe_1580_update_start_
      -- CP-element group 312: 	 branch_block_stmt_436/assign_stmt_1572_to_assign_stmt_1608/RPIPE_maxpool_input_pipe_1580_Sample/$exit
      -- CP-element group 312: 	 branch_block_stmt_436/assign_stmt_1572_to_assign_stmt_1608/RPIPE_maxpool_input_pipe_1580_Sample/ra
      -- CP-element group 312: 	 branch_block_stmt_436/assign_stmt_1572_to_assign_stmt_1608/RPIPE_maxpool_input_pipe_1580_Update/$entry
      -- CP-element group 312: 	 branch_block_stmt_436/assign_stmt_1572_to_assign_stmt_1608/RPIPE_maxpool_input_pipe_1580_Update/cr
      -- 
    ra_3352_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 312_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1580_inst_ack_0, ack => convolution3D_CP_1120_elements(312)); -- 
    cr_3356_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3356_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(312), ack => RPIPE_maxpool_input_pipe_1580_inst_req_1); -- 
    -- CP-element group 313:  fork  transition  input  output  bypass 
    -- CP-element group 313: predecessors 
    -- CP-element group 313: 	312 
    -- CP-element group 313: successors 
    -- CP-element group 313: 	314 
    -- CP-element group 313: 	316 
    -- CP-element group 313:  members (9) 
      -- CP-element group 313: 	 branch_block_stmt_436/assign_stmt_1572_to_assign_stmt_1608/RPIPE_maxpool_input_pipe_1580_update_completed_
      -- CP-element group 313: 	 branch_block_stmt_436/assign_stmt_1572_to_assign_stmt_1608/RPIPE_maxpool_input_pipe_1580_Update/$exit
      -- CP-element group 313: 	 branch_block_stmt_436/assign_stmt_1572_to_assign_stmt_1608/RPIPE_maxpool_input_pipe_1580_Update/ca
      -- CP-element group 313: 	 branch_block_stmt_436/assign_stmt_1572_to_assign_stmt_1608/WPIPE_maxpool_output_pipe_1582_sample_start_
      -- CP-element group 313: 	 branch_block_stmt_436/assign_stmt_1572_to_assign_stmt_1608/type_cast_1587_Sample/rr
      -- CP-element group 313: 	 branch_block_stmt_436/assign_stmt_1572_to_assign_stmt_1608/type_cast_1587_Sample/$entry
      -- CP-element group 313: 	 branch_block_stmt_436/assign_stmt_1572_to_assign_stmt_1608/type_cast_1587_sample_start_
      -- CP-element group 313: 	 branch_block_stmt_436/assign_stmt_1572_to_assign_stmt_1608/WPIPE_maxpool_output_pipe_1582_Sample/req
      -- CP-element group 313: 	 branch_block_stmt_436/assign_stmt_1572_to_assign_stmt_1608/WPIPE_maxpool_output_pipe_1582_Sample/$entry
      -- 
    ca_3357_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 313_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1580_inst_ack_1, ack => convolution3D_CP_1120_elements(313)); -- 
    req_3365_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3365_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(313), ack => WPIPE_maxpool_output_pipe_1582_inst_req_0); -- 
    rr_3379_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3379_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(313), ack => type_cast_1587_inst_req_0); -- 
    -- CP-element group 314:  transition  input  output  bypass 
    -- CP-element group 314: predecessors 
    -- CP-element group 314: 	313 
    -- CP-element group 314: successors 
    -- CP-element group 314: 	315 
    -- CP-element group 314:  members (6) 
      -- CP-element group 314: 	 branch_block_stmt_436/assign_stmt_1572_to_assign_stmt_1608/WPIPE_maxpool_output_pipe_1582_sample_completed_
      -- CP-element group 314: 	 branch_block_stmt_436/assign_stmt_1572_to_assign_stmt_1608/WPIPE_maxpool_output_pipe_1582_Update/req
      -- CP-element group 314: 	 branch_block_stmt_436/assign_stmt_1572_to_assign_stmt_1608/WPIPE_maxpool_output_pipe_1582_Update/$entry
      -- CP-element group 314: 	 branch_block_stmt_436/assign_stmt_1572_to_assign_stmt_1608/WPIPE_maxpool_output_pipe_1582_Sample/ack
      -- CP-element group 314: 	 branch_block_stmt_436/assign_stmt_1572_to_assign_stmt_1608/WPIPE_maxpool_output_pipe_1582_Sample/$exit
      -- CP-element group 314: 	 branch_block_stmt_436/assign_stmt_1572_to_assign_stmt_1608/WPIPE_maxpool_output_pipe_1582_update_start_
      -- 
    ack_3366_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 314_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1582_inst_ack_0, ack => convolution3D_CP_1120_elements(314)); -- 
    req_3370_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3370_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(314), ack => WPIPE_maxpool_output_pipe_1582_inst_req_1); -- 
    -- CP-element group 315:  transition  input  bypass 
    -- CP-element group 315: predecessors 
    -- CP-element group 315: 	314 
    -- CP-element group 315: successors 
    -- CP-element group 315: 	320 
    -- CP-element group 315:  members (3) 
      -- CP-element group 315: 	 branch_block_stmt_436/assign_stmt_1572_to_assign_stmt_1608/WPIPE_maxpool_output_pipe_1582_Update/ack
      -- CP-element group 315: 	 branch_block_stmt_436/assign_stmt_1572_to_assign_stmt_1608/WPIPE_maxpool_output_pipe_1582_Update/$exit
      -- CP-element group 315: 	 branch_block_stmt_436/assign_stmt_1572_to_assign_stmt_1608/WPIPE_maxpool_output_pipe_1582_update_completed_
      -- 
    ack_3371_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 315_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1582_inst_ack_1, ack => convolution3D_CP_1120_elements(315)); -- 
    -- CP-element group 316:  transition  input  bypass 
    -- CP-element group 316: predecessors 
    -- CP-element group 316: 	313 
    -- CP-element group 316: successors 
    -- CP-element group 316:  members (3) 
      -- CP-element group 316: 	 branch_block_stmt_436/assign_stmt_1572_to_assign_stmt_1608/type_cast_1587_Sample/ra
      -- CP-element group 316: 	 branch_block_stmt_436/assign_stmt_1572_to_assign_stmt_1608/type_cast_1587_Sample/$exit
      -- CP-element group 316: 	 branch_block_stmt_436/assign_stmt_1572_to_assign_stmt_1608/type_cast_1587_sample_completed_
      -- 
    ra_3380_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 316_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1587_inst_ack_0, ack => convolution3D_CP_1120_elements(316)); -- 
    -- CP-element group 317:  transition  input  bypass 
    -- CP-element group 317: predecessors 
    -- CP-element group 317: 	419 
    -- CP-element group 317: successors 
    -- CP-element group 317: 	320 
    -- CP-element group 317:  members (3) 
      -- CP-element group 317: 	 branch_block_stmt_436/assign_stmt_1572_to_assign_stmt_1608/type_cast_1587_Update/ca
      -- CP-element group 317: 	 branch_block_stmt_436/assign_stmt_1572_to_assign_stmt_1608/type_cast_1587_Update/$exit
      -- CP-element group 317: 	 branch_block_stmt_436/assign_stmt_1572_to_assign_stmt_1608/type_cast_1587_update_completed_
      -- 
    ca_3385_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 317_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1587_inst_ack_1, ack => convolution3D_CP_1120_elements(317)); -- 
    -- CP-element group 318:  transition  input  bypass 
    -- CP-element group 318: predecessors 
    -- CP-element group 318: 	419 
    -- CP-element group 318: successors 
    -- CP-element group 318:  members (3) 
      -- CP-element group 318: 	 branch_block_stmt_436/assign_stmt_1572_to_assign_stmt_1608/type_cast_1602_Sample/ra
      -- CP-element group 318: 	 branch_block_stmt_436/assign_stmt_1572_to_assign_stmt_1608/type_cast_1602_Sample/$exit
      -- CP-element group 318: 	 branch_block_stmt_436/assign_stmt_1572_to_assign_stmt_1608/type_cast_1602_sample_completed_
      -- 
    ra_3394_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 318_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1602_inst_ack_0, ack => convolution3D_CP_1120_elements(318)); -- 
    -- CP-element group 319:  transition  input  bypass 
    -- CP-element group 319: predecessors 
    -- CP-element group 319: 	419 
    -- CP-element group 319: successors 
    -- CP-element group 319: 	320 
    -- CP-element group 319:  members (3) 
      -- CP-element group 319: 	 branch_block_stmt_436/assign_stmt_1572_to_assign_stmt_1608/type_cast_1602_Update/ca
      -- CP-element group 319: 	 branch_block_stmt_436/assign_stmt_1572_to_assign_stmt_1608/type_cast_1602_Update/$exit
      -- CP-element group 319: 	 branch_block_stmt_436/assign_stmt_1572_to_assign_stmt_1608/type_cast_1602_update_completed_
      -- 
    ca_3399_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 319_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1602_inst_ack_1, ack => convolution3D_CP_1120_elements(319)); -- 
    -- CP-element group 320:  branch  join  transition  place  output  bypass 
    -- CP-element group 320: predecessors 
    -- CP-element group 320: 	315 
    -- CP-element group 320: 	317 
    -- CP-element group 320: 	319 
    -- CP-element group 320: successors 
    -- CP-element group 320: 	321 
    -- CP-element group 320: 	322 
    -- CP-element group 320:  members (10) 
      -- CP-element group 320: 	 branch_block_stmt_436/assign_stmt_1572_to_assign_stmt_1608__exit__
      -- CP-element group 320: 	 branch_block_stmt_436/if_stmt_1609__entry__
      -- CP-element group 320: 	 branch_block_stmt_436/R_cmpx_xi428_1610_place
      -- CP-element group 320: 	 branch_block_stmt_436/assign_stmt_1572_to_assign_stmt_1608/$exit
      -- CP-element group 320: 	 branch_block_stmt_436/if_stmt_1609_else_link/$entry
      -- CP-element group 320: 	 branch_block_stmt_436/if_stmt_1609_if_link/$entry
      -- CP-element group 320: 	 branch_block_stmt_436/if_stmt_1609_eval_test/branch_req
      -- CP-element group 320: 	 branch_block_stmt_436/if_stmt_1609_eval_test/$exit
      -- CP-element group 320: 	 branch_block_stmt_436/if_stmt_1609_eval_test/$entry
      -- CP-element group 320: 	 branch_block_stmt_436/if_stmt_1609_dead_link/$entry
      -- 
    branch_req_3407_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3407_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(320), ack => if_stmt_1609_branch_req_0); -- 
    convolution3D_cp_element_group_320: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_320"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(315) & convolution3D_CP_1120_elements(317) & convolution3D_CP_1120_elements(319);
      gj_convolution3D_cp_element_group_320 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(320), clk => clk, reset => reset); --
    end block;
    -- CP-element group 321:  fork  transition  place  input  output  bypass 
    -- CP-element group 321: predecessors 
    -- CP-element group 321: 	320 
    -- CP-element group 321: successors 
    -- CP-element group 321: 	410 
    -- CP-element group 321: 	412 
    -- CP-element group 321: 	413 
    -- CP-element group 321: 	409 
    -- CP-element group 321:  members (20) 
      -- CP-element group 321: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429
      -- CP-element group 321: 	 branch_block_stmt_436/if_stmt_1609_if_link/if_choice_transition
      -- CP-element group 321: 	 branch_block_stmt_436/if_stmt_1609_if_link/$exit
      -- CP-element group 321: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/$entry
      -- CP-element group 321: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1552/$entry
      -- CP-element group 321: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1552/phi_stmt_1552_sources/$entry
      -- CP-element group 321: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1552/phi_stmt_1552_sources/type_cast_1558/$entry
      -- CP-element group 321: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1552/phi_stmt_1552_sources/type_cast_1558/SplitProtocol/$entry
      -- CP-element group 321: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1552/phi_stmt_1552_sources/type_cast_1558/SplitProtocol/Sample/$entry
      -- CP-element group 321: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1552/phi_stmt_1552_sources/type_cast_1558/SplitProtocol/Sample/rr
      -- CP-element group 321: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1552/phi_stmt_1552_sources/type_cast_1558/SplitProtocol/Update/$entry
      -- CP-element group 321: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1552/phi_stmt_1552_sources/type_cast_1558/SplitProtocol/Update/cr
      -- CP-element group 321: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1559/$entry
      -- CP-element group 321: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1559/phi_stmt_1559_sources/$entry
      -- CP-element group 321: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1559/phi_stmt_1559_sources/type_cast_1565/$entry
      -- CP-element group 321: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1559/phi_stmt_1559_sources/type_cast_1565/SplitProtocol/$entry
      -- CP-element group 321: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1559/phi_stmt_1559_sources/type_cast_1565/SplitProtocol/Sample/$entry
      -- CP-element group 321: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1559/phi_stmt_1559_sources/type_cast_1565/SplitProtocol/Sample/rr
      -- CP-element group 321: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1559/phi_stmt_1559_sources/type_cast_1565/SplitProtocol/Update/$entry
      -- CP-element group 321: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1559/phi_stmt_1559_sources/type_cast_1565/SplitProtocol/Update/cr
      -- 
    if_choice_transition_3412_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 321_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1609_branch_ack_1, ack => convolution3D_CP_1120_elements(321)); -- 
    rr_4145_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4145_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(321), ack => type_cast_1558_inst_req_0); -- 
    cr_4150_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4150_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(321), ack => type_cast_1558_inst_req_1); -- 
    rr_4168_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4168_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(321), ack => type_cast_1565_inst_req_0); -- 
    cr_4173_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4173_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(321), ack => type_cast_1565_inst_req_1); -- 
    -- CP-element group 322:  fork  transition  place  input  output  bypass 
    -- CP-element group 322: predecessors 
    -- CP-element group 322: 	320 
    -- CP-element group 322: successors 
    -- CP-element group 322: 	420 
    -- CP-element group 322: 	421 
    -- CP-element group 322:  members (12) 
      -- CP-element group 322: 	 branch_block_stmt_436/forx_xbodyx_xi429_getRemainingElementsx_xexit437
      -- CP-element group 322: 	 branch_block_stmt_436/if_stmt_1609_else_link/else_choice_transition
      -- CP-element group 322: 	 branch_block_stmt_436/if_stmt_1609_else_link/$exit
      -- CP-element group 322: 	 branch_block_stmt_436/forx_xbodyx_xi429_getRemainingElementsx_xexit437_PhiReq/$entry
      -- CP-element group 322: 	 branch_block_stmt_436/forx_xbodyx_xi429_getRemainingElementsx_xexit437_PhiReq/phi_stmt_1616/$entry
      -- CP-element group 322: 	 branch_block_stmt_436/forx_xbodyx_xi429_getRemainingElementsx_xexit437_PhiReq/phi_stmt_1616/phi_stmt_1616_sources/$entry
      -- CP-element group 322: 	 branch_block_stmt_436/forx_xbodyx_xi429_getRemainingElementsx_xexit437_PhiReq/phi_stmt_1616/phi_stmt_1616_sources/type_cast_1619/$entry
      -- CP-element group 322: 	 branch_block_stmt_436/forx_xbodyx_xi429_getRemainingElementsx_xexit437_PhiReq/phi_stmt_1616/phi_stmt_1616_sources/type_cast_1619/SplitProtocol/$entry
      -- CP-element group 322: 	 branch_block_stmt_436/forx_xbodyx_xi429_getRemainingElementsx_xexit437_PhiReq/phi_stmt_1616/phi_stmt_1616_sources/type_cast_1619/SplitProtocol/Sample/$entry
      -- CP-element group 322: 	 branch_block_stmt_436/forx_xbodyx_xi429_getRemainingElementsx_xexit437_PhiReq/phi_stmt_1616/phi_stmt_1616_sources/type_cast_1619/SplitProtocol/Sample/rr
      -- CP-element group 322: 	 branch_block_stmt_436/forx_xbodyx_xi429_getRemainingElementsx_xexit437_PhiReq/phi_stmt_1616/phi_stmt_1616_sources/type_cast_1619/SplitProtocol/Update/$entry
      -- CP-element group 322: 	 branch_block_stmt_436/forx_xbodyx_xi429_getRemainingElementsx_xexit437_PhiReq/phi_stmt_1616/phi_stmt_1616_sources/type_cast_1619/SplitProtocol/Update/cr
      -- 
    else_choice_transition_3416_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 322_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1609_branch_ack_0, ack => convolution3D_CP_1120_elements(322)); -- 
    rr_4204_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4204_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(322), ack => type_cast_1619_inst_req_0); -- 
    cr_4209_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4209_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(322), ack => type_cast_1619_inst_req_1); -- 
    -- CP-element group 323:  transition  input  bypass 
    -- CP-element group 323: predecessors 
    -- CP-element group 323: 	423 
    -- CP-element group 323: successors 
    -- CP-element group 323: 	329 
    -- CP-element group 323:  members (3) 
      -- CP-element group 323: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/array_obj_ref_1648_final_index_sum_regn_Sample/ack
      -- CP-element group 323: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/array_obj_ref_1648_final_index_sum_regn_sample_complete
      -- CP-element group 323: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/array_obj_ref_1648_final_index_sum_regn_Sample/$exit
      -- 
    ack_3447_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 323_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1648_index_offset_ack_0, ack => convolution3D_CP_1120_elements(323)); -- 
    -- CP-element group 324:  transition  input  output  bypass 
    -- CP-element group 324: predecessors 
    -- CP-element group 324: 	423 
    -- CP-element group 324: successors 
    -- CP-element group 324: 	325 
    -- CP-element group 324:  members (11) 
      -- CP-element group 324: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/array_obj_ref_1648_offset_calculated
      -- CP-element group 324: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/array_obj_ref_1648_final_index_sum_regn_Update/$exit
      -- CP-element group 324: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/array_obj_ref_1648_root_address_calculated
      -- CP-element group 324: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/addr_of_1649_sample_start_
      -- CP-element group 324: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/addr_of_1649_request/req
      -- CP-element group 324: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/addr_of_1649_request/$entry
      -- CP-element group 324: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/array_obj_ref_1648_base_plus_offset/sum_rename_ack
      -- CP-element group 324: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/array_obj_ref_1648_base_plus_offset/sum_rename_req
      -- CP-element group 324: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/array_obj_ref_1648_base_plus_offset/$exit
      -- CP-element group 324: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/array_obj_ref_1648_base_plus_offset/$entry
      -- CP-element group 324: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/array_obj_ref_1648_final_index_sum_regn_Update/ack
      -- 
    ack_3452_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 324_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1648_index_offset_ack_1, ack => convolution3D_CP_1120_elements(324)); -- 
    req_3461_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3461_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(324), ack => addr_of_1649_final_reg_req_0); -- 
    -- CP-element group 325:  transition  input  bypass 
    -- CP-element group 325: predecessors 
    -- CP-element group 325: 	324 
    -- CP-element group 325: successors 
    -- CP-element group 325:  members (3) 
      -- CP-element group 325: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/addr_of_1649_sample_completed_
      -- CP-element group 325: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/addr_of_1649_request/ack
      -- CP-element group 325: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/addr_of_1649_request/$exit
      -- 
    ack_3462_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 325_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1649_final_reg_ack_0, ack => convolution3D_CP_1120_elements(325)); -- 
    -- CP-element group 326:  join  fork  transition  input  output  bypass 
    -- CP-element group 326: predecessors 
    -- CP-element group 326: 	423 
    -- CP-element group 326: successors 
    -- CP-element group 326: 	327 
    -- CP-element group 326:  members (28) 
      -- CP-element group 326: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/ptr_deref_1652_Sample/word_access_start/word_0/rr
      -- CP-element group 326: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/addr_of_1649_update_completed_
      -- CP-element group 326: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/ptr_deref_1652_Sample/word_access_start/word_0/$entry
      -- CP-element group 326: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/ptr_deref_1652_Sample/word_access_start/$entry
      -- CP-element group 326: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/ptr_deref_1652_Sample/ptr_deref_1652_Split/split_ack
      -- CP-element group 326: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/ptr_deref_1652_Sample/ptr_deref_1652_Split/split_req
      -- CP-element group 326: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/ptr_deref_1652_Sample/ptr_deref_1652_Split/$exit
      -- CP-element group 326: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/ptr_deref_1652_Sample/ptr_deref_1652_Split/$entry
      -- CP-element group 326: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/ptr_deref_1652_Sample/$entry
      -- CP-element group 326: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/ptr_deref_1652_word_addrgen/root_register_ack
      -- CP-element group 326: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/ptr_deref_1652_word_addrgen/root_register_req
      -- CP-element group 326: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/ptr_deref_1652_word_addrgen/$exit
      -- CP-element group 326: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/ptr_deref_1652_word_addrgen/$entry
      -- CP-element group 326: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/ptr_deref_1652_base_plus_offset/sum_rename_ack
      -- CP-element group 326: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/ptr_deref_1652_base_plus_offset/sum_rename_req
      -- CP-element group 326: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/ptr_deref_1652_base_plus_offset/$exit
      -- CP-element group 326: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/ptr_deref_1652_base_plus_offset/$entry
      -- CP-element group 326: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/ptr_deref_1652_base_addr_resize/base_resize_ack
      -- CP-element group 326: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/ptr_deref_1652_base_addr_resize/base_resize_req
      -- CP-element group 326: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/ptr_deref_1652_base_addr_resize/$exit
      -- CP-element group 326: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/ptr_deref_1652_base_addr_resize/$entry
      -- CP-element group 326: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/ptr_deref_1652_base_address_resized
      -- CP-element group 326: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/ptr_deref_1652_root_address_calculated
      -- CP-element group 326: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/ptr_deref_1652_word_address_calculated
      -- CP-element group 326: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/ptr_deref_1652_base_address_calculated
      -- CP-element group 326: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/ptr_deref_1652_sample_start_
      -- CP-element group 326: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/addr_of_1649_complete/ack
      -- CP-element group 326: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/addr_of_1649_complete/$exit
      -- 
    ack_3467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 326_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1649_final_reg_ack_1, ack => convolution3D_CP_1120_elements(326)); -- 
    rr_3505_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3505_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(326), ack => ptr_deref_1652_store_0_req_0); -- 
    -- CP-element group 327:  transition  input  bypass 
    -- CP-element group 327: predecessors 
    -- CP-element group 327: 	326 
    -- CP-element group 327: successors 
    -- CP-element group 327:  members (5) 
      -- CP-element group 327: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/ptr_deref_1652_Sample/word_access_start/word_0/ra
      -- CP-element group 327: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/ptr_deref_1652_Sample/word_access_start/word_0/$exit
      -- CP-element group 327: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/ptr_deref_1652_Sample/word_access_start/$exit
      -- CP-element group 327: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/ptr_deref_1652_Sample/$exit
      -- CP-element group 327: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/ptr_deref_1652_sample_completed_
      -- 
    ra_3506_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 327_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1652_store_0_ack_0, ack => convolution3D_CP_1120_elements(327)); -- 
    -- CP-element group 328:  transition  input  bypass 
    -- CP-element group 328: predecessors 
    -- CP-element group 328: 	423 
    -- CP-element group 328: successors 
    -- CP-element group 328: 	329 
    -- CP-element group 328:  members (5) 
      -- CP-element group 328: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/ptr_deref_1652_Update/$exit
      -- CP-element group 328: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/ptr_deref_1652_Update/word_access_complete/$exit
      -- CP-element group 328: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/ptr_deref_1652_update_completed_
      -- CP-element group 328: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/ptr_deref_1652_Update/word_access_complete/word_0/ca
      -- CP-element group 328: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/ptr_deref_1652_Update/word_access_complete/word_0/$exit
      -- 
    ca_3517_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 328_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1652_store_0_ack_1, ack => convolution3D_CP_1120_elements(328)); -- 
    -- CP-element group 329:  join  transition  place  bypass 
    -- CP-element group 329: predecessors 
    -- CP-element group 329: 	323 
    -- CP-element group 329: 	328 
    -- CP-element group 329: successors 
    -- CP-element group 329: 	424 
    -- CP-element group 329:  members (5) 
      -- CP-element group 329: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654__exit__
      -- CP-element group 329: 	 branch_block_stmt_436/getRemainingElementsx_xexit437_ifx_xend353
      -- CP-element group 329: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/$exit
      -- CP-element group 329: 	 branch_block_stmt_436/getRemainingElementsx_xexit437_ifx_xend353_PhiReq/$entry
      -- CP-element group 329: 	 branch_block_stmt_436/getRemainingElementsx_xexit437_ifx_xend353_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_329: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_329"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(323) & convolution3D_CP_1120_elements(328);
      gj_convolution3D_cp_element_group_329 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(329), clk => clk, reset => reset); --
    end block;
    -- CP-element group 330:  transition  input  bypass 
    -- CP-element group 330: predecessors 
    -- CP-element group 330: 	424 
    -- CP-element group 330: successors 
    -- CP-element group 330:  members (3) 
      -- CP-element group 330: 	 branch_block_stmt_436/call_stmt_1659/call_stmt_1659_Sample/cra
      -- CP-element group 330: 	 branch_block_stmt_436/call_stmt_1659/call_stmt_1659_Sample/$exit
      -- CP-element group 330: 	 branch_block_stmt_436/call_stmt_1659/call_stmt_1659_sample_completed_
      -- 
    cra_3529_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 330_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1659_call_ack_0, ack => convolution3D_CP_1120_elements(330)); -- 
    -- CP-element group 331:  fork  transition  place  input  output  bypass 
    -- CP-element group 331: predecessors 
    -- CP-element group 331: 	424 
    -- CP-element group 331: successors 
    -- CP-element group 331: 	332 
    -- CP-element group 331: 	334 
    -- CP-element group 331: 	336 
    -- CP-element group 331: 	337 
    -- CP-element group 331: 	338 
    -- CP-element group 331: 	339 
    -- CP-element group 331: 	340 
    -- CP-element group 331: 	341 
    -- CP-element group 331:  members (31) 
      -- CP-element group 331: 	 branch_block_stmt_436/assign_stmt_1665_to_assign_stmt_1723/WPIPE_num_out_pipe_1671_sample_start_
      -- CP-element group 331: 	 branch_block_stmt_436/call_stmt_1659__exit__
      -- CP-element group 331: 	 branch_block_stmt_436/assign_stmt_1665_to_assign_stmt_1723__entry__
      -- CP-element group 331: 	 branch_block_stmt_436/assign_stmt_1665_to_assign_stmt_1723/type_cast_1698_Sample/$entry
      -- CP-element group 331: 	 branch_block_stmt_436/assign_stmt_1665_to_assign_stmt_1723/type_cast_1698_Sample/rr
      -- CP-element group 331: 	 branch_block_stmt_436/assign_stmt_1665_to_assign_stmt_1723/type_cast_1708_update_start_
      -- CP-element group 331: 	 branch_block_stmt_436/assign_stmt_1665_to_assign_stmt_1723/type_cast_1698_Update/$entry
      -- CP-element group 331: 	 branch_block_stmt_436/assign_stmt_1665_to_assign_stmt_1723/type_cast_1698_Update/cr
      -- CP-element group 331: 	 branch_block_stmt_436/assign_stmt_1665_to_assign_stmt_1723/WPIPE_num_out_pipe_1671_Sample/$entry
      -- CP-element group 331: 	 branch_block_stmt_436/assign_stmt_1665_to_assign_stmt_1723/type_cast_1698_update_start_
      -- CP-element group 331: 	 branch_block_stmt_436/assign_stmt_1665_to_assign_stmt_1723/type_cast_1708_sample_start_
      -- CP-element group 331: 	 branch_block_stmt_436/assign_stmt_1665_to_assign_stmt_1723/$entry
      -- CP-element group 331: 	 branch_block_stmt_436/call_stmt_1659/call_stmt_1659_Update/cca
      -- CP-element group 331: 	 branch_block_stmt_436/assign_stmt_1665_to_assign_stmt_1723/type_cast_1717_Update/cr
      -- CP-element group 331: 	 branch_block_stmt_436/call_stmt_1659/call_stmt_1659_Update/$exit
      -- CP-element group 331: 	 branch_block_stmt_436/assign_stmt_1665_to_assign_stmt_1723/type_cast_1717_Update/$entry
      -- CP-element group 331: 	 branch_block_stmt_436/assign_stmt_1665_to_assign_stmt_1723/type_cast_1717_Sample/rr
      -- CP-element group 331: 	 branch_block_stmt_436/assign_stmt_1665_to_assign_stmt_1723/type_cast_1717_Sample/$entry
      -- CP-element group 331: 	 branch_block_stmt_436/call_stmt_1659/call_stmt_1659_update_completed_
      -- CP-element group 331: 	 branch_block_stmt_436/assign_stmt_1665_to_assign_stmt_1723/type_cast_1708_Sample/rr
      -- CP-element group 331: 	 branch_block_stmt_436/assign_stmt_1665_to_assign_stmt_1723/type_cast_1708_Sample/$entry
      -- CP-element group 331: 	 branch_block_stmt_436/assign_stmt_1665_to_assign_stmt_1723/type_cast_1717_update_start_
      -- CP-element group 331: 	 branch_block_stmt_436/assign_stmt_1665_to_assign_stmt_1723/type_cast_1698_sample_start_
      -- CP-element group 331: 	 branch_block_stmt_436/assign_stmt_1665_to_assign_stmt_1723/type_cast_1717_sample_start_
      -- CP-element group 331: 	 branch_block_stmt_436/call_stmt_1659/$exit
      -- CP-element group 331: 	 branch_block_stmt_436/assign_stmt_1665_to_assign_stmt_1723/WPIPE_maxpool_output_pipe_1674_Sample/req
      -- CP-element group 331: 	 branch_block_stmt_436/assign_stmt_1665_to_assign_stmt_1723/WPIPE_maxpool_output_pipe_1674_Sample/$entry
      -- CP-element group 331: 	 branch_block_stmt_436/assign_stmt_1665_to_assign_stmt_1723/type_cast_1708_Update/cr
      -- CP-element group 331: 	 branch_block_stmt_436/assign_stmt_1665_to_assign_stmt_1723/WPIPE_maxpool_output_pipe_1674_sample_start_
      -- CP-element group 331: 	 branch_block_stmt_436/assign_stmt_1665_to_assign_stmt_1723/type_cast_1708_Update/$entry
      -- CP-element group 331: 	 branch_block_stmt_436/assign_stmt_1665_to_assign_stmt_1723/WPIPE_num_out_pipe_1671_Sample/req
      -- 
    cca_3534_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 331_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1659_call_ack_1, ack => convolution3D_CP_1120_elements(331)); -- 
    rr_3573_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3573_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(331), ack => type_cast_1698_inst_req_0); -- 
    cr_3578_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3578_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(331), ack => type_cast_1698_inst_req_1); -- 
    cr_3606_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3606_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(331), ack => type_cast_1717_inst_req_1); -- 
    rr_3601_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3601_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(331), ack => type_cast_1717_inst_req_0); -- 
    rr_3587_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3587_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(331), ack => type_cast_1708_inst_req_0); -- 
    req_3559_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3559_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(331), ack => WPIPE_maxpool_output_pipe_1674_inst_req_0); -- 
    cr_3592_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3592_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(331), ack => type_cast_1708_inst_req_1); -- 
    req_3545_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3545_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(331), ack => WPIPE_num_out_pipe_1671_inst_req_0); -- 
    -- CP-element group 332:  transition  input  output  bypass 
    -- CP-element group 332: predecessors 
    -- CP-element group 332: 	331 
    -- CP-element group 332: successors 
    -- CP-element group 332: 	333 
    -- CP-element group 332:  members (6) 
      -- CP-element group 332: 	 branch_block_stmt_436/assign_stmt_1665_to_assign_stmt_1723/WPIPE_num_out_pipe_1671_sample_completed_
      -- CP-element group 332: 	 branch_block_stmt_436/assign_stmt_1665_to_assign_stmt_1723/WPIPE_num_out_pipe_1671_update_start_
      -- CP-element group 332: 	 branch_block_stmt_436/assign_stmt_1665_to_assign_stmt_1723/WPIPE_num_out_pipe_1671_Update/req
      -- CP-element group 332: 	 branch_block_stmt_436/assign_stmt_1665_to_assign_stmt_1723/WPIPE_num_out_pipe_1671_Update/$entry
      -- CP-element group 332: 	 branch_block_stmt_436/assign_stmt_1665_to_assign_stmt_1723/WPIPE_num_out_pipe_1671_Sample/ack
      -- CP-element group 332: 	 branch_block_stmt_436/assign_stmt_1665_to_assign_stmt_1723/WPIPE_num_out_pipe_1671_Sample/$exit
      -- 
    ack_3546_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 332_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_num_out_pipe_1671_inst_ack_0, ack => convolution3D_CP_1120_elements(332)); -- 
    req_3550_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3550_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(332), ack => WPIPE_num_out_pipe_1671_inst_req_1); -- 
    -- CP-element group 333:  transition  input  bypass 
    -- CP-element group 333: predecessors 
    -- CP-element group 333: 	332 
    -- CP-element group 333: successors 
    -- CP-element group 333: 	342 
    -- CP-element group 333:  members (3) 
      -- CP-element group 333: 	 branch_block_stmt_436/assign_stmt_1665_to_assign_stmt_1723/WPIPE_num_out_pipe_1671_update_completed_
      -- CP-element group 333: 	 branch_block_stmt_436/assign_stmt_1665_to_assign_stmt_1723/WPIPE_num_out_pipe_1671_Update/ack
      -- CP-element group 333: 	 branch_block_stmt_436/assign_stmt_1665_to_assign_stmt_1723/WPIPE_num_out_pipe_1671_Update/$exit
      -- 
    ack_3551_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 333_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_num_out_pipe_1671_inst_ack_1, ack => convolution3D_CP_1120_elements(333)); -- 
    -- CP-element group 334:  transition  input  output  bypass 
    -- CP-element group 334: predecessors 
    -- CP-element group 334: 	331 
    -- CP-element group 334: successors 
    -- CP-element group 334: 	335 
    -- CP-element group 334:  members (6) 
      -- CP-element group 334: 	 branch_block_stmt_436/assign_stmt_1665_to_assign_stmt_1723/WPIPE_maxpool_output_pipe_1674_Update/req
      -- CP-element group 334: 	 branch_block_stmt_436/assign_stmt_1665_to_assign_stmt_1723/WPIPE_maxpool_output_pipe_1674_Update/$entry
      -- CP-element group 334: 	 branch_block_stmt_436/assign_stmt_1665_to_assign_stmt_1723/WPIPE_maxpool_output_pipe_1674_Sample/ack
      -- CP-element group 334: 	 branch_block_stmt_436/assign_stmt_1665_to_assign_stmt_1723/WPIPE_maxpool_output_pipe_1674_Sample/$exit
      -- CP-element group 334: 	 branch_block_stmt_436/assign_stmt_1665_to_assign_stmt_1723/WPIPE_maxpool_output_pipe_1674_update_start_
      -- CP-element group 334: 	 branch_block_stmt_436/assign_stmt_1665_to_assign_stmt_1723/WPIPE_maxpool_output_pipe_1674_sample_completed_
      -- 
    ack_3560_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 334_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1674_inst_ack_0, ack => convolution3D_CP_1120_elements(334)); -- 
    req_3564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(334), ack => WPIPE_maxpool_output_pipe_1674_inst_req_1); -- 
    -- CP-element group 335:  transition  input  bypass 
    -- CP-element group 335: predecessors 
    -- CP-element group 335: 	334 
    -- CP-element group 335: successors 
    -- CP-element group 335: 	342 
    -- CP-element group 335:  members (3) 
      -- CP-element group 335: 	 branch_block_stmt_436/assign_stmt_1665_to_assign_stmt_1723/WPIPE_maxpool_output_pipe_1674_Update/ack
      -- CP-element group 335: 	 branch_block_stmt_436/assign_stmt_1665_to_assign_stmt_1723/WPIPE_maxpool_output_pipe_1674_Update/$exit
      -- CP-element group 335: 	 branch_block_stmt_436/assign_stmt_1665_to_assign_stmt_1723/WPIPE_maxpool_output_pipe_1674_update_completed_
      -- 
    ack_3565_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 335_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1674_inst_ack_1, ack => convolution3D_CP_1120_elements(335)); -- 
    -- CP-element group 336:  transition  input  bypass 
    -- CP-element group 336: predecessors 
    -- CP-element group 336: 	331 
    -- CP-element group 336: successors 
    -- CP-element group 336:  members (3) 
      -- CP-element group 336: 	 branch_block_stmt_436/assign_stmt_1665_to_assign_stmt_1723/type_cast_1698_Sample/$exit
      -- CP-element group 336: 	 branch_block_stmt_436/assign_stmt_1665_to_assign_stmt_1723/type_cast_1698_Sample/ra
      -- CP-element group 336: 	 branch_block_stmt_436/assign_stmt_1665_to_assign_stmt_1723/type_cast_1698_sample_completed_
      -- 
    ra_3574_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 336_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1698_inst_ack_0, ack => convolution3D_CP_1120_elements(336)); -- 
    -- CP-element group 337:  transition  input  bypass 
    -- CP-element group 337: predecessors 
    -- CP-element group 337: 	331 
    -- CP-element group 337: successors 
    -- CP-element group 337: 	342 
    -- CP-element group 337:  members (3) 
      -- CP-element group 337: 	 branch_block_stmt_436/assign_stmt_1665_to_assign_stmt_1723/type_cast_1698_update_completed_
      -- CP-element group 337: 	 branch_block_stmt_436/assign_stmt_1665_to_assign_stmt_1723/type_cast_1698_Update/$exit
      -- CP-element group 337: 	 branch_block_stmt_436/assign_stmt_1665_to_assign_stmt_1723/type_cast_1698_Update/ca
      -- 
    ca_3579_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 337_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1698_inst_ack_1, ack => convolution3D_CP_1120_elements(337)); -- 
    -- CP-element group 338:  transition  input  bypass 
    -- CP-element group 338: predecessors 
    -- CP-element group 338: 	331 
    -- CP-element group 338: successors 
    -- CP-element group 338:  members (3) 
      -- CP-element group 338: 	 branch_block_stmt_436/assign_stmt_1665_to_assign_stmt_1723/type_cast_1708_sample_completed_
      -- CP-element group 338: 	 branch_block_stmt_436/assign_stmt_1665_to_assign_stmt_1723/type_cast_1708_Sample/ra
      -- CP-element group 338: 	 branch_block_stmt_436/assign_stmt_1665_to_assign_stmt_1723/type_cast_1708_Sample/$exit
      -- 
    ra_3588_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 338_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1708_inst_ack_0, ack => convolution3D_CP_1120_elements(338)); -- 
    -- CP-element group 339:  transition  input  bypass 
    -- CP-element group 339: predecessors 
    -- CP-element group 339: 	331 
    -- CP-element group 339: successors 
    -- CP-element group 339: 	342 
    -- CP-element group 339:  members (3) 
      -- CP-element group 339: 	 branch_block_stmt_436/assign_stmt_1665_to_assign_stmt_1723/type_cast_1708_update_completed_
      -- CP-element group 339: 	 branch_block_stmt_436/assign_stmt_1665_to_assign_stmt_1723/type_cast_1708_Update/ca
      -- CP-element group 339: 	 branch_block_stmt_436/assign_stmt_1665_to_assign_stmt_1723/type_cast_1708_Update/$exit
      -- 
    ca_3593_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 339_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1708_inst_ack_1, ack => convolution3D_CP_1120_elements(339)); -- 
    -- CP-element group 340:  transition  input  bypass 
    -- CP-element group 340: predecessors 
    -- CP-element group 340: 	331 
    -- CP-element group 340: successors 
    -- CP-element group 340:  members (3) 
      -- CP-element group 340: 	 branch_block_stmt_436/assign_stmt_1665_to_assign_stmt_1723/type_cast_1717_Sample/ra
      -- CP-element group 340: 	 branch_block_stmt_436/assign_stmt_1665_to_assign_stmt_1723/type_cast_1717_Sample/$exit
      -- CP-element group 340: 	 branch_block_stmt_436/assign_stmt_1665_to_assign_stmt_1723/type_cast_1717_sample_completed_
      -- 
    ra_3602_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 340_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1717_inst_ack_0, ack => convolution3D_CP_1120_elements(340)); -- 
    -- CP-element group 341:  transition  input  bypass 
    -- CP-element group 341: predecessors 
    -- CP-element group 341: 	331 
    -- CP-element group 341: successors 
    -- CP-element group 341: 	342 
    -- CP-element group 341:  members (3) 
      -- CP-element group 341: 	 branch_block_stmt_436/assign_stmt_1665_to_assign_stmt_1723/type_cast_1717_Update/ca
      -- CP-element group 341: 	 branch_block_stmt_436/assign_stmt_1665_to_assign_stmt_1723/type_cast_1717_Update/$exit
      -- CP-element group 341: 	 branch_block_stmt_436/assign_stmt_1665_to_assign_stmt_1723/type_cast_1717_update_completed_
      -- 
    ca_3607_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 341_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1717_inst_ack_1, ack => convolution3D_CP_1120_elements(341)); -- 
    -- CP-element group 342:  join  transition  place  bypass 
    -- CP-element group 342: predecessors 
    -- CP-element group 342: 	333 
    -- CP-element group 342: 	335 
    -- CP-element group 342: 	337 
    -- CP-element group 342: 	339 
    -- CP-element group 342: 	341 
    -- CP-element group 342: successors 
    -- CP-element group 342: 	425 
    -- CP-element group 342:  members (6) 
      -- CP-element group 342: 	 branch_block_stmt_436/assign_stmt_1665_to_assign_stmt_1723__exit__
      -- CP-element group 342: 	 branch_block_stmt_436/ifx_xend353_whilex_xbody
      -- CP-element group 342: 	 branch_block_stmt_436/assign_stmt_1665_to_assign_stmt_1723/$exit
      -- CP-element group 342: 	 branch_block_stmt_436/ifx_xend353_whilex_xbody_PhiReq/$entry
      -- CP-element group 342: 	 branch_block_stmt_436/ifx_xend353_whilex_xbody_PhiReq/phi_stmt_1726/$entry
      -- CP-element group 342: 	 branch_block_stmt_436/ifx_xend353_whilex_xbody_PhiReq/phi_stmt_1726/phi_stmt_1726_sources/$entry
      -- 
    convolution3D_cp_element_group_342: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_342"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(333) & convolution3D_CP_1120_elements(335) & convolution3D_CP_1120_elements(337) & convolution3D_CP_1120_elements(339) & convolution3D_CP_1120_elements(341);
      gj_convolution3D_cp_element_group_342 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(342), clk => clk, reset => reset); --
    end block;
    -- CP-element group 343:  transition  input  bypass 
    -- CP-element group 343: predecessors 
    -- CP-element group 343: 	430 
    -- CP-element group 343: successors 
    -- CP-element group 343:  members (3) 
      -- CP-element group 343: 	 branch_block_stmt_436/assign_stmt_1738_to_assign_stmt_1772/type_cast_1746_Sample/$exit
      -- CP-element group 343: 	 branch_block_stmt_436/assign_stmt_1738_to_assign_stmt_1772/type_cast_1746_sample_completed_
      -- CP-element group 343: 	 branch_block_stmt_436/assign_stmt_1738_to_assign_stmt_1772/type_cast_1746_Sample/ra
      -- 
    ra_3619_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 343_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1746_inst_ack_0, ack => convolution3D_CP_1120_elements(343)); -- 
    -- CP-element group 344:  transition  input  bypass 
    -- CP-element group 344: predecessors 
    -- CP-element group 344: 	430 
    -- CP-element group 344: successors 
    -- CP-element group 344: 	347 
    -- CP-element group 344:  members (3) 
      -- CP-element group 344: 	 branch_block_stmt_436/assign_stmt_1738_to_assign_stmt_1772/type_cast_1746_update_completed_
      -- CP-element group 344: 	 branch_block_stmt_436/assign_stmt_1738_to_assign_stmt_1772/type_cast_1746_Update/ca
      -- CP-element group 344: 	 branch_block_stmt_436/assign_stmt_1738_to_assign_stmt_1772/type_cast_1746_Update/$exit
      -- 
    ca_3624_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 344_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1746_inst_ack_1, ack => convolution3D_CP_1120_elements(344)); -- 
    -- CP-element group 345:  transition  input  bypass 
    -- CP-element group 345: predecessors 
    -- CP-element group 345: 	430 
    -- CP-element group 345: successors 
    -- CP-element group 345:  members (3) 
      -- CP-element group 345: 	 branch_block_stmt_436/assign_stmt_1738_to_assign_stmt_1772/type_cast_1750_Sample/ra
      -- CP-element group 345: 	 branch_block_stmt_436/assign_stmt_1738_to_assign_stmt_1772/type_cast_1750_Sample/$exit
      -- CP-element group 345: 	 branch_block_stmt_436/assign_stmt_1738_to_assign_stmt_1772/type_cast_1750_sample_completed_
      -- 
    ra_3633_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 345_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1750_inst_ack_0, ack => convolution3D_CP_1120_elements(345)); -- 
    -- CP-element group 346:  transition  input  bypass 
    -- CP-element group 346: predecessors 
    -- CP-element group 346: 	430 
    -- CP-element group 346: successors 
    -- CP-element group 346: 	347 
    -- CP-element group 346:  members (3) 
      -- CP-element group 346: 	 branch_block_stmt_436/assign_stmt_1738_to_assign_stmt_1772/type_cast_1750_Update/ca
      -- CP-element group 346: 	 branch_block_stmt_436/assign_stmt_1738_to_assign_stmt_1772/type_cast_1750_Update/$exit
      -- CP-element group 346: 	 branch_block_stmt_436/assign_stmt_1738_to_assign_stmt_1772/type_cast_1750_update_completed_
      -- 
    ca_3638_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 346_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1750_inst_ack_1, ack => convolution3D_CP_1120_elements(346)); -- 
    -- CP-element group 347:  join  transition  output  bypass 
    -- CP-element group 347: predecessors 
    -- CP-element group 347: 	344 
    -- CP-element group 347: 	346 
    -- CP-element group 347: successors 
    -- CP-element group 347: 	348 
    -- CP-element group 347:  members (3) 
      -- CP-element group 347: 	 branch_block_stmt_436/assign_stmt_1738_to_assign_stmt_1772/call_stmt_1754_Sample/$entry
      -- CP-element group 347: 	 branch_block_stmt_436/assign_stmt_1738_to_assign_stmt_1772/call_stmt_1754_Sample/crr
      -- CP-element group 347: 	 branch_block_stmt_436/assign_stmt_1738_to_assign_stmt_1772/call_stmt_1754_sample_start_
      -- 
    crr_3646_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3646_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(347), ack => call_stmt_1754_call_req_0); -- 
    convolution3D_cp_element_group_347: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_347"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(344) & convolution3D_CP_1120_elements(346);
      gj_convolution3D_cp_element_group_347 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(347), clk => clk, reset => reset); --
    end block;
    -- CP-element group 348:  transition  input  bypass 
    -- CP-element group 348: predecessors 
    -- CP-element group 348: 	347 
    -- CP-element group 348: successors 
    -- CP-element group 348:  members (3) 
      -- CP-element group 348: 	 branch_block_stmt_436/assign_stmt_1738_to_assign_stmt_1772/call_stmt_1754_Sample/$exit
      -- CP-element group 348: 	 branch_block_stmt_436/assign_stmt_1738_to_assign_stmt_1772/call_stmt_1754_sample_completed_
      -- CP-element group 348: 	 branch_block_stmt_436/assign_stmt_1738_to_assign_stmt_1772/call_stmt_1754_Sample/cra
      -- 
    cra_3647_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 348_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1754_call_ack_0, ack => convolution3D_CP_1120_elements(348)); -- 
    -- CP-element group 349:  transition  input  bypass 
    -- CP-element group 349: predecessors 
    -- CP-element group 349: 	430 
    -- CP-element group 349: successors 
    -- CP-element group 349: 	352 
    -- CP-element group 349:  members (3) 
      -- CP-element group 349: 	 branch_block_stmt_436/assign_stmt_1738_to_assign_stmt_1772/call_stmt_1754_update_completed_
      -- CP-element group 349: 	 branch_block_stmt_436/assign_stmt_1738_to_assign_stmt_1772/call_stmt_1754_Update/$exit
      -- CP-element group 349: 	 branch_block_stmt_436/assign_stmt_1738_to_assign_stmt_1772/call_stmt_1754_Update/cca
      -- 
    cca_3652_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 349_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1754_call_ack_1, ack => convolution3D_CP_1120_elements(349)); -- 
    -- CP-element group 350:  transition  input  bypass 
    -- CP-element group 350: predecessors 
    -- CP-element group 350: 	430 
    -- CP-element group 350: successors 
    -- CP-element group 350:  members (3) 
      -- CP-element group 350: 	 branch_block_stmt_436/assign_stmt_1738_to_assign_stmt_1772/call_stmt_1761_Sample/cra
      -- CP-element group 350: 	 branch_block_stmt_436/assign_stmt_1738_to_assign_stmt_1772/call_stmt_1761_sample_completed_
      -- CP-element group 350: 	 branch_block_stmt_436/assign_stmt_1738_to_assign_stmt_1772/call_stmt_1761_Sample/$exit
      -- 
    cra_3661_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 350_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1761_call_ack_0, ack => convolution3D_CP_1120_elements(350)); -- 
    -- CP-element group 351:  transition  input  bypass 
    -- CP-element group 351: predecessors 
    -- CP-element group 351: 	430 
    -- CP-element group 351: successors 
    -- CP-element group 351: 	352 
    -- CP-element group 351:  members (3) 
      -- CP-element group 351: 	 branch_block_stmt_436/assign_stmt_1738_to_assign_stmt_1772/call_stmt_1761_Update/cca
      -- CP-element group 351: 	 branch_block_stmt_436/assign_stmt_1738_to_assign_stmt_1772/call_stmt_1761_update_completed_
      -- CP-element group 351: 	 branch_block_stmt_436/assign_stmt_1738_to_assign_stmt_1772/call_stmt_1761_Update/$exit
      -- 
    cca_3666_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 351_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1761_call_ack_1, ack => convolution3D_CP_1120_elements(351)); -- 
    -- CP-element group 352:  branch  join  transition  place  output  bypass 
    -- CP-element group 352: predecessors 
    -- CP-element group 352: 	349 
    -- CP-element group 352: 	351 
    -- CP-element group 352: successors 
    -- CP-element group 352: 	353 
    -- CP-element group 352: 	354 
    -- CP-element group 352:  members (10) 
      -- CP-element group 352: 	 branch_block_stmt_436/assign_stmt_1738_to_assign_stmt_1772__exit__
      -- CP-element group 352: 	 branch_block_stmt_436/if_stmt_1773__entry__
      -- CP-element group 352: 	 branch_block_stmt_436/R_exitcond5_1774_place
      -- CP-element group 352: 	 branch_block_stmt_436/if_stmt_1773_dead_link/$entry
      -- CP-element group 352: 	 branch_block_stmt_436/assign_stmt_1738_to_assign_stmt_1772/$exit
      -- CP-element group 352: 	 branch_block_stmt_436/if_stmt_1773_eval_test/$entry
      -- CP-element group 352: 	 branch_block_stmt_436/if_stmt_1773_eval_test/$exit
      -- CP-element group 352: 	 branch_block_stmt_436/if_stmt_1773_eval_test/branch_req
      -- CP-element group 352: 	 branch_block_stmt_436/if_stmt_1773_if_link/$entry
      -- CP-element group 352: 	 branch_block_stmt_436/if_stmt_1773_else_link/$entry
      -- 
    branch_req_3674_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3674_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(352), ack => if_stmt_1773_branch_req_0); -- 
    convolution3D_cp_element_group_352: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_352"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(349) & convolution3D_CP_1120_elements(351);
      gj_convolution3D_cp_element_group_352 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(352), clk => clk, reset => reset); --
    end block;
    -- CP-element group 353:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 353: predecessors 
    -- CP-element group 353: 	352 
    -- CP-element group 353: successors 
    -- CP-element group 353: 	355 
    -- CP-element group 353: 	356 
    -- CP-element group 353:  members (18) 
      -- CP-element group 353: 	 branch_block_stmt_436/merge_stmt_1779__exit__
      -- CP-element group 353: 	 branch_block_stmt_436/assign_stmt_1784__entry__
      -- CP-element group 353: 	 branch_block_stmt_436/whilex_xbody_whilex_xend
      -- CP-element group 353: 	 branch_block_stmt_436/if_stmt_1773_if_link/$exit
      -- CP-element group 353: 	 branch_block_stmt_436/if_stmt_1773_if_link/if_choice_transition
      -- CP-element group 353: 	 branch_block_stmt_436/assign_stmt_1784/$entry
      -- CP-element group 353: 	 branch_block_stmt_436/assign_stmt_1784/type_cast_1783_sample_start_
      -- CP-element group 353: 	 branch_block_stmt_436/assign_stmt_1784/type_cast_1783_update_start_
      -- CP-element group 353: 	 branch_block_stmt_436/assign_stmt_1784/type_cast_1783_Sample/$entry
      -- CP-element group 353: 	 branch_block_stmt_436/assign_stmt_1784/type_cast_1783_Sample/rr
      -- CP-element group 353: 	 branch_block_stmt_436/assign_stmt_1784/type_cast_1783_Update/$entry
      -- CP-element group 353: 	 branch_block_stmt_436/assign_stmt_1784/type_cast_1783_Update/cr
      -- CP-element group 353: 	 branch_block_stmt_436/whilex_xbody_whilex_xend_PhiReq/$entry
      -- CP-element group 353: 	 branch_block_stmt_436/whilex_xbody_whilex_xend_PhiReq/$exit
      -- CP-element group 353: 	 branch_block_stmt_436/merge_stmt_1779_PhiReqMerge
      -- CP-element group 353: 	 branch_block_stmt_436/merge_stmt_1779_PhiAck/$entry
      -- CP-element group 353: 	 branch_block_stmt_436/merge_stmt_1779_PhiAck/$exit
      -- CP-element group 353: 	 branch_block_stmt_436/merge_stmt_1779_PhiAck/dummy
      -- 
    if_choice_transition_3679_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 353_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1773_branch_ack_1, ack => convolution3D_CP_1120_elements(353)); -- 
    rr_3696_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3696_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(353), ack => type_cast_1783_inst_req_0); -- 
    cr_3701_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3701_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(353), ack => type_cast_1783_inst_req_1); -- 
    -- CP-element group 354:  fork  transition  place  input  output  bypass 
    -- CP-element group 354: predecessors 
    -- CP-element group 354: 	352 
    -- CP-element group 354: successors 
    -- CP-element group 354: 	426 
    -- CP-element group 354: 	427 
    -- CP-element group 354:  members (12) 
      -- CP-element group 354: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody
      -- CP-element group 354: 	 branch_block_stmt_436/if_stmt_1773_else_link/$exit
      -- CP-element group 354: 	 branch_block_stmt_436/if_stmt_1773_else_link/else_choice_transition
      -- CP-element group 354: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/$entry
      -- CP-element group 354: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1726/$entry
      -- CP-element group 354: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1726/phi_stmt_1726_sources/$entry
      -- CP-element group 354: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1726/phi_stmt_1726_sources/type_cast_1729/$entry
      -- CP-element group 354: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1726/phi_stmt_1726_sources/type_cast_1729/SplitProtocol/$entry
      -- CP-element group 354: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1726/phi_stmt_1726_sources/type_cast_1729/SplitProtocol/Sample/$entry
      -- CP-element group 354: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1726/phi_stmt_1726_sources/type_cast_1729/SplitProtocol/Sample/rr
      -- CP-element group 354: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1726/phi_stmt_1726_sources/type_cast_1729/SplitProtocol/Update/$entry
      -- CP-element group 354: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1726/phi_stmt_1726_sources/type_cast_1729/SplitProtocol/Update/cr
      -- 
    else_choice_transition_3683_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 354_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1773_branch_ack_0, ack => convolution3D_CP_1120_elements(354)); -- 
    rr_4257_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4257_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(354), ack => type_cast_1729_inst_req_0); -- 
    cr_4262_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4262_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(354), ack => type_cast_1729_inst_req_1); -- 
    -- CP-element group 355:  transition  input  bypass 
    -- CP-element group 355: predecessors 
    -- CP-element group 355: 	353 
    -- CP-element group 355: successors 
    -- CP-element group 355:  members (3) 
      -- CP-element group 355: 	 branch_block_stmt_436/assign_stmt_1784/type_cast_1783_sample_completed_
      -- CP-element group 355: 	 branch_block_stmt_436/assign_stmt_1784/type_cast_1783_Sample/$exit
      -- CP-element group 355: 	 branch_block_stmt_436/assign_stmt_1784/type_cast_1783_Sample/ra
      -- 
    ra_3697_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 355_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1783_inst_ack_0, ack => convolution3D_CP_1120_elements(355)); -- 
    -- CP-element group 356:  fork  transition  place  input  output  bypass 
    -- CP-element group 356: predecessors 
    -- CP-element group 356: 	353 
    -- CP-element group 356: successors 
    -- CP-element group 356: 	357 
    -- CP-element group 356: 	358 
    -- CP-element group 356: 	360 
    -- CP-element group 356:  members (16) 
      -- CP-element group 356: 	 branch_block_stmt_436/assign_stmt_1784__exit__
      -- CP-element group 356: 	 branch_block_stmt_436/call_stmt_1787_to_assign_stmt_1800__entry__
      -- CP-element group 356: 	 branch_block_stmt_436/assign_stmt_1784/$exit
      -- CP-element group 356: 	 branch_block_stmt_436/assign_stmt_1784/type_cast_1783_update_completed_
      -- CP-element group 356: 	 branch_block_stmt_436/assign_stmt_1784/type_cast_1783_Update/$exit
      -- CP-element group 356: 	 branch_block_stmt_436/assign_stmt_1784/type_cast_1783_Update/ca
      -- CP-element group 356: 	 branch_block_stmt_436/call_stmt_1787_to_assign_stmt_1800/$entry
      -- CP-element group 356: 	 branch_block_stmt_436/call_stmt_1787_to_assign_stmt_1800/call_stmt_1787_sample_start_
      -- CP-element group 356: 	 branch_block_stmt_436/call_stmt_1787_to_assign_stmt_1800/call_stmt_1787_update_start_
      -- CP-element group 356: 	 branch_block_stmt_436/call_stmt_1787_to_assign_stmt_1800/call_stmt_1787_Sample/$entry
      -- CP-element group 356: 	 branch_block_stmt_436/call_stmt_1787_to_assign_stmt_1800/call_stmt_1787_Sample/crr
      -- CP-element group 356: 	 branch_block_stmt_436/call_stmt_1787_to_assign_stmt_1800/call_stmt_1787_Update/$entry
      -- CP-element group 356: 	 branch_block_stmt_436/call_stmt_1787_to_assign_stmt_1800/call_stmt_1787_Update/ccr
      -- CP-element group 356: 	 branch_block_stmt_436/call_stmt_1787_to_assign_stmt_1800/type_cast_1791_update_start_
      -- CP-element group 356: 	 branch_block_stmt_436/call_stmt_1787_to_assign_stmt_1800/type_cast_1791_Update/$entry
      -- CP-element group 356: 	 branch_block_stmt_436/call_stmt_1787_to_assign_stmt_1800/type_cast_1791_Update/cr
      -- 
    ca_3702_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 356_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1783_inst_ack_1, ack => convolution3D_CP_1120_elements(356)); -- 
    crr_3713_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3713_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(356), ack => call_stmt_1787_call_req_0); -- 
    ccr_3718_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3718_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(356), ack => call_stmt_1787_call_req_1); -- 
    cr_3732_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3732_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(356), ack => type_cast_1791_inst_req_1); -- 
    -- CP-element group 357:  transition  input  bypass 
    -- CP-element group 357: predecessors 
    -- CP-element group 357: 	356 
    -- CP-element group 357: successors 
    -- CP-element group 357:  members (3) 
      -- CP-element group 357: 	 branch_block_stmt_436/call_stmt_1787_to_assign_stmt_1800/call_stmt_1787_sample_completed_
      -- CP-element group 357: 	 branch_block_stmt_436/call_stmt_1787_to_assign_stmt_1800/call_stmt_1787_Sample/$exit
      -- CP-element group 357: 	 branch_block_stmt_436/call_stmt_1787_to_assign_stmt_1800/call_stmt_1787_Sample/cra
      -- 
    cra_3714_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 357_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1787_call_ack_0, ack => convolution3D_CP_1120_elements(357)); -- 
    -- CP-element group 358:  transition  input  output  bypass 
    -- CP-element group 358: predecessors 
    -- CP-element group 358: 	356 
    -- CP-element group 358: successors 
    -- CP-element group 358: 	359 
    -- CP-element group 358:  members (6) 
      -- CP-element group 358: 	 branch_block_stmt_436/call_stmt_1787_to_assign_stmt_1800/call_stmt_1787_update_completed_
      -- CP-element group 358: 	 branch_block_stmt_436/call_stmt_1787_to_assign_stmt_1800/call_stmt_1787_Update/$exit
      -- CP-element group 358: 	 branch_block_stmt_436/call_stmt_1787_to_assign_stmt_1800/call_stmt_1787_Update/cca
      -- CP-element group 358: 	 branch_block_stmt_436/call_stmt_1787_to_assign_stmt_1800/type_cast_1791_sample_start_
      -- CP-element group 358: 	 branch_block_stmt_436/call_stmt_1787_to_assign_stmt_1800/type_cast_1791_Sample/$entry
      -- CP-element group 358: 	 branch_block_stmt_436/call_stmt_1787_to_assign_stmt_1800/type_cast_1791_Sample/rr
      -- 
    cca_3719_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 358_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1787_call_ack_1, ack => convolution3D_CP_1120_elements(358)); -- 
    rr_3727_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3727_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(358), ack => type_cast_1791_inst_req_0); -- 
    -- CP-element group 359:  transition  input  bypass 
    -- CP-element group 359: predecessors 
    -- CP-element group 359: 	358 
    -- CP-element group 359: successors 
    -- CP-element group 359:  members (3) 
      -- CP-element group 359: 	 branch_block_stmt_436/call_stmt_1787_to_assign_stmt_1800/type_cast_1791_sample_completed_
      -- CP-element group 359: 	 branch_block_stmt_436/call_stmt_1787_to_assign_stmt_1800/type_cast_1791_Sample/$exit
      -- CP-element group 359: 	 branch_block_stmt_436/call_stmt_1787_to_assign_stmt_1800/type_cast_1791_Sample/ra
      -- 
    ra_3728_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 359_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1791_inst_ack_0, ack => convolution3D_CP_1120_elements(359)); -- 
    -- CP-element group 360:  transition  input  output  bypass 
    -- CP-element group 360: predecessors 
    -- CP-element group 360: 	356 
    -- CP-element group 360: successors 
    -- CP-element group 360: 	361 
    -- CP-element group 360:  members (6) 
      -- CP-element group 360: 	 branch_block_stmt_436/call_stmt_1787_to_assign_stmt_1800/type_cast_1791_update_completed_
      -- CP-element group 360: 	 branch_block_stmt_436/call_stmt_1787_to_assign_stmt_1800/type_cast_1791_Update/$exit
      -- CP-element group 360: 	 branch_block_stmt_436/call_stmt_1787_to_assign_stmt_1800/type_cast_1791_Update/ca
      -- CP-element group 360: 	 branch_block_stmt_436/call_stmt_1787_to_assign_stmt_1800/WPIPE_elapsed_time_pipe_1798_sample_start_
      -- CP-element group 360: 	 branch_block_stmt_436/call_stmt_1787_to_assign_stmt_1800/WPIPE_elapsed_time_pipe_1798_Sample/$entry
      -- CP-element group 360: 	 branch_block_stmt_436/call_stmt_1787_to_assign_stmt_1800/WPIPE_elapsed_time_pipe_1798_Sample/req
      -- 
    ca_3733_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 360_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1791_inst_ack_1, ack => convolution3D_CP_1120_elements(360)); -- 
    req_3741_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3741_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(360), ack => WPIPE_elapsed_time_pipe_1798_inst_req_0); -- 
    -- CP-element group 361:  transition  input  output  bypass 
    -- CP-element group 361: predecessors 
    -- CP-element group 361: 	360 
    -- CP-element group 361: successors 
    -- CP-element group 361: 	362 
    -- CP-element group 361:  members (6) 
      -- CP-element group 361: 	 branch_block_stmt_436/call_stmt_1787_to_assign_stmt_1800/WPIPE_elapsed_time_pipe_1798_sample_completed_
      -- CP-element group 361: 	 branch_block_stmt_436/call_stmt_1787_to_assign_stmt_1800/WPIPE_elapsed_time_pipe_1798_update_start_
      -- CP-element group 361: 	 branch_block_stmt_436/call_stmt_1787_to_assign_stmt_1800/WPIPE_elapsed_time_pipe_1798_Sample/$exit
      -- CP-element group 361: 	 branch_block_stmt_436/call_stmt_1787_to_assign_stmt_1800/WPIPE_elapsed_time_pipe_1798_Sample/ack
      -- CP-element group 361: 	 branch_block_stmt_436/call_stmt_1787_to_assign_stmt_1800/WPIPE_elapsed_time_pipe_1798_Update/$entry
      -- CP-element group 361: 	 branch_block_stmt_436/call_stmt_1787_to_assign_stmt_1800/WPIPE_elapsed_time_pipe_1798_Update/req
      -- 
    ack_3742_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 361_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_elapsed_time_pipe_1798_inst_ack_0, ack => convolution3D_CP_1120_elements(361)); -- 
    req_3746_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3746_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(361), ack => WPIPE_elapsed_time_pipe_1798_inst_req_1); -- 
    -- CP-element group 362:  transition  place  input  bypass 
    -- CP-element group 362: predecessors 
    -- CP-element group 362: 	361 
    -- CP-element group 362: successors 
    -- CP-element group 362:  members (16) 
      -- CP-element group 362: 	 $exit
      -- CP-element group 362: 	 branch_block_stmt_436/$exit
      -- CP-element group 362: 	 branch_block_stmt_436/branch_block_stmt_436__exit__
      -- CP-element group 362: 	 branch_block_stmt_436/call_stmt_1787_to_assign_stmt_1800__exit__
      -- CP-element group 362: 	 branch_block_stmt_436/return__
      -- CP-element group 362: 	 branch_block_stmt_436/merge_stmt_1803__exit__
      -- CP-element group 362: 	 branch_block_stmt_436/merge_stmt_1803_PhiReqMerge
      -- CP-element group 362: 	 branch_block_stmt_436/call_stmt_1787_to_assign_stmt_1800/$exit
      -- CP-element group 362: 	 branch_block_stmt_436/call_stmt_1787_to_assign_stmt_1800/WPIPE_elapsed_time_pipe_1798_update_completed_
      -- CP-element group 362: 	 branch_block_stmt_436/call_stmt_1787_to_assign_stmt_1800/WPIPE_elapsed_time_pipe_1798_Update/$exit
      -- CP-element group 362: 	 branch_block_stmt_436/call_stmt_1787_to_assign_stmt_1800/WPIPE_elapsed_time_pipe_1798_Update/ack
      -- CP-element group 362: 	 branch_block_stmt_436/return___PhiReq/$entry
      -- CP-element group 362: 	 branch_block_stmt_436/return___PhiReq/$exit
      -- CP-element group 362: 	 branch_block_stmt_436/merge_stmt_1803_PhiAck/$entry
      -- CP-element group 362: 	 branch_block_stmt_436/merge_stmt_1803_PhiAck/$exit
      -- CP-element group 362: 	 branch_block_stmt_436/merge_stmt_1803_PhiAck/dummy
      -- 
    ack_3747_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 362_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_elapsed_time_pipe_1798_inst_ack_1, ack => convolution3D_CP_1120_elements(362)); -- 
    -- CP-element group 363:  transition  output  delay-element  bypass 
    -- CP-element group 363: predecessors 
    -- CP-element group 363: 	133 
    -- CP-element group 363: successors 
    -- CP-element group 363: 	367 
    -- CP-element group 363:  members (5) 
      -- CP-element group 363: 	 branch_block_stmt_436/bbx_xnph449_forx_xbody_PhiReq/$exit
      -- CP-element group 363: 	 branch_block_stmt_436/bbx_xnph449_forx_xbody_PhiReq/phi_stmt_793/$exit
      -- CP-element group 363: 	 branch_block_stmt_436/bbx_xnph449_forx_xbody_PhiReq/phi_stmt_793/phi_stmt_793_sources/$exit
      -- CP-element group 363: 	 branch_block_stmt_436/bbx_xnph449_forx_xbody_PhiReq/phi_stmt_793/phi_stmt_793_sources/type_cast_797_konst_delay_trans
      -- CP-element group 363: 	 branch_block_stmt_436/bbx_xnph449_forx_xbody_PhiReq/phi_stmt_793/phi_stmt_793_req
      -- 
    phi_stmt_793_req_3770_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_793_req_3770_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(363), ack => phi_stmt_793_req_0); -- 
    -- Element group convolution3D_CP_1120_elements(363) is a control-delay.
    cp_element_363_delay: control_delay_element  generic map(name => " 363_delay", delay_value => 1)  port map(req => convolution3D_CP_1120_elements(133), ack => convolution3D_CP_1120_elements(363), clk => clk, reset =>reset);
    -- CP-element group 364:  transition  input  bypass 
    -- CP-element group 364: predecessors 
    -- CP-element group 364: 	198 
    -- CP-element group 364: successors 
    -- CP-element group 364: 	366 
    -- CP-element group 364:  members (2) 
      -- CP-element group 364: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_793/phi_stmt_793_sources/type_cast_799/SplitProtocol/Sample/$exit
      -- CP-element group 364: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_793/phi_stmt_793_sources/type_cast_799/SplitProtocol/Sample/ra
      -- 
    ra_3790_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 364_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_799_inst_ack_0, ack => convolution3D_CP_1120_elements(364)); -- 
    -- CP-element group 365:  transition  input  bypass 
    -- CP-element group 365: predecessors 
    -- CP-element group 365: 	198 
    -- CP-element group 365: successors 
    -- CP-element group 365: 	366 
    -- CP-element group 365:  members (2) 
      -- CP-element group 365: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_793/phi_stmt_793_sources/type_cast_799/SplitProtocol/Update/$exit
      -- CP-element group 365: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_793/phi_stmt_793_sources/type_cast_799/SplitProtocol/Update/ca
      -- 
    ca_3795_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 365_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_799_inst_ack_1, ack => convolution3D_CP_1120_elements(365)); -- 
    -- CP-element group 366:  join  transition  output  bypass 
    -- CP-element group 366: predecessors 
    -- CP-element group 366: 	364 
    -- CP-element group 366: 	365 
    -- CP-element group 366: successors 
    -- CP-element group 366: 	367 
    -- CP-element group 366:  members (6) 
      -- CP-element group 366: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 366: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_793/$exit
      -- CP-element group 366: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_793/phi_stmt_793_sources/$exit
      -- CP-element group 366: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_793/phi_stmt_793_sources/type_cast_799/$exit
      -- CP-element group 366: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_793/phi_stmt_793_sources/type_cast_799/SplitProtocol/$exit
      -- CP-element group 366: 	 branch_block_stmt_436/forx_xbody_forx_xbody_PhiReq/phi_stmt_793/phi_stmt_793_req
      -- 
    phi_stmt_793_req_3796_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_793_req_3796_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(366), ack => phi_stmt_793_req_1); -- 
    convolution3D_cp_element_group_366: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_366"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(364) & convolution3D_CP_1120_elements(365);
      gj_convolution3D_cp_element_group_366 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(366), clk => clk, reset => reset); --
    end block;
    -- CP-element group 367:  merge  transition  place  bypass 
    -- CP-element group 367: predecessors 
    -- CP-element group 367: 	363 
    -- CP-element group 367: 	366 
    -- CP-element group 367: successors 
    -- CP-element group 367: 	368 
    -- CP-element group 367:  members (2) 
      -- CP-element group 367: 	 branch_block_stmt_436/merge_stmt_792_PhiReqMerge
      -- CP-element group 367: 	 branch_block_stmt_436/merge_stmt_792_PhiAck/$entry
      -- 
    convolution3D_CP_1120_elements(367) <= OrReduce(convolution3D_CP_1120_elements(363) & convolution3D_CP_1120_elements(366));
    -- CP-element group 368:  fork  transition  place  input  output  bypass 
    -- CP-element group 368: predecessors 
    -- CP-element group 368: 	367 
    -- CP-element group 368: successors 
    -- CP-element group 368: 	134 
    -- CP-element group 368: 	135 
    -- CP-element group 368: 	137 
    -- CP-element group 368: 	138 
    -- CP-element group 368: 	143 
    -- CP-element group 368: 	150 
    -- CP-element group 368: 	157 
    -- CP-element group 368: 	164 
    -- CP-element group 368: 	171 
    -- CP-element group 368: 	178 
    -- CP-element group 368: 	185 
    -- CP-element group 368: 	192 
    -- CP-element group 368: 	195 
    -- CP-element group 368:  members (56) 
      -- CP-element group 368: 	 branch_block_stmt_436/merge_stmt_792__exit__
      -- CP-element group 368: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979__entry__
      -- CP-element group 368: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/ptr_deref_966_Update/$entry
      -- CP-element group 368: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/ptr_deref_966_Update/word_access_complete/$entry
      -- CP-element group 368: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_937_Update/cr
      -- CP-element group 368: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/ptr_deref_966_Update/word_access_complete/word_0/cr
      -- CP-element group 368: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/ptr_deref_966_Update/word_access_complete/word_0/$entry
      -- CP-element group 368: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_937_Update/$entry
      -- CP-element group 368: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/ptr_deref_966_update_start_
      -- CP-element group 368: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_958_Update/cr
      -- CP-element group 368: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_958_Update/$entry
      -- CP-element group 368: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_937_update_start_
      -- CP-element group 368: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/$entry
      -- CP-element group 368: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/addr_of_806_update_start_
      -- CP-element group 368: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/array_obj_ref_805_index_resized_1
      -- CP-element group 368: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_958_update_start_
      -- CP-element group 368: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/array_obj_ref_805_index_scaled_1
      -- CP-element group 368: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/array_obj_ref_805_index_computed_1
      -- CP-element group 368: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/array_obj_ref_805_index_resize_1/$entry
      -- CP-element group 368: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/array_obj_ref_805_index_resize_1/$exit
      -- CP-element group 368: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/array_obj_ref_805_index_resize_1/index_resize_req
      -- CP-element group 368: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/array_obj_ref_805_index_resize_1/index_resize_ack
      -- CP-element group 368: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/array_obj_ref_805_index_scale_1/$entry
      -- CP-element group 368: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/array_obj_ref_805_index_scale_1/$exit
      -- CP-element group 368: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/array_obj_ref_805_index_scale_1/scale_rename_req
      -- CP-element group 368: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/array_obj_ref_805_index_scale_1/scale_rename_ack
      -- CP-element group 368: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/array_obj_ref_805_final_index_sum_regn_update_start
      -- CP-element group 368: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/array_obj_ref_805_final_index_sum_regn_Sample/$entry
      -- CP-element group 368: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/array_obj_ref_805_final_index_sum_regn_Sample/req
      -- CP-element group 368: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/array_obj_ref_805_final_index_sum_regn_Update/$entry
      -- CP-element group 368: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/array_obj_ref_805_final_index_sum_regn_Update/req
      -- CP-element group 368: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/addr_of_806_complete/$entry
      -- CP-element group 368: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/addr_of_806_complete/req
      -- CP-element group 368: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_809_sample_start_
      -- CP-element group 368: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_809_Sample/$entry
      -- CP-element group 368: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/RPIPE_maxpool_input_pipe_809_Sample/rr
      -- CP-element group 368: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_816_update_start_
      -- CP-element group 368: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_816_Update/$entry
      -- CP-element group 368: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_816_Update/cr
      -- CP-element group 368: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_832_update_start_
      -- CP-element group 368: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_832_Update/$entry
      -- CP-element group 368: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_832_Update/cr
      -- CP-element group 368: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_853_update_start_
      -- CP-element group 368: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_853_Update/$entry
      -- CP-element group 368: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_853_Update/cr
      -- CP-element group 368: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_874_update_start_
      -- CP-element group 368: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_874_Update/$entry
      -- CP-element group 368: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_874_Update/cr
      -- CP-element group 368: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_895_update_start_
      -- CP-element group 368: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_895_Update/$entry
      -- CP-element group 368: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_895_Update/cr
      -- CP-element group 368: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_916_update_start_
      -- CP-element group 368: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_916_Update/$entry
      -- CP-element group 368: 	 branch_block_stmt_436/assign_stmt_807_to_assign_stmt_979/type_cast_916_Update/cr
      -- CP-element group 368: 	 branch_block_stmt_436/merge_stmt_792_PhiAck/$exit
      -- CP-element group 368: 	 branch_block_stmt_436/merge_stmt_792_PhiAck/phi_stmt_793_ack
      -- 
    phi_stmt_793_ack_3801_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 368_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_793_ack_0, ack => convolution3D_CP_1120_elements(368)); -- 
    cr_2362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(368), ack => type_cast_937_inst_req_1); -- 
    cr_2454_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2454_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(368), ack => ptr_deref_966_store_0_req_1); -- 
    cr_2404_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2404_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(368), ack => type_cast_958_inst_req_1); -- 
    req_2048_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2048_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(368), ack => array_obj_ref_805_index_offset_req_0); -- 
    req_2053_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2053_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(368), ack => array_obj_ref_805_index_offset_req_1); -- 
    req_2068_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2068_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(368), ack => addr_of_806_final_reg_req_1); -- 
    rr_2077_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2077_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(368), ack => RPIPE_maxpool_input_pipe_809_inst_req_0); -- 
    cr_2110_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2110_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(368), ack => type_cast_816_inst_req_1); -- 
    cr_2152_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2152_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(368), ack => type_cast_832_inst_req_1); -- 
    cr_2194_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2194_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(368), ack => type_cast_853_inst_req_1); -- 
    cr_2236_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2236_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(368), ack => type_cast_874_inst_req_1); -- 
    cr_2278_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2278_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(368), ack => type_cast_895_inst_req_1); -- 
    cr_2320_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2320_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(368), ack => type_cast_916_inst_req_1); -- 
    -- CP-element group 369:  transition  output  delay-element  bypass 
    -- CP-element group 369: predecessors 
    -- CP-element group 369: 	123 
    -- CP-element group 369: successors 
    -- CP-element group 369: 	373 
    -- CP-element group 369:  members (5) 
      -- CP-element group 369: 	 branch_block_stmt_436/entry_forx_xend_PhiReq/$exit
      -- CP-element group 369: 	 branch_block_stmt_436/entry_forx_xend_PhiReq/phi_stmt_1011/$exit
      -- CP-element group 369: 	 branch_block_stmt_436/entry_forx_xend_PhiReq/phi_stmt_1011/phi_stmt_1011_sources/$exit
      -- CP-element group 369: 	 branch_block_stmt_436/entry_forx_xend_PhiReq/phi_stmt_1011/phi_stmt_1011_sources/type_cast_1017_konst_delay_trans
      -- CP-element group 369: 	 branch_block_stmt_436/entry_forx_xend_PhiReq/phi_stmt_1011/phi_stmt_1011_req
      -- 
    phi_stmt_1011_req_3824_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1011_req_3824_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(369), ack => phi_stmt_1011_req_1); -- 
    -- Element group convolution3D_CP_1120_elements(369) is a control-delay.
    cp_element_369_delay: control_delay_element  generic map(name => " 369_delay", delay_value => 1)  port map(req => convolution3D_CP_1120_elements(123), ack => convolution3D_CP_1120_elements(369), clk => clk, reset =>reset);
    -- CP-element group 370:  transition  input  bypass 
    -- CP-element group 370: predecessors 
    -- CP-element group 370: 	197 
    -- CP-element group 370: successors 
    -- CP-element group 370: 	372 
    -- CP-element group 370:  members (2) 
      -- CP-element group 370: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1011/phi_stmt_1011_sources/type_cast_1014/SplitProtocol/Sample/$exit
      -- CP-element group 370: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1011/phi_stmt_1011_sources/type_cast_1014/SplitProtocol/Sample/ra
      -- 
    ra_3844_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 370_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1014_inst_ack_0, ack => convolution3D_CP_1120_elements(370)); -- 
    -- CP-element group 371:  transition  input  bypass 
    -- CP-element group 371: predecessors 
    -- CP-element group 371: 	197 
    -- CP-element group 371: successors 
    -- CP-element group 371: 	372 
    -- CP-element group 371:  members (2) 
      -- CP-element group 371: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1011/phi_stmt_1011_sources/type_cast_1014/SplitProtocol/Update/$exit
      -- CP-element group 371: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1011/phi_stmt_1011_sources/type_cast_1014/SplitProtocol/Update/ca
      -- 
    ca_3849_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 371_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1014_inst_ack_1, ack => convolution3D_CP_1120_elements(371)); -- 
    -- CP-element group 372:  join  transition  output  bypass 
    -- CP-element group 372: predecessors 
    -- CP-element group 372: 	370 
    -- CP-element group 372: 	371 
    -- CP-element group 372: successors 
    -- CP-element group 372: 	373 
    -- CP-element group 372:  members (6) 
      -- CP-element group 372: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/$exit
      -- CP-element group 372: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1011/$exit
      -- CP-element group 372: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1011/phi_stmt_1011_sources/$exit
      -- CP-element group 372: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1011/phi_stmt_1011_sources/type_cast_1014/$exit
      -- CP-element group 372: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1011/phi_stmt_1011_sources/type_cast_1014/SplitProtocol/$exit
      -- CP-element group 372: 	 branch_block_stmt_436/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_1011/phi_stmt_1011_req
      -- 
    phi_stmt_1011_req_3850_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1011_req_3850_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(372), ack => phi_stmt_1011_req_0); -- 
    convolution3D_cp_element_group_372: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_372"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(370) & convolution3D_CP_1120_elements(371);
      gj_convolution3D_cp_element_group_372 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(372), clk => clk, reset => reset); --
    end block;
    -- CP-element group 373:  merge  transition  place  bypass 
    -- CP-element group 373: predecessors 
    -- CP-element group 373: 	369 
    -- CP-element group 373: 	372 
    -- CP-element group 373: successors 
    -- CP-element group 373: 	374 
    -- CP-element group 373:  members (2) 
      -- CP-element group 373: 	 branch_block_stmt_436/merge_stmt_1010_PhiReqMerge
      -- CP-element group 373: 	 branch_block_stmt_436/merge_stmt_1010_PhiAck/$entry
      -- 
    convolution3D_CP_1120_elements(373) <= OrReduce(convolution3D_CP_1120_elements(369) & convolution3D_CP_1120_elements(372));
    -- CP-element group 374:  branch  transition  place  input  output  bypass 
    -- CP-element group 374: predecessors 
    -- CP-element group 374: 	373 
    -- CP-element group 374: successors 
    -- CP-element group 374: 	199 
    -- CP-element group 374: 	200 
    -- CP-element group 374:  members (15) 
      -- CP-element group 374: 	 branch_block_stmt_436/merge_stmt_1010__exit__
      -- CP-element group 374: 	 branch_block_stmt_436/assign_stmt_1024_to_assign_stmt_1030__entry__
      -- CP-element group 374: 	 branch_block_stmt_436/assign_stmt_1024_to_assign_stmt_1030__exit__
      -- CP-element group 374: 	 branch_block_stmt_436/if_stmt_1031__entry__
      -- CP-element group 374: 	 branch_block_stmt_436/if_stmt_1031_else_link/$entry
      -- CP-element group 374: 	 branch_block_stmt_436/if_stmt_1031_if_link/$entry
      -- CP-element group 374: 	 branch_block_stmt_436/if_stmt_1031_eval_test/branch_req
      -- CP-element group 374: 	 branch_block_stmt_436/if_stmt_1031_eval_test/$exit
      -- CP-element group 374: 	 branch_block_stmt_436/R_tobool_1032_place
      -- CP-element group 374: 	 branch_block_stmt_436/if_stmt_1031_eval_test/$entry
      -- CP-element group 374: 	 branch_block_stmt_436/if_stmt_1031_dead_link/$entry
      -- CP-element group 374: 	 branch_block_stmt_436/assign_stmt_1024_to_assign_stmt_1030/$exit
      -- CP-element group 374: 	 branch_block_stmt_436/assign_stmt_1024_to_assign_stmt_1030/$entry
      -- CP-element group 374: 	 branch_block_stmt_436/merge_stmt_1010_PhiAck/$exit
      -- CP-element group 374: 	 branch_block_stmt_436/merge_stmt_1010_PhiAck/phi_stmt_1011_ack
      -- 
    phi_stmt_1011_ack_3855_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 374_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1011_ack_0, ack => convolution3D_CP_1120_elements(374)); -- 
    branch_req_2488_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2488_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(374), ack => if_stmt_1031_branch_req_0); -- 
    -- CP-element group 375:  transition  output  delay-element  bypass 
    -- CP-element group 375: predecessors 
    -- CP-element group 375: 	200 
    -- CP-element group 375: successors 
    -- CP-element group 375: 	377 
    -- CP-element group 375:  members (4) 
      -- CP-element group 375: 	 branch_block_stmt_436/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1052/$exit
      -- CP-element group 375: 	 branch_block_stmt_436/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1052/phi_stmt_1052_sources/$exit
      -- CP-element group 375: 	 branch_block_stmt_436/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1052/phi_stmt_1052_sources/type_cast_1056_konst_delay_trans
      -- CP-element group 375: 	 branch_block_stmt_436/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1052/phi_stmt_1052_req
      -- 
    phi_stmt_1052_req_3878_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1052_req_3878_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(375), ack => phi_stmt_1052_req_0); -- 
    -- Element group convolution3D_CP_1120_elements(375) is a control-delay.
    cp_element_375_delay: control_delay_element  generic map(name => " 375_delay", delay_value => 1)  port map(req => convolution3D_CP_1120_elements(200), ack => convolution3D_CP_1120_elements(375), clk => clk, reset =>reset);
    -- CP-element group 376:  transition  output  delay-element  bypass 
    -- CP-element group 376: predecessors 
    -- CP-element group 376: 	200 
    -- CP-element group 376: successors 
    -- CP-element group 376: 	377 
    -- CP-element group 376:  members (4) 
      -- CP-element group 376: 	 branch_block_stmt_436/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1059/$exit
      -- CP-element group 376: 	 branch_block_stmt_436/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1059/phi_stmt_1059_sources/$exit
      -- CP-element group 376: 	 branch_block_stmt_436/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1059/phi_stmt_1059_sources/type_cast_1063_konst_delay_trans
      -- CP-element group 376: 	 branch_block_stmt_436/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1059/phi_stmt_1059_req
      -- 
    phi_stmt_1059_req_3886_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1059_req_3886_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(376), ack => phi_stmt_1059_req_0); -- 
    -- Element group convolution3D_CP_1120_elements(376) is a control-delay.
    cp_element_376_delay: control_delay_element  generic map(name => " 376_delay", delay_value => 1)  port map(req => convolution3D_CP_1120_elements(200), ack => convolution3D_CP_1120_elements(376), clk => clk, reset =>reset);
    -- CP-element group 377:  join  transition  bypass 
    -- CP-element group 377: predecessors 
    -- CP-element group 377: 	375 
    -- CP-element group 377: 	376 
    -- CP-element group 377: successors 
    -- CP-element group 377: 	385 
    -- CP-element group 377:  members (1) 
      -- CP-element group 377: 	 branch_block_stmt_436/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_377: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_377"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(375) & convolution3D_CP_1120_elements(376);
      gj_convolution3D_cp_element_group_377 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(377), clk => clk, reset => reset); --
    end block;
    -- CP-element group 378:  transition  input  bypass 
    -- CP-element group 378: predecessors 
    -- CP-element group 378: 	210 
    -- CP-element group 378: successors 
    -- CP-element group 378: 	380 
    -- CP-element group 378:  members (2) 
      -- CP-element group 378: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1052/phi_stmt_1052_sources/type_cast_1058/SplitProtocol/Sample/$exit
      -- CP-element group 378: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1052/phi_stmt_1052_sources/type_cast_1058/SplitProtocol/Sample/ra
      -- 
    ra_3906_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 378_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1058_inst_ack_0, ack => convolution3D_CP_1120_elements(378)); -- 
    -- CP-element group 379:  transition  input  bypass 
    -- CP-element group 379: predecessors 
    -- CP-element group 379: 	210 
    -- CP-element group 379: successors 
    -- CP-element group 379: 	380 
    -- CP-element group 379:  members (2) 
      -- CP-element group 379: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1052/phi_stmt_1052_sources/type_cast_1058/SplitProtocol/Update/$exit
      -- CP-element group 379: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1052/phi_stmt_1052_sources/type_cast_1058/SplitProtocol/Update/ca
      -- 
    ca_3911_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 379_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1058_inst_ack_1, ack => convolution3D_CP_1120_elements(379)); -- 
    -- CP-element group 380:  join  transition  output  bypass 
    -- CP-element group 380: predecessors 
    -- CP-element group 380: 	378 
    -- CP-element group 380: 	379 
    -- CP-element group 380: successors 
    -- CP-element group 380: 	384 
    -- CP-element group 380:  members (5) 
      -- CP-element group 380: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1052/$exit
      -- CP-element group 380: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1052/phi_stmt_1052_sources/$exit
      -- CP-element group 380: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1052/phi_stmt_1052_sources/type_cast_1058/$exit
      -- CP-element group 380: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1052/phi_stmt_1052_sources/type_cast_1058/SplitProtocol/$exit
      -- CP-element group 380: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1052/phi_stmt_1052_req
      -- 
    phi_stmt_1052_req_3912_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1052_req_3912_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(380), ack => phi_stmt_1052_req_1); -- 
    convolution3D_cp_element_group_380: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_380"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(378) & convolution3D_CP_1120_elements(379);
      gj_convolution3D_cp_element_group_380 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(380), clk => clk, reset => reset); --
    end block;
    -- CP-element group 381:  transition  input  bypass 
    -- CP-element group 381: predecessors 
    -- CP-element group 381: 	210 
    -- CP-element group 381: successors 
    -- CP-element group 381: 	383 
    -- CP-element group 381:  members (2) 
      -- CP-element group 381: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1059/phi_stmt_1059_sources/type_cast_1065/SplitProtocol/Sample/$exit
      -- CP-element group 381: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1059/phi_stmt_1059_sources/type_cast_1065/SplitProtocol/Sample/ra
      -- 
    ra_3929_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 381_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1065_inst_ack_0, ack => convolution3D_CP_1120_elements(381)); -- 
    -- CP-element group 382:  transition  input  bypass 
    -- CP-element group 382: predecessors 
    -- CP-element group 382: 	210 
    -- CP-element group 382: successors 
    -- CP-element group 382: 	383 
    -- CP-element group 382:  members (2) 
      -- CP-element group 382: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1059/phi_stmt_1059_sources/type_cast_1065/SplitProtocol/Update/$exit
      -- CP-element group 382: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1059/phi_stmt_1059_sources/type_cast_1065/SplitProtocol/Update/ca
      -- 
    ca_3934_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 382_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1065_inst_ack_1, ack => convolution3D_CP_1120_elements(382)); -- 
    -- CP-element group 383:  join  transition  output  bypass 
    -- CP-element group 383: predecessors 
    -- CP-element group 383: 	381 
    -- CP-element group 383: 	382 
    -- CP-element group 383: successors 
    -- CP-element group 383: 	384 
    -- CP-element group 383:  members (5) 
      -- CP-element group 383: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1059/$exit
      -- CP-element group 383: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1059/phi_stmt_1059_sources/$exit
      -- CP-element group 383: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1059/phi_stmt_1059_sources/type_cast_1065/$exit
      -- CP-element group 383: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1059/phi_stmt_1059_sources/type_cast_1065/SplitProtocol/$exit
      -- CP-element group 383: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1059/phi_stmt_1059_req
      -- 
    phi_stmt_1059_req_3935_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1059_req_3935_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(383), ack => phi_stmt_1059_req_1); -- 
    convolution3D_cp_element_group_383: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_383"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(381) & convolution3D_CP_1120_elements(382);
      gj_convolution3D_cp_element_group_383 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(383), clk => clk, reset => reset); --
    end block;
    -- CP-element group 384:  join  transition  bypass 
    -- CP-element group 384: predecessors 
    -- CP-element group 384: 	380 
    -- CP-element group 384: 	383 
    -- CP-element group 384: successors 
    -- CP-element group 384: 	385 
    -- CP-element group 384:  members (1) 
      -- CP-element group 384: 	 branch_block_stmt_436/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_384: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_384"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(380) & convolution3D_CP_1120_elements(383);
      gj_convolution3D_cp_element_group_384 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(384), clk => clk, reset => reset); --
    end block;
    -- CP-element group 385:  merge  fork  transition  place  bypass 
    -- CP-element group 385: predecessors 
    -- CP-element group 385: 	377 
    -- CP-element group 385: 	384 
    -- CP-element group 385: successors 
    -- CP-element group 385: 	386 
    -- CP-element group 385: 	387 
    -- CP-element group 385:  members (2) 
      -- CP-element group 385: 	 branch_block_stmt_436/merge_stmt_1051_PhiReqMerge
      -- CP-element group 385: 	 branch_block_stmt_436/merge_stmt_1051_PhiAck/$entry
      -- 
    convolution3D_CP_1120_elements(385) <= OrReduce(convolution3D_CP_1120_elements(377) & convolution3D_CP_1120_elements(384));
    -- CP-element group 386:  transition  input  bypass 
    -- CP-element group 386: predecessors 
    -- CP-element group 386: 	385 
    -- CP-element group 386: successors 
    -- CP-element group 386: 	388 
    -- CP-element group 386:  members (1) 
      -- CP-element group 386: 	 branch_block_stmt_436/merge_stmt_1051_PhiAck/phi_stmt_1052_ack
      -- 
    phi_stmt_1052_ack_3940_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 386_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1052_ack_0, ack => convolution3D_CP_1120_elements(386)); -- 
    -- CP-element group 387:  transition  input  bypass 
    -- CP-element group 387: predecessors 
    -- CP-element group 387: 	385 
    -- CP-element group 387: successors 
    -- CP-element group 387: 	388 
    -- CP-element group 387:  members (1) 
      -- CP-element group 387: 	 branch_block_stmt_436/merge_stmt_1051_PhiAck/phi_stmt_1059_ack
      -- 
    phi_stmt_1059_ack_3941_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 387_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1059_ack_0, ack => convolution3D_CP_1120_elements(387)); -- 
    -- CP-element group 388:  join  fork  transition  place  output  bypass 
    -- CP-element group 388: predecessors 
    -- CP-element group 388: 	386 
    -- CP-element group 388: 	387 
    -- CP-element group 388: successors 
    -- CP-element group 388: 	201 
    -- CP-element group 388: 	206 
    -- CP-element group 388: 	207 
    -- CP-element group 388: 	208 
    -- CP-element group 388:  members (16) 
      -- CP-element group 388: 	 branch_block_stmt_436/assign_stmt_1072_to_assign_stmt_1108/type_cast_1102_Update/$entry
      -- CP-element group 388: 	 branch_block_stmt_436/assign_stmt_1072_to_assign_stmt_1108/type_cast_1102_Update/cr
      -- CP-element group 388: 	 branch_block_stmt_436/merge_stmt_1051__exit__
      -- CP-element group 388: 	 branch_block_stmt_436/assign_stmt_1072_to_assign_stmt_1108__entry__
      -- CP-element group 388: 	 branch_block_stmt_436/assign_stmt_1072_to_assign_stmt_1108/type_cast_1102_Sample/rr
      -- CP-element group 388: 	 branch_block_stmt_436/assign_stmt_1072_to_assign_stmt_1108/RPIPE_maxpool_input_pipe_1080_Sample/rr
      -- CP-element group 388: 	 branch_block_stmt_436/assign_stmt_1072_to_assign_stmt_1108/RPIPE_maxpool_input_pipe_1080_Sample/$entry
      -- CP-element group 388: 	 branch_block_stmt_436/assign_stmt_1072_to_assign_stmt_1108/type_cast_1102_Sample/$entry
      -- CP-element group 388: 	 branch_block_stmt_436/assign_stmt_1072_to_assign_stmt_1108/type_cast_1102_update_start_
      -- CP-element group 388: 	 branch_block_stmt_436/assign_stmt_1072_to_assign_stmt_1108/RPIPE_maxpool_input_pipe_1080_sample_start_
      -- CP-element group 388: 	 branch_block_stmt_436/assign_stmt_1072_to_assign_stmt_1108/$entry
      -- CP-element group 388: 	 branch_block_stmt_436/assign_stmt_1072_to_assign_stmt_1108/type_cast_1102_sample_start_
      -- CP-element group 388: 	 branch_block_stmt_436/assign_stmt_1072_to_assign_stmt_1108/type_cast_1087_Update/cr
      -- CP-element group 388: 	 branch_block_stmt_436/assign_stmt_1072_to_assign_stmt_1108/type_cast_1087_Update/$entry
      -- CP-element group 388: 	 branch_block_stmt_436/assign_stmt_1072_to_assign_stmt_1108/type_cast_1087_update_start_
      -- CP-element group 388: 	 branch_block_stmt_436/merge_stmt_1051_PhiAck/$exit
      -- 
    cr_2560_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2560_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(388), ack => type_cast_1102_inst_req_1); -- 
    rr_2555_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2555_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(388), ack => type_cast_1102_inst_req_0); -- 
    rr_2513_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2513_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(388), ack => RPIPE_maxpool_input_pipe_1080_inst_req_0); -- 
    cr_2546_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2546_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(388), ack => type_cast_1087_inst_req_1); -- 
    convolution3D_cp_element_group_388: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_388"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(386) & convolution3D_CP_1120_elements(387);
      gj_convolution3D_cp_element_group_388 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(388), clk => clk, reset => reset); --
    end block;
    -- CP-element group 389:  transition  input  bypass 
    -- CP-element group 389: predecessors 
    -- CP-element group 389: 	211 
    -- CP-element group 389: successors 
    -- CP-element group 389: 	391 
    -- CP-element group 389:  members (2) 
      -- CP-element group 389: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1116/phi_stmt_1116_sources/type_cast_1119/SplitProtocol/Sample/$exit
      -- CP-element group 389: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1116/phi_stmt_1116_sources/type_cast_1119/SplitProtocol/Sample/ra
      -- 
    ra_3965_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 389_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1119_inst_ack_0, ack => convolution3D_CP_1120_elements(389)); -- 
    -- CP-element group 390:  transition  input  bypass 
    -- CP-element group 390: predecessors 
    -- CP-element group 390: 	211 
    -- CP-element group 390: successors 
    -- CP-element group 390: 	391 
    -- CP-element group 390:  members (2) 
      -- CP-element group 390: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1116/phi_stmt_1116_sources/type_cast_1119/SplitProtocol/Update/$exit
      -- CP-element group 390: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1116/phi_stmt_1116_sources/type_cast_1119/SplitProtocol/Update/ca
      -- 
    ca_3970_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 390_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1119_inst_ack_1, ack => convolution3D_CP_1120_elements(390)); -- 
    -- CP-element group 391:  join  transition  place  output  bypass 
    -- CP-element group 391: predecessors 
    -- CP-element group 391: 	389 
    -- CP-element group 391: 	390 
    -- CP-element group 391: successors 
    -- CP-element group 391: 	392 
    -- CP-element group 391:  members (8) 
      -- CP-element group 391: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/$exit
      -- CP-element group 391: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1116/$exit
      -- CP-element group 391: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1116/phi_stmt_1116_sources/$exit
      -- CP-element group 391: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1116/phi_stmt_1116_sources/type_cast_1119/$exit
      -- CP-element group 391: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1116/phi_stmt_1116_sources/type_cast_1119/SplitProtocol/$exit
      -- CP-element group 391: 	 branch_block_stmt_436/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1116/phi_stmt_1116_req
      -- CP-element group 391: 	 branch_block_stmt_436/merge_stmt_1115_PhiReqMerge
      -- CP-element group 391: 	 branch_block_stmt_436/merge_stmt_1115_PhiAck/$entry
      -- 
    phi_stmt_1116_req_3971_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1116_req_3971_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(391), ack => phi_stmt_1116_req_0); -- 
    convolution3D_cp_element_group_391: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_391"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(389) & convolution3D_CP_1120_elements(390);
      gj_convolution3D_cp_element_group_391 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(391), clk => clk, reset => reset); --
    end block;
    -- CP-element group 392:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 392: predecessors 
    -- CP-element group 392: 	391 
    -- CP-element group 392: successors 
    -- CP-element group 392: 	212 
    -- CP-element group 392: 	213 
    -- CP-element group 392: 	215 
    -- CP-element group 392: 	217 
    -- CP-element group 392:  members (29) 
      -- CP-element group 392: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/array_obj_ref_1148_index_resize_1/index_resize_ack
      -- CP-element group 392: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/array_obj_ref_1148_index_scale_1/$entry
      -- CP-element group 392: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/array_obj_ref_1148_index_scale_1/$exit
      -- CP-element group 392: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/array_obj_ref_1148_index_resize_1/index_resize_req
      -- CP-element group 392: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/array_obj_ref_1148_index_resize_1/$exit
      -- CP-element group 392: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/array_obj_ref_1148_final_index_sum_regn_Sample/$entry
      -- CP-element group 392: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/array_obj_ref_1148_index_computed_1
      -- CP-element group 392: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/array_obj_ref_1148_index_resize_1/$entry
      -- CP-element group 392: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/array_obj_ref_1148_index_scaled_1
      -- CP-element group 392: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/array_obj_ref_1148_index_resized_1
      -- CP-element group 392: 	 branch_block_stmt_436/merge_stmt_1115__exit__
      -- CP-element group 392: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154__entry__
      -- CP-element group 392: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/array_obj_ref_1148_index_scale_1/scale_rename_req
      -- CP-element group 392: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/array_obj_ref_1148_index_scale_1/scale_rename_ack
      -- CP-element group 392: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/array_obj_ref_1148_final_index_sum_regn_Sample/req
      -- CP-element group 392: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/array_obj_ref_1148_final_index_sum_regn_update_start
      -- CP-element group 392: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/addr_of_1149_update_start_
      -- CP-element group 392: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/$entry
      -- CP-element group 392: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/array_obj_ref_1148_final_index_sum_regn_Update/req
      -- CP-element group 392: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/ptr_deref_1152_update_start_
      -- CP-element group 392: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/ptr_deref_1152_Update/word_access_complete/word_0/cr
      -- CP-element group 392: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/ptr_deref_1152_Update/word_access_complete/word_0/$entry
      -- CP-element group 392: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/ptr_deref_1152_Update/word_access_complete/$entry
      -- CP-element group 392: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/ptr_deref_1152_Update/$entry
      -- CP-element group 392: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/addr_of_1149_complete/req
      -- CP-element group 392: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/addr_of_1149_complete/$entry
      -- CP-element group 392: 	 branch_block_stmt_436/assign_stmt_1126_to_assign_stmt_1154/array_obj_ref_1148_final_index_sum_regn_Update/$entry
      -- CP-element group 392: 	 branch_block_stmt_436/merge_stmt_1115_PhiAck/$exit
      -- CP-element group 392: 	 branch_block_stmt_436/merge_stmt_1115_PhiAck/phi_stmt_1116_ack
      -- 
    phi_stmt_1116_ack_3976_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 392_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1116_ack_0, ack => convolution3D_CP_1120_elements(392)); -- 
    req_2608_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2608_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(392), ack => array_obj_ref_1148_index_offset_req_0); -- 
    req_2613_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2613_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(392), ack => array_obj_ref_1148_index_offset_req_1); -- 
    cr_2678_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2678_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(392), ack => ptr_deref_1152_store_0_req_1); -- 
    req_2628_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2628_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(392), ack => addr_of_1149_final_reg_req_1); -- 
    -- CP-element group 393:  merge  fork  transition  place  output  bypass 
    -- CP-element group 393: predecessors 
    -- CP-element group 393: 	199 
    -- CP-element group 393: 	218 
    -- CP-element group 393: successors 
    -- CP-element group 393: 	219 
    -- CP-element group 393: 	220 
    -- CP-element group 393: 	221 
    -- CP-element group 393: 	222 
    -- CP-element group 393: 	223 
    -- CP-element group 393: 	224 
    -- CP-element group 393: 	225 
    -- CP-element group 393: 	226 
    -- CP-element group 393:  members (31) 
      -- CP-element group 393: 	 branch_block_stmt_436/assign_stmt_1160_to_assign_stmt_1208/type_cast_1159_Update/cr
      -- CP-element group 393: 	 branch_block_stmt_436/assign_stmt_1160_to_assign_stmt_1208/type_cast_1159_Update/$entry
      -- CP-element group 393: 	 branch_block_stmt_436/assign_stmt_1160_to_assign_stmt_1208/type_cast_1171_sample_start_
      -- CP-element group 393: 	 branch_block_stmt_436/assign_stmt_1160_to_assign_stmt_1208/type_cast_1167_update_start_
      -- CP-element group 393: 	 branch_block_stmt_436/assign_stmt_1160_to_assign_stmt_1208/type_cast_1171_update_start_
      -- CP-element group 393: 	 branch_block_stmt_436/assign_stmt_1160_to_assign_stmt_1208/type_cast_1171_Update/cr
      -- CP-element group 393: 	 branch_block_stmt_436/assign_stmt_1160_to_assign_stmt_1208/type_cast_1163_Update/cr
      -- CP-element group 393: 	 branch_block_stmt_436/assign_stmt_1160_to_assign_stmt_1208/type_cast_1159_Sample/rr
      -- CP-element group 393: 	 branch_block_stmt_436/assign_stmt_1160_to_assign_stmt_1208/type_cast_1167_Update/$entry
      -- CP-element group 393: 	 branch_block_stmt_436/assign_stmt_1160_to_assign_stmt_1208/type_cast_1167_sample_start_
      -- CP-element group 393: 	 branch_block_stmt_436/merge_stmt_1156__exit__
      -- CP-element group 393: 	 branch_block_stmt_436/assign_stmt_1160_to_assign_stmt_1208__entry__
      -- CP-element group 393: 	 branch_block_stmt_436/assign_stmt_1160_to_assign_stmt_1208/type_cast_1171_Sample/$entry
      -- CP-element group 393: 	 branch_block_stmt_436/assign_stmt_1160_to_assign_stmt_1208/type_cast_1163_sample_start_
      -- CP-element group 393: 	 branch_block_stmt_436/assign_stmt_1160_to_assign_stmt_1208/type_cast_1159_Sample/$entry
      -- CP-element group 393: 	 branch_block_stmt_436/assign_stmt_1160_to_assign_stmt_1208/type_cast_1167_Sample/$entry
      -- CP-element group 393: 	 branch_block_stmt_436/assign_stmt_1160_to_assign_stmt_1208/type_cast_1163_Update/$entry
      -- CP-element group 393: 	 branch_block_stmt_436/assign_stmt_1160_to_assign_stmt_1208/type_cast_1159_update_start_
      -- CP-element group 393: 	 branch_block_stmt_436/assign_stmt_1160_to_assign_stmt_1208/type_cast_1171_Update/$entry
      -- CP-element group 393: 	 branch_block_stmt_436/assign_stmt_1160_to_assign_stmt_1208/type_cast_1163_Sample/rr
      -- CP-element group 393: 	 branch_block_stmt_436/assign_stmt_1160_to_assign_stmt_1208/type_cast_1159_sample_start_
      -- CP-element group 393: 	 branch_block_stmt_436/assign_stmt_1160_to_assign_stmt_1208/$entry
      -- CP-element group 393: 	 branch_block_stmt_436/assign_stmt_1160_to_assign_stmt_1208/type_cast_1167_Update/cr
      -- CP-element group 393: 	 branch_block_stmt_436/assign_stmt_1160_to_assign_stmt_1208/type_cast_1163_Sample/$entry
      -- CP-element group 393: 	 branch_block_stmt_436/assign_stmt_1160_to_assign_stmt_1208/type_cast_1163_update_start_
      -- CP-element group 393: 	 branch_block_stmt_436/assign_stmt_1160_to_assign_stmt_1208/type_cast_1167_Sample/rr
      -- CP-element group 393: 	 branch_block_stmt_436/assign_stmt_1160_to_assign_stmt_1208/type_cast_1171_Sample/rr
      -- CP-element group 393: 	 branch_block_stmt_436/merge_stmt_1156_PhiReqMerge
      -- CP-element group 393: 	 branch_block_stmt_436/merge_stmt_1156_PhiAck/$entry
      -- CP-element group 393: 	 branch_block_stmt_436/merge_stmt_1156_PhiAck/$exit
      -- CP-element group 393: 	 branch_block_stmt_436/merge_stmt_1156_PhiAck/dummy
      -- 
    cr_2695_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2695_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(393), ack => type_cast_1159_inst_req_1); -- 
    cr_2737_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2737_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(393), ack => type_cast_1171_inst_req_1); -- 
    cr_2709_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2709_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(393), ack => type_cast_1163_inst_req_1); -- 
    rr_2690_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2690_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(393), ack => type_cast_1159_inst_req_0); -- 
    rr_2704_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2704_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(393), ack => type_cast_1163_inst_req_0); -- 
    cr_2723_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2723_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(393), ack => type_cast_1167_inst_req_1); -- 
    rr_2718_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2718_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(393), ack => type_cast_1167_inst_req_0); -- 
    rr_2732_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2732_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(393), ack => type_cast_1171_inst_req_0); -- 
    convolution3D_CP_1120_elements(393) <= OrReduce(convolution3D_CP_1120_elements(199) & convolution3D_CP_1120_elements(218));
    -- CP-element group 394:  transition  output  delay-element  bypass 
    -- CP-element group 394: predecessors 
    -- CP-element group 394: 	242 
    -- CP-element group 394: successors 
    -- CP-element group 394: 	398 
    -- CP-element group 394:  members (5) 
      -- CP-element group 394: 	 branch_block_stmt_436/bbx_xnph_forx_xbody257_PhiReq/$exit
      -- CP-element group 394: 	 branch_block_stmt_436/bbx_xnph_forx_xbody257_PhiReq/phi_stmt_1289/$exit
      -- CP-element group 394: 	 branch_block_stmt_436/bbx_xnph_forx_xbody257_PhiReq/phi_stmt_1289/phi_stmt_1289_sources/$exit
      -- CP-element group 394: 	 branch_block_stmt_436/bbx_xnph_forx_xbody257_PhiReq/phi_stmt_1289/phi_stmt_1289_sources/type_cast_1293_konst_delay_trans
      -- CP-element group 394: 	 branch_block_stmt_436/bbx_xnph_forx_xbody257_PhiReq/phi_stmt_1289/phi_stmt_1289_req
      -- 
    phi_stmt_1289_req_4010_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1289_req_4010_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(394), ack => phi_stmt_1289_req_0); -- 
    -- Element group convolution3D_CP_1120_elements(394) is a control-delay.
    cp_element_394_delay: control_delay_element  generic map(name => " 394_delay", delay_value => 1)  port map(req => convolution3D_CP_1120_elements(242), ack => convolution3D_CP_1120_elements(394), clk => clk, reset =>reset);
    -- CP-element group 395:  transition  input  bypass 
    -- CP-element group 395: predecessors 
    -- CP-element group 395: 	307 
    -- CP-element group 395: successors 
    -- CP-element group 395: 	397 
    -- CP-element group 395:  members (2) 
      -- CP-element group 395: 	 branch_block_stmt_436/forx_xbody257_forx_xbody257_PhiReq/phi_stmt_1289/phi_stmt_1289_sources/type_cast_1295/SplitProtocol/Sample/$exit
      -- CP-element group 395: 	 branch_block_stmt_436/forx_xbody257_forx_xbody257_PhiReq/phi_stmt_1289/phi_stmt_1289_sources/type_cast_1295/SplitProtocol/Sample/ra
      -- 
    ra_4030_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 395_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1295_inst_ack_0, ack => convolution3D_CP_1120_elements(395)); -- 
    -- CP-element group 396:  transition  input  bypass 
    -- CP-element group 396: predecessors 
    -- CP-element group 396: 	307 
    -- CP-element group 396: successors 
    -- CP-element group 396: 	397 
    -- CP-element group 396:  members (2) 
      -- CP-element group 396: 	 branch_block_stmt_436/forx_xbody257_forx_xbody257_PhiReq/phi_stmt_1289/phi_stmt_1289_sources/type_cast_1295/SplitProtocol/Update/$exit
      -- CP-element group 396: 	 branch_block_stmt_436/forx_xbody257_forx_xbody257_PhiReq/phi_stmt_1289/phi_stmt_1289_sources/type_cast_1295/SplitProtocol/Update/ca
      -- 
    ca_4035_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 396_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1295_inst_ack_1, ack => convolution3D_CP_1120_elements(396)); -- 
    -- CP-element group 397:  join  transition  output  bypass 
    -- CP-element group 397: predecessors 
    -- CP-element group 397: 	395 
    -- CP-element group 397: 	396 
    -- CP-element group 397: successors 
    -- CP-element group 397: 	398 
    -- CP-element group 397:  members (6) 
      -- CP-element group 397: 	 branch_block_stmt_436/forx_xbody257_forx_xbody257_PhiReq/$exit
      -- CP-element group 397: 	 branch_block_stmt_436/forx_xbody257_forx_xbody257_PhiReq/phi_stmt_1289/$exit
      -- CP-element group 397: 	 branch_block_stmt_436/forx_xbody257_forx_xbody257_PhiReq/phi_stmt_1289/phi_stmt_1289_sources/$exit
      -- CP-element group 397: 	 branch_block_stmt_436/forx_xbody257_forx_xbody257_PhiReq/phi_stmt_1289/phi_stmt_1289_sources/type_cast_1295/$exit
      -- CP-element group 397: 	 branch_block_stmt_436/forx_xbody257_forx_xbody257_PhiReq/phi_stmt_1289/phi_stmt_1289_sources/type_cast_1295/SplitProtocol/$exit
      -- CP-element group 397: 	 branch_block_stmt_436/forx_xbody257_forx_xbody257_PhiReq/phi_stmt_1289/phi_stmt_1289_req
      -- 
    phi_stmt_1289_req_4036_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1289_req_4036_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(397), ack => phi_stmt_1289_req_1); -- 
    convolution3D_cp_element_group_397: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_397"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(395) & convolution3D_CP_1120_elements(396);
      gj_convolution3D_cp_element_group_397 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(397), clk => clk, reset => reset); --
    end block;
    -- CP-element group 398:  merge  transition  place  bypass 
    -- CP-element group 398: predecessors 
    -- CP-element group 398: 	394 
    -- CP-element group 398: 	397 
    -- CP-element group 398: successors 
    -- CP-element group 398: 	399 
    -- CP-element group 398:  members (2) 
      -- CP-element group 398: 	 branch_block_stmt_436/merge_stmt_1288_PhiReqMerge
      -- CP-element group 398: 	 branch_block_stmt_436/merge_stmt_1288_PhiAck/$entry
      -- 
    convolution3D_CP_1120_elements(398) <= OrReduce(convolution3D_CP_1120_elements(394) & convolution3D_CP_1120_elements(397));
    -- CP-element group 399:  fork  transition  place  input  output  bypass 
    -- CP-element group 399: predecessors 
    -- CP-element group 399: 	398 
    -- CP-element group 399: successors 
    -- CP-element group 399: 	243 
    -- CP-element group 399: 	244 
    -- CP-element group 399: 	246 
    -- CP-element group 399: 	247 
    -- CP-element group 399: 	252 
    -- CP-element group 399: 	259 
    -- CP-element group 399: 	266 
    -- CP-element group 399: 	273 
    -- CP-element group 399: 	280 
    -- CP-element group 399: 	287 
    -- CP-element group 399: 	294 
    -- CP-element group 399: 	301 
    -- CP-element group 399: 	304 
    -- CP-element group 399:  members (56) 
      -- CP-element group 399: 	 branch_block_stmt_436/merge_stmt_1288__exit__
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475__entry__
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/$entry
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/addr_of_1302_update_start_
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/array_obj_ref_1301_index_resized_1
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/array_obj_ref_1301_index_scaled_1
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/array_obj_ref_1301_index_computed_1
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/array_obj_ref_1301_index_resize_1/$entry
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/array_obj_ref_1301_index_resize_1/$exit
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/array_obj_ref_1301_index_resize_1/index_resize_req
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/array_obj_ref_1301_index_resize_1/index_resize_ack
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/array_obj_ref_1301_index_scale_1/$entry
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/array_obj_ref_1301_index_scale_1/$exit
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/array_obj_ref_1301_index_scale_1/scale_rename_req
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/array_obj_ref_1301_index_scale_1/scale_rename_ack
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/array_obj_ref_1301_final_index_sum_regn_update_start
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/array_obj_ref_1301_final_index_sum_regn_Sample/$entry
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/array_obj_ref_1301_final_index_sum_regn_Sample/req
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/array_obj_ref_1301_final_index_sum_regn_Update/$entry
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/array_obj_ref_1301_final_index_sum_regn_Update/req
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/addr_of_1302_complete/$entry
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/addr_of_1302_complete/req
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1305_sample_start_
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1305_Sample/$entry
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/RPIPE_maxpool_input_pipe_1305_Sample/rr
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1312_update_start_
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1312_Update/$entry
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1312_Update/cr
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1328_update_start_
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1328_Update/$entry
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1328_Update/cr
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1349_update_start_
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1349_Update/$entry
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1349_Update/cr
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1370_update_start_
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1370_Update/$entry
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1370_Update/cr
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1391_update_start_
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1391_Update/$entry
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1391_Update/cr
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1412_update_start_
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1412_Update/$entry
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1412_Update/cr
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1433_update_start_
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1433_Update/$entry
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1433_Update/cr
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1454_update_start_
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1454_Update/$entry
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/type_cast_1454_Update/cr
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/ptr_deref_1462_update_start_
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/ptr_deref_1462_Update/$entry
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/ptr_deref_1462_Update/word_access_complete/$entry
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/ptr_deref_1462_Update/word_access_complete/word_0/$entry
      -- CP-element group 399: 	 branch_block_stmt_436/assign_stmt_1303_to_assign_stmt_1475/ptr_deref_1462_Update/word_access_complete/word_0/cr
      -- CP-element group 399: 	 branch_block_stmt_436/merge_stmt_1288_PhiAck/$exit
      -- CP-element group 399: 	 branch_block_stmt_436/merge_stmt_1288_PhiAck/phi_stmt_1289_ack
      -- 
    phi_stmt_1289_ack_4041_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 399_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1289_ack_0, ack => convolution3D_CP_1120_elements(399)); -- 
    req_2872_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2872_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(399), ack => array_obj_ref_1301_index_offset_req_0); -- 
    req_2877_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2877_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(399), ack => array_obj_ref_1301_index_offset_req_1); -- 
    req_2892_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2892_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(399), ack => addr_of_1302_final_reg_req_1); -- 
    rr_2901_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2901_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(399), ack => RPIPE_maxpool_input_pipe_1305_inst_req_0); -- 
    cr_2934_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2934_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(399), ack => type_cast_1312_inst_req_1); -- 
    cr_2976_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2976_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(399), ack => type_cast_1328_inst_req_1); -- 
    cr_3018_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3018_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(399), ack => type_cast_1349_inst_req_1); -- 
    cr_3060_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3060_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(399), ack => type_cast_1370_inst_req_1); -- 
    cr_3102_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3102_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(399), ack => type_cast_1391_inst_req_1); -- 
    cr_3144_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3144_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(399), ack => type_cast_1412_inst_req_1); -- 
    cr_3186_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3186_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(399), ack => type_cast_1433_inst_req_1); -- 
    cr_3228_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3228_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(399), ack => type_cast_1454_inst_req_1); -- 
    cr_3278_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3278_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(399), ack => ptr_deref_1462_store_0_req_1); -- 
    -- CP-element group 400:  transition  input  bypass 
    -- CP-element group 400: predecessors 
    -- CP-element group 400: 	306 
    -- CP-element group 400: successors 
    -- CP-element group 400: 	402 
    -- CP-element group 400:  members (2) 
      -- CP-element group 400: 	 branch_block_stmt_436/forx_xcond250x_xforx_xend341_crit_edge_forx_xend341_PhiReq/phi_stmt_1507/phi_stmt_1507_sources/type_cast_1510/SplitProtocol/Sample/$exit
      -- CP-element group 400: 	 branch_block_stmt_436/forx_xcond250x_xforx_xend341_crit_edge_forx_xend341_PhiReq/phi_stmt_1507/phi_stmt_1507_sources/type_cast_1510/SplitProtocol/Sample/ra
      -- 
    ra_4073_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 400_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1510_inst_ack_0, ack => convolution3D_CP_1120_elements(400)); -- 
    -- CP-element group 401:  transition  input  bypass 
    -- CP-element group 401: predecessors 
    -- CP-element group 401: 	306 
    -- CP-element group 401: successors 
    -- CP-element group 401: 	402 
    -- CP-element group 401:  members (2) 
      -- CP-element group 401: 	 branch_block_stmt_436/forx_xcond250x_xforx_xend341_crit_edge_forx_xend341_PhiReq/phi_stmt_1507/phi_stmt_1507_sources/type_cast_1510/SplitProtocol/Update/$exit
      -- CP-element group 401: 	 branch_block_stmt_436/forx_xcond250x_xforx_xend341_crit_edge_forx_xend341_PhiReq/phi_stmt_1507/phi_stmt_1507_sources/type_cast_1510/SplitProtocol/Update/ca
      -- 
    ca_4078_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 401_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1510_inst_ack_1, ack => convolution3D_CP_1120_elements(401)); -- 
    -- CP-element group 402:  join  transition  output  bypass 
    -- CP-element group 402: predecessors 
    -- CP-element group 402: 	400 
    -- CP-element group 402: 	401 
    -- CP-element group 402: successors 
    -- CP-element group 402: 	404 
    -- CP-element group 402:  members (6) 
      -- CP-element group 402: 	 branch_block_stmt_436/forx_xcond250x_xforx_xend341_crit_edge_forx_xend341_PhiReq/$exit
      -- CP-element group 402: 	 branch_block_stmt_436/forx_xcond250x_xforx_xend341_crit_edge_forx_xend341_PhiReq/phi_stmt_1507/$exit
      -- CP-element group 402: 	 branch_block_stmt_436/forx_xcond250x_xforx_xend341_crit_edge_forx_xend341_PhiReq/phi_stmt_1507/phi_stmt_1507_sources/$exit
      -- CP-element group 402: 	 branch_block_stmt_436/forx_xcond250x_xforx_xend341_crit_edge_forx_xend341_PhiReq/phi_stmt_1507/phi_stmt_1507_sources/type_cast_1510/$exit
      -- CP-element group 402: 	 branch_block_stmt_436/forx_xcond250x_xforx_xend341_crit_edge_forx_xend341_PhiReq/phi_stmt_1507/phi_stmt_1507_sources/type_cast_1510/SplitProtocol/$exit
      -- CP-element group 402: 	 branch_block_stmt_436/forx_xcond250x_xforx_xend341_crit_edge_forx_xend341_PhiReq/phi_stmt_1507/phi_stmt_1507_req
      -- 
    phi_stmt_1507_req_4079_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1507_req_4079_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(402), ack => phi_stmt_1507_req_0); -- 
    convolution3D_cp_element_group_402: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_402"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(400) & convolution3D_CP_1120_elements(401);
      gj_convolution3D_cp_element_group_402 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(402), clk => clk, reset => reset); --
    end block;
    -- CP-element group 403:  transition  output  delay-element  bypass 
    -- CP-element group 403: predecessors 
    -- CP-element group 403: 	229 
    -- CP-element group 403: successors 
    -- CP-element group 403: 	404 
    -- CP-element group 403:  members (5) 
      -- CP-element group 403: 	 branch_block_stmt_436/ifx_xend_forx_xend341_PhiReq/$exit
      -- CP-element group 403: 	 branch_block_stmt_436/ifx_xend_forx_xend341_PhiReq/phi_stmt_1507/$exit
      -- CP-element group 403: 	 branch_block_stmt_436/ifx_xend_forx_xend341_PhiReq/phi_stmt_1507/phi_stmt_1507_sources/$exit
      -- CP-element group 403: 	 branch_block_stmt_436/ifx_xend_forx_xend341_PhiReq/phi_stmt_1507/phi_stmt_1507_sources/type_cast_1513_konst_delay_trans
      -- CP-element group 403: 	 branch_block_stmt_436/ifx_xend_forx_xend341_PhiReq/phi_stmt_1507/phi_stmt_1507_req
      -- 
    phi_stmt_1507_req_4090_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1507_req_4090_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(403), ack => phi_stmt_1507_req_1); -- 
    -- Element group convolution3D_CP_1120_elements(403) is a control-delay.
    cp_element_403_delay: control_delay_element  generic map(name => " 403_delay", delay_value => 1)  port map(req => convolution3D_CP_1120_elements(229), ack => convolution3D_CP_1120_elements(403), clk => clk, reset =>reset);
    -- CP-element group 404:  merge  transition  place  bypass 
    -- CP-element group 404: predecessors 
    -- CP-element group 404: 	402 
    -- CP-element group 404: 	403 
    -- CP-element group 404: successors 
    -- CP-element group 404: 	405 
    -- CP-element group 404:  members (2) 
      -- CP-element group 404: 	 branch_block_stmt_436/merge_stmt_1506_PhiReqMerge
      -- CP-element group 404: 	 branch_block_stmt_436/merge_stmt_1506_PhiAck/$entry
      -- 
    convolution3D_CP_1120_elements(404) <= OrReduce(convolution3D_CP_1120_elements(402) & convolution3D_CP_1120_elements(403));
    -- CP-element group 405:  branch  transition  place  input  output  bypass 
    -- CP-element group 405: predecessors 
    -- CP-element group 405: 	404 
    -- CP-element group 405: successors 
    -- CP-element group 405: 	308 
    -- CP-element group 405: 	309 
    -- CP-element group 405:  members (15) 
      -- CP-element group 405: 	 branch_block_stmt_436/merge_stmt_1506__exit__
      -- CP-element group 405: 	 branch_block_stmt_436/assign_stmt_1520_to_assign_stmt_1526__entry__
      -- CP-element group 405: 	 branch_block_stmt_436/assign_stmt_1520_to_assign_stmt_1526__exit__
      -- CP-element group 405: 	 branch_block_stmt_436/if_stmt_1527__entry__
      -- CP-element group 405: 	 branch_block_stmt_436/assign_stmt_1520_to_assign_stmt_1526/$entry
      -- CP-element group 405: 	 branch_block_stmt_436/assign_stmt_1520_to_assign_stmt_1526/$exit
      -- CP-element group 405: 	 branch_block_stmt_436/if_stmt_1527_dead_link/$entry
      -- CP-element group 405: 	 branch_block_stmt_436/R_tobool344_1528_place
      -- CP-element group 405: 	 branch_block_stmt_436/if_stmt_1527_else_link/$entry
      -- CP-element group 405: 	 branch_block_stmt_436/if_stmt_1527_if_link/$entry
      -- CP-element group 405: 	 branch_block_stmt_436/if_stmt_1527_eval_test/branch_req
      -- CP-element group 405: 	 branch_block_stmt_436/if_stmt_1527_eval_test/$exit
      -- CP-element group 405: 	 branch_block_stmt_436/if_stmt_1527_eval_test/$entry
      -- CP-element group 405: 	 branch_block_stmt_436/merge_stmt_1506_PhiAck/$exit
      -- CP-element group 405: 	 branch_block_stmt_436/merge_stmt_1506_PhiAck/phi_stmt_1507_ack
      -- 
    phi_stmt_1507_ack_4095_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 405_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1507_ack_0, ack => convolution3D_CP_1120_elements(405)); -- 
    branch_req_3312_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3312_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(405), ack => if_stmt_1527_branch_req_0); -- 
    -- CP-element group 406:  transition  output  delay-element  bypass 
    -- CP-element group 406: predecessors 
    -- CP-element group 406: 	311 
    -- CP-element group 406: successors 
    -- CP-element group 406: 	408 
    -- CP-element group 406:  members (4) 
      -- CP-element group 406: 	 branch_block_stmt_436/bbx_xnphx_xi420_forx_xbodyx_xi429_PhiReq/phi_stmt_1552/$exit
      -- CP-element group 406: 	 branch_block_stmt_436/bbx_xnphx_xi420_forx_xbodyx_xi429_PhiReq/phi_stmt_1552/phi_stmt_1552_sources/$exit
      -- CP-element group 406: 	 branch_block_stmt_436/bbx_xnphx_xi420_forx_xbodyx_xi429_PhiReq/phi_stmt_1552/phi_stmt_1552_sources/type_cast_1556_konst_delay_trans
      -- CP-element group 406: 	 branch_block_stmt_436/bbx_xnphx_xi420_forx_xbodyx_xi429_PhiReq/phi_stmt_1552/phi_stmt_1552_req
      -- 
    phi_stmt_1552_req_4118_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1552_req_4118_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(406), ack => phi_stmt_1552_req_0); -- 
    -- Element group convolution3D_CP_1120_elements(406) is a control-delay.
    cp_element_406_delay: control_delay_element  generic map(name => " 406_delay", delay_value => 1)  port map(req => convolution3D_CP_1120_elements(311), ack => convolution3D_CP_1120_elements(406), clk => clk, reset =>reset);
    -- CP-element group 407:  transition  output  delay-element  bypass 
    -- CP-element group 407: predecessors 
    -- CP-element group 407: 	311 
    -- CP-element group 407: successors 
    -- CP-element group 407: 	408 
    -- CP-element group 407:  members (4) 
      -- CP-element group 407: 	 branch_block_stmt_436/bbx_xnphx_xi420_forx_xbodyx_xi429_PhiReq/phi_stmt_1559/$exit
      -- CP-element group 407: 	 branch_block_stmt_436/bbx_xnphx_xi420_forx_xbodyx_xi429_PhiReq/phi_stmt_1559/phi_stmt_1559_sources/$exit
      -- CP-element group 407: 	 branch_block_stmt_436/bbx_xnphx_xi420_forx_xbodyx_xi429_PhiReq/phi_stmt_1559/phi_stmt_1559_sources/type_cast_1563_konst_delay_trans
      -- CP-element group 407: 	 branch_block_stmt_436/bbx_xnphx_xi420_forx_xbodyx_xi429_PhiReq/phi_stmt_1559/phi_stmt_1559_req
      -- 
    phi_stmt_1559_req_4126_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1559_req_4126_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(407), ack => phi_stmt_1559_req_0); -- 
    -- Element group convolution3D_CP_1120_elements(407) is a control-delay.
    cp_element_407_delay: control_delay_element  generic map(name => " 407_delay", delay_value => 1)  port map(req => convolution3D_CP_1120_elements(311), ack => convolution3D_CP_1120_elements(407), clk => clk, reset =>reset);
    -- CP-element group 408:  join  transition  bypass 
    -- CP-element group 408: predecessors 
    -- CP-element group 408: 	406 
    -- CP-element group 408: 	407 
    -- CP-element group 408: successors 
    -- CP-element group 408: 	416 
    -- CP-element group 408:  members (1) 
      -- CP-element group 408: 	 branch_block_stmt_436/bbx_xnphx_xi420_forx_xbodyx_xi429_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_408: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_408"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(406) & convolution3D_CP_1120_elements(407);
      gj_convolution3D_cp_element_group_408 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(408), clk => clk, reset => reset); --
    end block;
    -- CP-element group 409:  transition  input  bypass 
    -- CP-element group 409: predecessors 
    -- CP-element group 409: 	321 
    -- CP-element group 409: successors 
    -- CP-element group 409: 	411 
    -- CP-element group 409:  members (2) 
      -- CP-element group 409: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1552/phi_stmt_1552_sources/type_cast_1558/SplitProtocol/Sample/$exit
      -- CP-element group 409: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1552/phi_stmt_1552_sources/type_cast_1558/SplitProtocol/Sample/ra
      -- 
    ra_4146_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 409_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1558_inst_ack_0, ack => convolution3D_CP_1120_elements(409)); -- 
    -- CP-element group 410:  transition  input  bypass 
    -- CP-element group 410: predecessors 
    -- CP-element group 410: 	321 
    -- CP-element group 410: successors 
    -- CP-element group 410: 	411 
    -- CP-element group 410:  members (2) 
      -- CP-element group 410: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1552/phi_stmt_1552_sources/type_cast_1558/SplitProtocol/Update/$exit
      -- CP-element group 410: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1552/phi_stmt_1552_sources/type_cast_1558/SplitProtocol/Update/ca
      -- 
    ca_4151_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 410_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1558_inst_ack_1, ack => convolution3D_CP_1120_elements(410)); -- 
    -- CP-element group 411:  join  transition  output  bypass 
    -- CP-element group 411: predecessors 
    -- CP-element group 411: 	410 
    -- CP-element group 411: 	409 
    -- CP-element group 411: successors 
    -- CP-element group 411: 	415 
    -- CP-element group 411:  members (5) 
      -- CP-element group 411: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1552/$exit
      -- CP-element group 411: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1552/phi_stmt_1552_sources/$exit
      -- CP-element group 411: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1552/phi_stmt_1552_sources/type_cast_1558/$exit
      -- CP-element group 411: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1552/phi_stmt_1552_sources/type_cast_1558/SplitProtocol/$exit
      -- CP-element group 411: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1552/phi_stmt_1552_req
      -- 
    phi_stmt_1552_req_4152_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1552_req_4152_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(411), ack => phi_stmt_1552_req_1); -- 
    convolution3D_cp_element_group_411: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_411"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(410) & convolution3D_CP_1120_elements(409);
      gj_convolution3D_cp_element_group_411 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(411), clk => clk, reset => reset); --
    end block;
    -- CP-element group 412:  transition  input  bypass 
    -- CP-element group 412: predecessors 
    -- CP-element group 412: 	321 
    -- CP-element group 412: successors 
    -- CP-element group 412: 	414 
    -- CP-element group 412:  members (2) 
      -- CP-element group 412: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1559/phi_stmt_1559_sources/type_cast_1565/SplitProtocol/Sample/$exit
      -- CP-element group 412: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1559/phi_stmt_1559_sources/type_cast_1565/SplitProtocol/Sample/ra
      -- 
    ra_4169_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 412_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1565_inst_ack_0, ack => convolution3D_CP_1120_elements(412)); -- 
    -- CP-element group 413:  transition  input  bypass 
    -- CP-element group 413: predecessors 
    -- CP-element group 413: 	321 
    -- CP-element group 413: successors 
    -- CP-element group 413: 	414 
    -- CP-element group 413:  members (2) 
      -- CP-element group 413: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1559/phi_stmt_1559_sources/type_cast_1565/SplitProtocol/Update/$exit
      -- CP-element group 413: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1559/phi_stmt_1559_sources/type_cast_1565/SplitProtocol/Update/ca
      -- 
    ca_4174_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 413_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1565_inst_ack_1, ack => convolution3D_CP_1120_elements(413)); -- 
    -- CP-element group 414:  join  transition  output  bypass 
    -- CP-element group 414: predecessors 
    -- CP-element group 414: 	412 
    -- CP-element group 414: 	413 
    -- CP-element group 414: successors 
    -- CP-element group 414: 	415 
    -- CP-element group 414:  members (5) 
      -- CP-element group 414: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1559/$exit
      -- CP-element group 414: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1559/phi_stmt_1559_sources/$exit
      -- CP-element group 414: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1559/phi_stmt_1559_sources/type_cast_1565/$exit
      -- CP-element group 414: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1559/phi_stmt_1559_sources/type_cast_1565/SplitProtocol/$exit
      -- CP-element group 414: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/phi_stmt_1559/phi_stmt_1559_req
      -- 
    phi_stmt_1559_req_4175_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1559_req_4175_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(414), ack => phi_stmt_1559_req_1); -- 
    convolution3D_cp_element_group_414: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_414"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(412) & convolution3D_CP_1120_elements(413);
      gj_convolution3D_cp_element_group_414 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(414), clk => clk, reset => reset); --
    end block;
    -- CP-element group 415:  join  transition  bypass 
    -- CP-element group 415: predecessors 
    -- CP-element group 415: 	411 
    -- CP-element group 415: 	414 
    -- CP-element group 415: successors 
    -- CP-element group 415: 	416 
    -- CP-element group 415:  members (1) 
      -- CP-element group 415: 	 branch_block_stmt_436/forx_xbodyx_xi429_forx_xbodyx_xi429_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_415: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_415"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(411) & convolution3D_CP_1120_elements(414);
      gj_convolution3D_cp_element_group_415 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(415), clk => clk, reset => reset); --
    end block;
    -- CP-element group 416:  merge  fork  transition  place  bypass 
    -- CP-element group 416: predecessors 
    -- CP-element group 416: 	415 
    -- CP-element group 416: 	408 
    -- CP-element group 416: successors 
    -- CP-element group 416: 	417 
    -- CP-element group 416: 	418 
    -- CP-element group 416:  members (2) 
      -- CP-element group 416: 	 branch_block_stmt_436/merge_stmt_1551_PhiReqMerge
      -- CP-element group 416: 	 branch_block_stmt_436/merge_stmt_1551_PhiAck/$entry
      -- 
    convolution3D_CP_1120_elements(416) <= OrReduce(convolution3D_CP_1120_elements(415) & convolution3D_CP_1120_elements(408));
    -- CP-element group 417:  transition  input  bypass 
    -- CP-element group 417: predecessors 
    -- CP-element group 417: 	416 
    -- CP-element group 417: successors 
    -- CP-element group 417: 	419 
    -- CP-element group 417:  members (1) 
      -- CP-element group 417: 	 branch_block_stmt_436/merge_stmt_1551_PhiAck/phi_stmt_1552_ack
      -- 
    phi_stmt_1552_ack_4180_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 417_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1552_ack_0, ack => convolution3D_CP_1120_elements(417)); -- 
    -- CP-element group 418:  transition  input  bypass 
    -- CP-element group 418: predecessors 
    -- CP-element group 418: 	416 
    -- CP-element group 418: successors 
    -- CP-element group 418: 	419 
    -- CP-element group 418:  members (1) 
      -- CP-element group 418: 	 branch_block_stmt_436/merge_stmt_1551_PhiAck/phi_stmt_1559_ack
      -- 
    phi_stmt_1559_ack_4181_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 418_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1559_ack_0, ack => convolution3D_CP_1120_elements(418)); -- 
    -- CP-element group 419:  join  fork  transition  place  output  bypass 
    -- CP-element group 419: predecessors 
    -- CP-element group 419: 	417 
    -- CP-element group 419: 	418 
    -- CP-element group 419: successors 
    -- CP-element group 419: 	312 
    -- CP-element group 419: 	317 
    -- CP-element group 419: 	318 
    -- CP-element group 419: 	319 
    -- CP-element group 419:  members (16) 
      -- CP-element group 419: 	 branch_block_stmt_436/merge_stmt_1551__exit__
      -- CP-element group 419: 	 branch_block_stmt_436/assign_stmt_1572_to_assign_stmt_1608__entry__
      -- CP-element group 419: 	 branch_block_stmt_436/assign_stmt_1572_to_assign_stmt_1608/RPIPE_maxpool_input_pipe_1580_Sample/$entry
      -- CP-element group 419: 	 branch_block_stmt_436/assign_stmt_1572_to_assign_stmt_1608/RPIPE_maxpool_input_pipe_1580_Sample/rr
      -- CP-element group 419: 	 branch_block_stmt_436/assign_stmt_1572_to_assign_stmt_1608/RPIPE_maxpool_input_pipe_1580_sample_start_
      -- CP-element group 419: 	 branch_block_stmt_436/assign_stmt_1572_to_assign_stmt_1608/$entry
      -- CP-element group 419: 	 branch_block_stmt_436/assign_stmt_1572_to_assign_stmt_1608/type_cast_1602_Update/cr
      -- CP-element group 419: 	 branch_block_stmt_436/assign_stmt_1572_to_assign_stmt_1608/type_cast_1602_Update/$entry
      -- CP-element group 419: 	 branch_block_stmt_436/assign_stmt_1572_to_assign_stmt_1608/type_cast_1602_Sample/rr
      -- CP-element group 419: 	 branch_block_stmt_436/assign_stmt_1572_to_assign_stmt_1608/type_cast_1602_Sample/$entry
      -- CP-element group 419: 	 branch_block_stmt_436/assign_stmt_1572_to_assign_stmt_1608/type_cast_1602_update_start_
      -- CP-element group 419: 	 branch_block_stmt_436/assign_stmt_1572_to_assign_stmt_1608/type_cast_1602_sample_start_
      -- CP-element group 419: 	 branch_block_stmt_436/assign_stmt_1572_to_assign_stmt_1608/type_cast_1587_Update/cr
      -- CP-element group 419: 	 branch_block_stmt_436/assign_stmt_1572_to_assign_stmt_1608/type_cast_1587_Update/$entry
      -- CP-element group 419: 	 branch_block_stmt_436/assign_stmt_1572_to_assign_stmt_1608/type_cast_1587_update_start_
      -- CP-element group 419: 	 branch_block_stmt_436/merge_stmt_1551_PhiAck/$exit
      -- 
    rr_3351_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3351_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(419), ack => RPIPE_maxpool_input_pipe_1580_inst_req_0); -- 
    cr_3398_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3398_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(419), ack => type_cast_1602_inst_req_1); -- 
    rr_3393_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3393_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(419), ack => type_cast_1602_inst_req_0); -- 
    cr_3384_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3384_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(419), ack => type_cast_1587_inst_req_1); -- 
    convolution3D_cp_element_group_419: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_419"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(417) & convolution3D_CP_1120_elements(418);
      gj_convolution3D_cp_element_group_419 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(419), clk => clk, reset => reset); --
    end block;
    -- CP-element group 420:  transition  input  bypass 
    -- CP-element group 420: predecessors 
    -- CP-element group 420: 	322 
    -- CP-element group 420: successors 
    -- CP-element group 420: 	422 
    -- CP-element group 420:  members (2) 
      -- CP-element group 420: 	 branch_block_stmt_436/forx_xbodyx_xi429_getRemainingElementsx_xexit437_PhiReq/phi_stmt_1616/phi_stmt_1616_sources/type_cast_1619/SplitProtocol/Sample/$exit
      -- CP-element group 420: 	 branch_block_stmt_436/forx_xbodyx_xi429_getRemainingElementsx_xexit437_PhiReq/phi_stmt_1616/phi_stmt_1616_sources/type_cast_1619/SplitProtocol/Sample/ra
      -- 
    ra_4205_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 420_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1619_inst_ack_0, ack => convolution3D_CP_1120_elements(420)); -- 
    -- CP-element group 421:  transition  input  bypass 
    -- CP-element group 421: predecessors 
    -- CP-element group 421: 	322 
    -- CP-element group 421: successors 
    -- CP-element group 421: 	422 
    -- CP-element group 421:  members (2) 
      -- CP-element group 421: 	 branch_block_stmt_436/forx_xbodyx_xi429_getRemainingElementsx_xexit437_PhiReq/phi_stmt_1616/phi_stmt_1616_sources/type_cast_1619/SplitProtocol/Update/$exit
      -- CP-element group 421: 	 branch_block_stmt_436/forx_xbodyx_xi429_getRemainingElementsx_xexit437_PhiReq/phi_stmt_1616/phi_stmt_1616_sources/type_cast_1619/SplitProtocol/Update/ca
      -- 
    ca_4210_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 421_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1619_inst_ack_1, ack => convolution3D_CP_1120_elements(421)); -- 
    -- CP-element group 422:  join  transition  place  output  bypass 
    -- CP-element group 422: predecessors 
    -- CP-element group 422: 	420 
    -- CP-element group 422: 	421 
    -- CP-element group 422: successors 
    -- CP-element group 422: 	423 
    -- CP-element group 422:  members (8) 
      -- CP-element group 422: 	 branch_block_stmt_436/forx_xbodyx_xi429_getRemainingElementsx_xexit437_PhiReq/$exit
      -- CP-element group 422: 	 branch_block_stmt_436/forx_xbodyx_xi429_getRemainingElementsx_xexit437_PhiReq/phi_stmt_1616/$exit
      -- CP-element group 422: 	 branch_block_stmt_436/forx_xbodyx_xi429_getRemainingElementsx_xexit437_PhiReq/phi_stmt_1616/phi_stmt_1616_sources/$exit
      -- CP-element group 422: 	 branch_block_stmt_436/forx_xbodyx_xi429_getRemainingElementsx_xexit437_PhiReq/phi_stmt_1616/phi_stmt_1616_sources/type_cast_1619/$exit
      -- CP-element group 422: 	 branch_block_stmt_436/forx_xbodyx_xi429_getRemainingElementsx_xexit437_PhiReq/phi_stmt_1616/phi_stmt_1616_sources/type_cast_1619/SplitProtocol/$exit
      -- CP-element group 422: 	 branch_block_stmt_436/forx_xbodyx_xi429_getRemainingElementsx_xexit437_PhiReq/phi_stmt_1616/phi_stmt_1616_req
      -- CP-element group 422: 	 branch_block_stmt_436/merge_stmt_1615_PhiReqMerge
      -- CP-element group 422: 	 branch_block_stmt_436/merge_stmt_1615_PhiAck/$entry
      -- 
    phi_stmt_1616_req_4211_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1616_req_4211_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(422), ack => phi_stmt_1616_req_0); -- 
    convolution3D_cp_element_group_422: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_422"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(420) & convolution3D_CP_1120_elements(421);
      gj_convolution3D_cp_element_group_422 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(422), clk => clk, reset => reset); --
    end block;
    -- CP-element group 423:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 423: predecessors 
    -- CP-element group 423: 	422 
    -- CP-element group 423: successors 
    -- CP-element group 423: 	323 
    -- CP-element group 423: 	324 
    -- CP-element group 423: 	326 
    -- CP-element group 423: 	328 
    -- CP-element group 423:  members (29) 
      -- CP-element group 423: 	 branch_block_stmt_436/merge_stmt_1615__exit__
      -- CP-element group 423: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654__entry__
      -- CP-element group 423: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/array_obj_ref_1648_final_index_sum_regn_Update/$entry
      -- CP-element group 423: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/array_obj_ref_1648_index_resized_1
      -- CP-element group 423: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/array_obj_ref_1648_index_scaled_1
      -- CP-element group 423: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/ptr_deref_1652_Update/$entry
      -- CP-element group 423: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/array_obj_ref_1648_index_computed_1
      -- CP-element group 423: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/array_obj_ref_1648_index_resize_1/$entry
      -- CP-element group 423: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/array_obj_ref_1648_index_resize_1/$exit
      -- CP-element group 423: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/array_obj_ref_1648_index_resize_1/index_resize_req
      -- CP-element group 423: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/array_obj_ref_1648_index_resize_1/index_resize_ack
      -- CP-element group 423: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/array_obj_ref_1648_index_scale_1/$entry
      -- CP-element group 423: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/array_obj_ref_1648_index_scale_1/$exit
      -- CP-element group 423: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/array_obj_ref_1648_index_scale_1/scale_rename_req
      -- CP-element group 423: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/ptr_deref_1652_Update/word_access_complete/$entry
      -- CP-element group 423: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/array_obj_ref_1648_index_scale_1/scale_rename_ack
      -- CP-element group 423: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/array_obj_ref_1648_final_index_sum_regn_update_start
      -- CP-element group 423: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/ptr_deref_1652_Update/word_access_complete/word_0/$entry
      -- CP-element group 423: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/array_obj_ref_1648_final_index_sum_regn_Sample/req
      -- CP-element group 423: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/array_obj_ref_1648_final_index_sum_regn_Sample/$entry
      -- CP-element group 423: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/addr_of_1649_update_start_
      -- CP-element group 423: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/$entry
      -- CP-element group 423: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/ptr_deref_1652_update_start_
      -- CP-element group 423: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/addr_of_1649_complete/req
      -- CP-element group 423: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/addr_of_1649_complete/$entry
      -- CP-element group 423: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/ptr_deref_1652_Update/word_access_complete/word_0/cr
      -- CP-element group 423: 	 branch_block_stmt_436/assign_stmt_1626_to_assign_stmt_1654/array_obj_ref_1648_final_index_sum_regn_Update/req
      -- CP-element group 423: 	 branch_block_stmt_436/merge_stmt_1615_PhiAck/$exit
      -- CP-element group 423: 	 branch_block_stmt_436/merge_stmt_1615_PhiAck/phi_stmt_1616_ack
      -- 
    phi_stmt_1616_ack_4216_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 423_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1616_ack_0, ack => convolution3D_CP_1120_elements(423)); -- 
    req_3446_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3446_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(423), ack => array_obj_ref_1648_index_offset_req_0); -- 
    req_3466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(423), ack => addr_of_1649_final_reg_req_1); -- 
    cr_3516_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3516_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(423), ack => ptr_deref_1652_store_0_req_1); -- 
    req_3451_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3451_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(423), ack => array_obj_ref_1648_index_offset_req_1); -- 
    -- CP-element group 424:  merge  fork  transition  place  output  bypass 
    -- CP-element group 424: predecessors 
    -- CP-element group 424: 	308 
    -- CP-element group 424: 	329 
    -- CP-element group 424: successors 
    -- CP-element group 424: 	330 
    -- CP-element group 424: 	331 
    -- CP-element group 424:  members (13) 
      -- CP-element group 424: 	 branch_block_stmt_436/merge_stmt_1656__exit__
      -- CP-element group 424: 	 branch_block_stmt_436/call_stmt_1659__entry__
      -- CP-element group 424: 	 branch_block_stmt_436/call_stmt_1659/call_stmt_1659_Update/ccr
      -- CP-element group 424: 	 branch_block_stmt_436/call_stmt_1659/call_stmt_1659_Update/$entry
      -- CP-element group 424: 	 branch_block_stmt_436/call_stmt_1659/call_stmt_1659_Sample/crr
      -- CP-element group 424: 	 branch_block_stmt_436/call_stmt_1659/call_stmt_1659_Sample/$entry
      -- CP-element group 424: 	 branch_block_stmt_436/call_stmt_1659/call_stmt_1659_update_start_
      -- CP-element group 424: 	 branch_block_stmt_436/call_stmt_1659/call_stmt_1659_sample_start_
      -- CP-element group 424: 	 branch_block_stmt_436/call_stmt_1659/$entry
      -- CP-element group 424: 	 branch_block_stmt_436/merge_stmt_1656_PhiReqMerge
      -- CP-element group 424: 	 branch_block_stmt_436/merge_stmt_1656_PhiAck/$entry
      -- CP-element group 424: 	 branch_block_stmt_436/merge_stmt_1656_PhiAck/$exit
      -- CP-element group 424: 	 branch_block_stmt_436/merge_stmt_1656_PhiAck/dummy
      -- 
    ccr_3533_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3533_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(424), ack => call_stmt_1659_call_req_1); -- 
    crr_3528_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3528_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(424), ack => call_stmt_1659_call_req_0); -- 
    convolution3D_CP_1120_elements(424) <= OrReduce(convolution3D_CP_1120_elements(308) & convolution3D_CP_1120_elements(329));
    -- CP-element group 425:  transition  output  delay-element  bypass 
    -- CP-element group 425: predecessors 
    -- CP-element group 425: 	342 
    -- CP-element group 425: successors 
    -- CP-element group 425: 	429 
    -- CP-element group 425:  members (5) 
      -- CP-element group 425: 	 branch_block_stmt_436/ifx_xend353_whilex_xbody_PhiReq/$exit
      -- CP-element group 425: 	 branch_block_stmt_436/ifx_xend353_whilex_xbody_PhiReq/phi_stmt_1726/$exit
      -- CP-element group 425: 	 branch_block_stmt_436/ifx_xend353_whilex_xbody_PhiReq/phi_stmt_1726/phi_stmt_1726_sources/$exit
      -- CP-element group 425: 	 branch_block_stmt_436/ifx_xend353_whilex_xbody_PhiReq/phi_stmt_1726/phi_stmt_1726_sources/type_cast_1732_konst_delay_trans
      -- CP-element group 425: 	 branch_block_stmt_436/ifx_xend353_whilex_xbody_PhiReq/phi_stmt_1726/phi_stmt_1726_req
      -- 
    phi_stmt_1726_req_4238_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1726_req_4238_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(425), ack => phi_stmt_1726_req_1); -- 
    -- Element group convolution3D_CP_1120_elements(425) is a control-delay.
    cp_element_425_delay: control_delay_element  generic map(name => " 425_delay", delay_value => 1)  port map(req => convolution3D_CP_1120_elements(342), ack => convolution3D_CP_1120_elements(425), clk => clk, reset =>reset);
    -- CP-element group 426:  transition  input  bypass 
    -- CP-element group 426: predecessors 
    -- CP-element group 426: 	354 
    -- CP-element group 426: successors 
    -- CP-element group 426: 	428 
    -- CP-element group 426:  members (2) 
      -- CP-element group 426: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1726/phi_stmt_1726_sources/type_cast_1729/SplitProtocol/Sample/$exit
      -- CP-element group 426: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1726/phi_stmt_1726_sources/type_cast_1729/SplitProtocol/Sample/ra
      -- 
    ra_4258_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 426_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1729_inst_ack_0, ack => convolution3D_CP_1120_elements(426)); -- 
    -- CP-element group 427:  transition  input  bypass 
    -- CP-element group 427: predecessors 
    -- CP-element group 427: 	354 
    -- CP-element group 427: successors 
    -- CP-element group 427: 	428 
    -- CP-element group 427:  members (2) 
      -- CP-element group 427: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1726/phi_stmt_1726_sources/type_cast_1729/SplitProtocol/Update/$exit
      -- CP-element group 427: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1726/phi_stmt_1726_sources/type_cast_1729/SplitProtocol/Update/ca
      -- 
    ca_4263_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 427_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1729_inst_ack_1, ack => convolution3D_CP_1120_elements(427)); -- 
    -- CP-element group 428:  join  transition  output  bypass 
    -- CP-element group 428: predecessors 
    -- CP-element group 428: 	426 
    -- CP-element group 428: 	427 
    -- CP-element group 428: successors 
    -- CP-element group 428: 	429 
    -- CP-element group 428:  members (6) 
      -- CP-element group 428: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/$exit
      -- CP-element group 428: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1726/$exit
      -- CP-element group 428: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1726/phi_stmt_1726_sources/$exit
      -- CP-element group 428: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1726/phi_stmt_1726_sources/type_cast_1729/$exit
      -- CP-element group 428: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1726/phi_stmt_1726_sources/type_cast_1729/SplitProtocol/$exit
      -- CP-element group 428: 	 branch_block_stmt_436/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1726/phi_stmt_1726_req
      -- 
    phi_stmt_1726_req_4264_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1726_req_4264_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(428), ack => phi_stmt_1726_req_0); -- 
    convolution3D_cp_element_group_428: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_428"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1120_elements(426) & convolution3D_CP_1120_elements(427);
      gj_convolution3D_cp_element_group_428 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1120_elements(428), clk => clk, reset => reset); --
    end block;
    -- CP-element group 429:  merge  transition  place  bypass 
    -- CP-element group 429: predecessors 
    -- CP-element group 429: 	425 
    -- CP-element group 429: 	428 
    -- CP-element group 429: successors 
    -- CP-element group 429: 	430 
    -- CP-element group 429:  members (2) 
      -- CP-element group 429: 	 branch_block_stmt_436/merge_stmt_1725_PhiReqMerge
      -- CP-element group 429: 	 branch_block_stmt_436/merge_stmt_1725_PhiAck/$entry
      -- 
    convolution3D_CP_1120_elements(429) <= OrReduce(convolution3D_CP_1120_elements(425) & convolution3D_CP_1120_elements(428));
    -- CP-element group 430:  fork  transition  place  input  output  bypass 
    -- CP-element group 430: predecessors 
    -- CP-element group 430: 	429 
    -- CP-element group 430: successors 
    -- CP-element group 430: 	343 
    -- CP-element group 430: 	344 
    -- CP-element group 430: 	345 
    -- CP-element group 430: 	346 
    -- CP-element group 430: 	349 
    -- CP-element group 430: 	350 
    -- CP-element group 430: 	351 
    -- CP-element group 430:  members (26) 
      -- CP-element group 430: 	 branch_block_stmt_436/merge_stmt_1725__exit__
      -- CP-element group 430: 	 branch_block_stmt_436/assign_stmt_1738_to_assign_stmt_1772__entry__
      -- CP-element group 430: 	 branch_block_stmt_436/assign_stmt_1738_to_assign_stmt_1772/type_cast_1746_Sample/$entry
      -- CP-element group 430: 	 branch_block_stmt_436/assign_stmt_1738_to_assign_stmt_1772/call_stmt_1761_update_start_
      -- CP-element group 430: 	 branch_block_stmt_436/assign_stmt_1738_to_assign_stmt_1772/call_stmt_1761_Update/$entry
      -- CP-element group 430: 	 branch_block_stmt_436/assign_stmt_1738_to_assign_stmt_1772/type_cast_1746_Sample/rr
      -- CP-element group 430: 	 branch_block_stmt_436/assign_stmt_1738_to_assign_stmt_1772/call_stmt_1754_Update/ccr
      -- CP-element group 430: 	 branch_block_stmt_436/assign_stmt_1738_to_assign_stmt_1772/type_cast_1746_update_start_
      -- CP-element group 430: 	 branch_block_stmt_436/assign_stmt_1738_to_assign_stmt_1772/call_stmt_1761_Update/ccr
      -- CP-element group 430: 	 branch_block_stmt_436/assign_stmt_1738_to_assign_stmt_1772/call_stmt_1754_update_start_
      -- CP-element group 430: 	 branch_block_stmt_436/assign_stmt_1738_to_assign_stmt_1772/type_cast_1746_sample_start_
      -- CP-element group 430: 	 branch_block_stmt_436/assign_stmt_1738_to_assign_stmt_1772/$entry
      -- CP-element group 430: 	 branch_block_stmt_436/assign_stmt_1738_to_assign_stmt_1772/call_stmt_1761_Sample/crr
      -- CP-element group 430: 	 branch_block_stmt_436/assign_stmt_1738_to_assign_stmt_1772/call_stmt_1754_Update/$entry
      -- CP-element group 430: 	 branch_block_stmt_436/assign_stmt_1738_to_assign_stmt_1772/type_cast_1750_Update/cr
      -- CP-element group 430: 	 branch_block_stmt_436/assign_stmt_1738_to_assign_stmt_1772/type_cast_1750_Update/$entry
      -- CP-element group 430: 	 branch_block_stmt_436/assign_stmt_1738_to_assign_stmt_1772/type_cast_1750_Sample/rr
      -- CP-element group 430: 	 branch_block_stmt_436/assign_stmt_1738_to_assign_stmt_1772/call_stmt_1761_sample_start_
      -- CP-element group 430: 	 branch_block_stmt_436/assign_stmt_1738_to_assign_stmt_1772/call_stmt_1761_Sample/$entry
      -- CP-element group 430: 	 branch_block_stmt_436/assign_stmt_1738_to_assign_stmt_1772/type_cast_1750_Sample/$entry
      -- CP-element group 430: 	 branch_block_stmt_436/assign_stmt_1738_to_assign_stmt_1772/type_cast_1750_update_start_
      -- CP-element group 430: 	 branch_block_stmt_436/assign_stmt_1738_to_assign_stmt_1772/type_cast_1750_sample_start_
      -- CP-element group 430: 	 branch_block_stmt_436/assign_stmt_1738_to_assign_stmt_1772/type_cast_1746_Update/cr
      -- CP-element group 430: 	 branch_block_stmt_436/assign_stmt_1738_to_assign_stmt_1772/type_cast_1746_Update/$entry
      -- CP-element group 430: 	 branch_block_stmt_436/merge_stmt_1725_PhiAck/$exit
      -- CP-element group 430: 	 branch_block_stmt_436/merge_stmt_1725_PhiAck/phi_stmt_1726_ack
      -- 
    phi_stmt_1726_ack_4269_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 430_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1726_ack_0, ack => convolution3D_CP_1120_elements(430)); -- 
    rr_3618_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3618_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(430), ack => type_cast_1746_inst_req_0); -- 
    ccr_3651_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3651_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(430), ack => call_stmt_1754_call_req_1); -- 
    ccr_3665_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3665_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(430), ack => call_stmt_1761_call_req_1); -- 
    crr_3660_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3660_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(430), ack => call_stmt_1761_call_req_0); -- 
    cr_3637_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3637_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(430), ack => type_cast_1750_inst_req_1); -- 
    rr_3632_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3632_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(430), ack => type_cast_1750_inst_req_0); -- 
    cr_3623_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3623_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1120_elements(430), ack => type_cast_1746_inst_req_1); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i64_i64_1006_wire : std_logic_vector(63 downto 0);
    signal ASHR_i64_i64_1200_wire : std_logic_vector(63 downto 0);
    signal ASHR_i64_i64_1502_wire : std_logic_vector(63 downto 0);
    signal Bx_xnot_1126 : std_logic_vector(63 downto 0);
    signal R_indvar476_1300_resized : std_logic_vector(13 downto 0);
    signal R_indvar476_1300_scaled : std_logic_vector(13 downto 0);
    signal R_indvar490_804_resized : std_logic_vector(13 downto 0);
    signal R_indvar490_804_scaled : std_logic_vector(13 downto 0);
    signal R_ix_x0x_xlcssa_1147_resized : std_logic_vector(13 downto 0);
    signal R_ix_x0x_xlcssa_1147_scaled : std_logic_vector(13 downto 0);
    signal R_ix_x1x_xlcssa_1647_resized : std_logic_vector(13 downto 0);
    signal R_ix_x1x_xlcssa_1647_scaled : std_logic_vector(13 downto 0);
    signal add117_653 : std_logic_vector(15 downto 0);
    signal add135_684 : std_logic_vector(15 downto 0);
    signal add1519x_xi434_1632 : std_logic_vector(63 downto 0);
    signal add1519x_xi_1132 : std_logic_vector(63 downto 0);
    signal add166_838 : std_logic_vector(63 downto 0);
    signal add176_859 : std_logic_vector(63 downto 0);
    signal add186_880 : std_logic_vector(63 downto 0);
    signal add196_901 : std_logic_vector(63 downto 0);
    signal add206_922 : std_logic_vector(63 downto 0);
    signal add216_943 : std_logic_vector(63 downto 0);
    signal add226_964 : std_logic_vector(63 downto 0);
    signal add273_1334 : std_logic_vector(63 downto 0);
    signal add27_498 : std_logic_vector(15 downto 0);
    signal add283_1355 : std_logic_vector(63 downto 0);
    signal add293_1376 : std_logic_vector(63 downto 0);
    signal add303_1397 : std_logic_vector(63 downto 0);
    signal add313_1418 : std_logic_vector(63 downto 0);
    signal add323_1439 : std_logic_vector(63 downto 0);
    signal add333_1460 : std_logic_vector(63 downto 0);
    signal add45_529 : std_logic_vector(15 downto 0);
    signal add63_560 : std_logic_vector(15 downto 0);
    signal add81_591 : std_logic_vector(15 downto 0);
    signal add99_622 : std_logic_vector(15 downto 0);
    signal add_467 : std_logic_vector(31 downto 0);
    signal addx_xi425_1593 : std_logic_vector(63 downto 0);
    signal addx_xi_1093 : std_logic_vector(63 downto 0);
    signal and343_1520 : std_logic_vector(63 downto 0);
    signal and_1024 : std_logic_vector(63 downto 0);
    signal array_obj_ref_1148_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1148_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1148_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1148_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1148_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1148_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1301_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1301_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1301_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1301_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1301_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1301_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1648_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1648_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1648_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1648_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1648_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1648_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_805_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_805_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_805_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_805_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_805_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_805_root_address : std_logic_vector(13 downto 0);
    signal arrayidx237_1150 : std_logic_vector(31 downto 0);
    signal arrayidx337_1303 : std_logic_vector(31 downto 0);
    signal arrayidx352_1650 : std_logic_vector(31 downto 0);
    signal arrayidx_807 : std_logic_vector(31 downto 0);
    signal call104_625 : std_logic_vector(7 downto 0);
    signal call113_641 : std_logic_vector(7 downto 0);
    signal call122_656 : std_logic_vector(7 downto 0);
    signal call131_672 : std_logic_vector(7 downto 0);
    signal call14_470 : std_logic_vector(7 downto 0);
    signal call153_810 : std_logic_vector(7 downto 0);
    signal call161_826 : std_logic_vector(7 downto 0);
    signal call171_847 : std_logic_vector(7 downto 0);
    signal call181_868 : std_logic_vector(7 downto 0);
    signal call191_889 : std_logic_vector(7 downto 0);
    signal call201_910 : std_logic_vector(7 downto 0);
    signal call211_931 : std_logic_vector(7 downto 0);
    signal call221_952 : std_logic_vector(7 downto 0);
    signal call23_486 : std_logic_vector(7 downto 0);
    signal call260_1306 : std_logic_vector(7 downto 0);
    signal call268_1322 : std_logic_vector(7 downto 0);
    signal call278_1343 : std_logic_vector(7 downto 0);
    signal call288_1364 : std_logic_vector(7 downto 0);
    signal call298_1385 : std_logic_vector(7 downto 0);
    signal call308_1406 : std_logic_vector(7 downto 0);
    signal call318_1427 : std_logic_vector(7 downto 0);
    signal call328_1448 : std_logic_vector(7 downto 0);
    signal call32_501 : std_logic_vector(7 downto 0);
    signal call355_1659 : std_logic_vector(63 downto 0);
    signal call410_1787 : std_logic_vector(63 downto 0);
    signal call41_517 : std_logic_vector(7 downto 0);
    signal call50_532 : std_logic_vector(7 downto 0);
    signal call59_548 : std_logic_vector(7 downto 0);
    signal call68_563 : std_logic_vector(7 downto 0);
    signal call6_455 : std_logic_vector(7 downto 0);
    signal call77_579 : std_logic_vector(7 downto 0);
    signal call86_594 : std_logic_vector(7 downto 0);
    signal call95_610 : std_logic_vector(7 downto 0);
    signal call_439 : std_logic_vector(7 downto 0);
    signal callx_xi423_1581 : std_logic_vector(7 downto 0);
    signal callx_xi_1081 : std_logic_vector(7 downto 0);
    signal cmp255443_1208 : std_logic_vector(0 downto 0);
    signal cmp447_714 : std_logic_vector(0 downto 0);
    signal cmpx_xi428_1608 : std_logic_vector(0 downto 0);
    signal cmpx_xi_1108 : std_logic_vector(0 downto 0);
    signal conv109_632 : std_logic_vector(15 downto 0);
    signal conv116_648 : std_logic_vector(15 downto 0);
    signal conv127_663 : std_logic_vector(15 downto 0);
    signal conv134_679 : std_logic_vector(15 downto 0);
    signal conv141_688 : std_logic_vector(31 downto 0);
    signal conv143_692 : std_logic_vector(31 downto 0);
    signal conv145_708 : std_logic_vector(63 downto 0);
    signal conv156_817 : std_logic_vector(63 downto 0);
    signal conv165_833 : std_logic_vector(63 downto 0);
    signal conv175_854 : std_logic_vector(63 downto 0);
    signal conv185_875 : std_logic_vector(63 downto 0);
    signal conv195_896 : std_logic_vector(63 downto 0);
    signal conv19_477 : std_logic_vector(15 downto 0);
    signal conv205_917 : std_logic_vector(63 downto 0);
    signal conv215_938 : std_logic_vector(63 downto 0);
    signal conv225_959 : std_logic_vector(63 downto 0);
    signal conv239_1160 : std_logic_vector(63 downto 0);
    signal conv241_1164 : std_logic_vector(63 downto 0);
    signal conv244_1168 : std_logic_vector(63 downto 0);
    signal conv247_1172 : std_logic_vector(63 downto 0);
    signal conv249_1202 : std_logic_vector(63 downto 0);
    signal conv263_1313 : std_logic_vector(63 downto 0);
    signal conv26_493 : std_logic_vector(15 downto 0);
    signal conv272_1329 : std_logic_vector(63 downto 0);
    signal conv282_1350 : std_logic_vector(63 downto 0);
    signal conv292_1371 : std_logic_vector(63 downto 0);
    signal conv2x_xi418_1543 : std_logic_vector(31 downto 0);
    signal conv2x_xi_1043 : std_logic_vector(31 downto 0);
    signal conv302_1392 : std_logic_vector(63 downto 0);
    signal conv312_1413 : std_logic_vector(63 downto 0);
    signal conv322_1434 : std_logic_vector(63 downto 0);
    signal conv332_1455 : std_logic_vector(63 downto 0);
    signal conv356_1784 : std_logic_vector(63 downto 0);
    signal conv37_508 : std_logic_vector(15 downto 0);
    signal conv381_1747 : std_logic_vector(63 downto 0);
    signal conv387_1751 : std_logic_vector(63 downto 0);
    signal conv3_446 : std_logic_vector(31 downto 0);
    signal conv411_1792 : std_logic_vector(63 downto 0);
    signal conv44_524 : std_logic_vector(15 downto 0);
    signal conv55_539 : std_logic_vector(15 downto 0);
    signal conv62_555 : std_logic_vector(15 downto 0);
    signal conv73_570 : std_logic_vector(15 downto 0);
    signal conv80_586 : std_logic_vector(15 downto 0);
    signal conv8x_xi424_1588 : std_logic_vector(63 downto 0);
    signal conv8x_xi_1088 : std_logic_vector(63 downto 0);
    signal conv91_601 : std_logic_vector(15 downto 0);
    signal conv98_617 : std_logic_vector(15 downto 0);
    signal conv9_462 : std_logic_vector(31 downto 0);
    signal convx_xi427_1603 : std_logic_vector(31 downto 0);
    signal convx_xi_1103 : std_logic_vector(31 downto 0);
    signal elementx_x024x_xi422_1559 : std_logic_vector(63 downto 0);
    signal elementx_x024x_xi_1059 : std_logic_vector(63 downto 0);
    signal exitcond32_979 : std_logic_vector(0 downto 0);
    signal exitcond5_1772 : std_logic_vector(0 downto 0);
    signal exitcond_1475 : std_logic_vector(0 downto 0);
    signal iNsTr_120_1539 : std_logic_vector(63 downto 0);
    signal iNsTr_128_1578 : std_logic_vector(15 downto 0);
    signal iNsTr_138_1626 : std_logic_vector(63 downto 0);
    signal iNsTr_82_1078 : std_logic_vector(15 downto 0);
    signal indvar476_1289 : std_logic_vector(63 downto 0);
    signal indvar490_793 : std_logic_vector(63 downto 0);
    signal indvar_1726 : std_logic_vector(31 downto 0);
    signal indvarx_xnext477_1470 : std_logic_vector(63 downto 0);
    signal indvarx_xnext491_974 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_1767 : std_logic_vector(31 downto 0);
    signal ix_x0x_xlcssa_1011 : std_logic_vector(63 downto 0);
    signal ix_x1x_xlcssa_1507 : std_logic_vector(63 downto 0);
    signal mul144_702 : std_logic_vector(31 downto 0);
    signal mul242_1177 : std_logic_vector(63 downto 0);
    signal mul245_1182 : std_logic_vector(63 downto 0);
    signal mul248_1187 : std_logic_vector(63 downto 0);
    signal mul362_1665 : std_logic_vector(15 downto 0);
    signal mul375_1670 : std_logic_vector(15 downto 0);
    signal mul380_1738 : std_logic_vector(31 downto 0);
    signal mul386_1743 : std_logic_vector(31 downto 0);
    signal mul_697 : std_logic_vector(31 downto 0);
    signal nx_x025x_xi421_1552 : std_logic_vector(15 downto 0);
    signal nx_x025x_xi_1052 : std_logic_vector(15 downto 0);
    signal phitmp451_1504 : std_logic_vector(63 downto 0);
    signal phitmp_1008 : std_logic_vector(63 downto 0);
    signal ptr_deref_1152_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1152_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1152_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1152_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1152_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1152_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1462_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1462_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1462_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1462_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1462_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1462_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1652_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1652_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1652_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1652_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1652_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1652_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_966_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_966_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_966_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_966_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_966_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_966_word_offset_0 : std_logic_vector(13 downto 0);
    signal sext_1193 : std_logic_vector(63 downto 0);
    signal sh_promx_xi435_1638 : std_logic_vector(63 downto 0);
    signal sh_promx_xi_1138 : std_logic_vector(63 downto 0);
    signal shl110_638 : std_logic_vector(15 downto 0);
    signal shl11x_xi426_1599 : std_logic_vector(63 downto 0);
    signal shl11x_xi426x_xlcssa_1616 : std_logic_vector(63 downto 0);
    signal shl11x_xi_1099 : std_logic_vector(63 downto 0);
    signal shl11x_xix_xlcssa_1116 : std_logic_vector(63 downto 0);
    signal shl128_669 : std_logic_vector(15 downto 0);
    signal shl158_823 : std_logic_vector(63 downto 0);
    signal shl168_844 : std_logic_vector(63 downto 0);
    signal shl178_865 : std_logic_vector(63 downto 0);
    signal shl17x_xi436_1643 : std_logic_vector(63 downto 0);
    signal shl17x_xi_1143 : std_logic_vector(63 downto 0);
    signal shl188_886 : std_logic_vector(63 downto 0);
    signal shl198_907 : std_logic_vector(63 downto 0);
    signal shl208_928 : std_logic_vector(63 downto 0);
    signal shl20_483 : std_logic_vector(15 downto 0);
    signal shl218_949 : std_logic_vector(63 downto 0);
    signal shl265_1319 : std_logic_vector(63 downto 0);
    signal shl275_1340 : std_logic_vector(63 downto 0);
    signal shl285_1361 : std_logic_vector(63 downto 0);
    signal shl295_1382 : std_logic_vector(63 downto 0);
    signal shl305_1403 : std_logic_vector(63 downto 0);
    signal shl315_1424 : std_logic_vector(63 downto 0);
    signal shl325_1445 : std_logic_vector(63 downto 0);
    signal shl38_514 : std_logic_vector(15 downto 0);
    signal shl56_545 : std_logic_vector(15 downto 0);
    signal shl74_576 : std_logic_vector(15 downto 0);
    signal shl92_607 : std_logic_vector(15 downto 0);
    signal shl_452 : std_logic_vector(31 downto 0);
    signal shlx_xi419_1549 : std_logic_vector(31 downto 0);
    signal shlx_xi_1049 : std_logic_vector(31 downto 0);
    signal sub395_1689 : std_logic_vector(15 downto 0);
    signal sub415_1797 : std_logic_vector(63 downto 0);
    signal sub_1683 : std_logic_vector(15 downto 0);
    signal tmp12_1231 : std_logic_vector(63 downto 0);
    signal tmp13_1235 : std_logic_vector(63 downto 0);
    signal tmp14_1240 : std_logic_vector(63 downto 0);
    signal tmp15_1244 : std_logic_vector(63 downto 0);
    signal tmp16_1249 : std_logic_vector(63 downto 0);
    signal tmp17_1253 : std_logic_vector(63 downto 0);
    signal tmp18_1258 : std_logic_vector(63 downto 0);
    signal tmp19_1262 : std_logic_vector(31 downto 0);
    signal tmp20_1267 : std_logic_vector(63 downto 0);
    signal tmp21_1273 : std_logic_vector(63 downto 0);
    signal tmp22_1279 : std_logic_vector(0 downto 0);
    signal tmp24_752 : std_logic_vector(31 downto 0);
    signal tmp25_757 : std_logic_vector(31 downto 0);
    signal tmp26_761 : std_logic_vector(31 downto 0);
    signal tmp27_766 : std_logic_vector(31 downto 0);
    signal tmp28_771 : std_logic_vector(63 downto 0);
    signal tmp29_777 : std_logic_vector(63 downto 0);
    signal tmp30_783 : std_logic_vector(0 downto 0);
    signal tmp3_1699 : std_logic_vector(31 downto 0);
    signal tmp452_1572 : std_logic_vector(15 downto 0);
    signal tmp453_1695 : std_logic_vector(15 downto 0);
    signal tmp471_1221 : std_logic_vector(63 downto 0);
    signal tmp472_1227 : std_logic_vector(0 downto 0);
    signal tmp473_1495 : std_logic_vector(63 downto 0);
    signal tmp480_726 : std_logic_vector(31 downto 0);
    signal tmp482_731 : std_logic_vector(31 downto 0);
    signal tmp483_736 : std_logic_vector(63 downto 0);
    signal tmp484_742 : std_logic_vector(63 downto 0);
    signal tmp485_748 : std_logic_vector(0 downto 0);
    signal tmp487_999 : std_logic_vector(63 downto 0);
    signal tmp4_1705 : std_logic_vector(31 downto 0);
    signal tmp6_1709 : std_logic_vector(31 downto 0);
    signal tmp7_1714 : std_logic_vector(15 downto 0);
    signal tmp8_1718 : std_logic_vector(31 downto 0);
    signal tmp9_1723 : std_logic_vector(31 downto 0);
    signal tmp_1072 : std_logic_vector(15 downto 0);
    signal tobool344_1526 : std_logic_vector(0 downto 0);
    signal tobool_1030 : std_logic_vector(0 downto 0);
    signal type_cast_1002_wire : std_logic_vector(63 downto 0);
    signal type_cast_1005_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1014_wire : std_logic_vector(63 downto 0);
    signal type_cast_1017_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1022_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1028_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1041_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1047_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1056_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1058_wire : std_logic_vector(15 downto 0);
    signal type_cast_1063_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1065_wire : std_logic_vector(63 downto 0);
    signal type_cast_1070_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1076_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1097_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1119_wire : std_logic_vector(63 downto 0);
    signal type_cast_1124_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1130_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1136_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1191_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1196_wire : std_logic_vector(63 downto 0);
    signal type_cast_1199_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1206_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1219_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1225_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1265_wire : std_logic_vector(63 downto 0);
    signal type_cast_1271_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1277_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1284_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1293_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1295_wire : std_logic_vector(63 downto 0);
    signal type_cast_1317_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1338_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1359_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1380_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1401_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1422_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1443_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1468_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1487_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1493_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1498_wire : std_logic_vector(63 downto 0);
    signal type_cast_1501_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1510_wire : std_logic_vector(63 downto 0);
    signal type_cast_1513_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1518_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1524_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1537_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1547_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1556_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1558_wire : std_logic_vector(15 downto 0);
    signal type_cast_1563_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1565_wire : std_logic_vector(63 downto 0);
    signal type_cast_1570_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1576_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1597_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1619_wire : std_logic_vector(63 downto 0);
    signal type_cast_1624_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1630_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1636_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1676_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1681_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1687_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1693_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1703_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1729_wire : std_logic_vector(31 downto 0);
    signal type_cast_1732_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1765_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1782_wire : std_logic_vector(63 downto 0);
    signal type_cast_1790_wire : std_logic_vector(63 downto 0);
    signal type_cast_450_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_481_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_512_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_543_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_574_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_605_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_636_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_667_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_706_wire : std_logic_vector(63 downto 0);
    signal type_cast_712_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_734_wire : std_logic_vector(63 downto 0);
    signal type_cast_740_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_746_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_769_wire : std_logic_vector(63 downto 0);
    signal type_cast_775_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_781_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_788_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_797_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_799_wire : std_logic_vector(63 downto 0);
    signal type_cast_821_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_842_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_863_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_884_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_905_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_926_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_947_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_972_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_991_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_997_wire_constant : std_logic_vector(63 downto 0);
    signal umax23_1286 : std_logic_vector(63 downto 0);
    signal umax31_790 : std_logic_vector(63 downto 0);
    signal umax486_993 : std_logic_vector(63 downto 0);
    signal umax_1489 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    array_obj_ref_1148_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1148_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1148_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1148_resized_base_address <= "00000000000000";
    array_obj_ref_1301_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1301_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1301_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1301_resized_base_address <= "00000000000000";
    array_obj_ref_1648_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1648_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1648_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1648_resized_base_address <= "00000000000000";
    array_obj_ref_805_constant_part_of_offset <= "00000000000000";
    array_obj_ref_805_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_805_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_805_resized_base_address <= "00000000000000";
    ptr_deref_1152_word_offset_0 <= "00000000000000";
    ptr_deref_1462_word_offset_0 <= "00000000000000";
    ptr_deref_1652_word_offset_0 <= "00000000000000";
    ptr_deref_966_word_offset_0 <= "00000000000000";
    type_cast_1005_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1017_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1022_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    type_cast_1028_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1041_wire_constant <= "00000000000000000000000000000001";
    type_cast_1047_wire_constant <= "00000000000000000000000000000110";
    type_cast_1056_wire_constant <= "0000000000000000";
    type_cast_1063_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1070_wire_constant <= "0000000000000001";
    type_cast_1076_wire_constant <= "0000000000000001";
    type_cast_1097_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1124_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000100";
    type_cast_1130_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1136_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1191_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1199_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1206_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    type_cast_1219_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_1225_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1271_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_1277_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1284_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1293_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1317_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1338_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1359_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1380_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1401_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1422_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1443_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1468_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1487_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1493_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1501_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1513_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1518_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    type_cast_1524_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1537_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1547_wire_constant <= "00000000000000000000000000000110";
    type_cast_1556_wire_constant <= "0000000000000000";
    type_cast_1563_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1570_wire_constant <= "0000000000000001";
    type_cast_1576_wire_constant <= "0000000000000001";
    type_cast_1597_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1624_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000100";
    type_cast_1630_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1636_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1676_wire_constant <= "00101100";
    type_cast_1681_wire_constant <= "1111111111111111";
    type_cast_1687_wire_constant <= "1111111111111111";
    type_cast_1693_wire_constant <= "1111111111111111";
    type_cast_1703_wire_constant <= "00000000000000000000000000000001";
    type_cast_1732_wire_constant <= "00000000000000000000000000000000";
    type_cast_1765_wire_constant <= "00000000000000000000000000000001";
    type_cast_450_wire_constant <= "00000000000000000000000000001000";
    type_cast_481_wire_constant <= "0000000000001000";
    type_cast_512_wire_constant <= "0000000000001000";
    type_cast_543_wire_constant <= "0000000000001000";
    type_cast_574_wire_constant <= "0000000000001000";
    type_cast_605_wire_constant <= "0000000000001000";
    type_cast_636_wire_constant <= "0000000000001000";
    type_cast_667_wire_constant <= "0000000000001000";
    type_cast_712_wire_constant <= "00000000000000000000000000000011";
    type_cast_740_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_746_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_775_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_781_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_788_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_797_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_821_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_842_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_863_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_884_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_905_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_926_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_947_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_972_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_991_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_997_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    phi_stmt_1011: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1014_wire & type_cast_1017_wire_constant;
      req <= phi_stmt_1011_req_0 & phi_stmt_1011_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1011",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1011_ack_0,
          idata => idata,
          odata => ix_x0x_xlcssa_1011,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1011
    phi_stmt_1052: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1056_wire_constant & type_cast_1058_wire;
      req <= phi_stmt_1052_req_0 & phi_stmt_1052_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1052",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1052_ack_0,
          idata => idata,
          odata => nx_x025x_xi_1052,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1052
    phi_stmt_1059: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1063_wire_constant & type_cast_1065_wire;
      req <= phi_stmt_1059_req_0 & phi_stmt_1059_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1059",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1059_ack_0,
          idata => idata,
          odata => elementx_x024x_xi_1059,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1059
    phi_stmt_1116: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_1119_wire;
      req(0) <= phi_stmt_1116_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1116",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1116_ack_0,
          idata => idata,
          odata => shl11x_xix_xlcssa_1116,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1116
    phi_stmt_1289: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1293_wire_constant & type_cast_1295_wire;
      req <= phi_stmt_1289_req_0 & phi_stmt_1289_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1289",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1289_ack_0,
          idata => idata,
          odata => indvar476_1289,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1289
    phi_stmt_1507: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1510_wire & type_cast_1513_wire_constant;
      req <= phi_stmt_1507_req_0 & phi_stmt_1507_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1507",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1507_ack_0,
          idata => idata,
          odata => ix_x1x_xlcssa_1507,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1507
    phi_stmt_1552: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1556_wire_constant & type_cast_1558_wire;
      req <= phi_stmt_1552_req_0 & phi_stmt_1552_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1552",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1552_ack_0,
          idata => idata,
          odata => nx_x025x_xi421_1552,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1552
    phi_stmt_1559: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1563_wire_constant & type_cast_1565_wire;
      req <= phi_stmt_1559_req_0 & phi_stmt_1559_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1559",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1559_ack_0,
          idata => idata,
          odata => elementx_x024x_xi422_1559,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1559
    phi_stmt_1616: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_1619_wire;
      req(0) <= phi_stmt_1616_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1616",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1616_ack_0,
          idata => idata,
          odata => shl11x_xi426x_xlcssa_1616,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1616
    phi_stmt_1726: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1729_wire & type_cast_1732_wire_constant;
      req <= phi_stmt_1726_req_0 & phi_stmt_1726_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1726",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1726_ack_0,
          idata => idata,
          odata => indvar_1726,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1726
    phi_stmt_793: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_797_wire_constant & type_cast_799_wire;
      req <= phi_stmt_793_req_0 & phi_stmt_793_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_793",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_793_ack_0,
          idata => idata,
          odata => indvar490_793,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_793
    -- flow-through select operator MUX_1285_inst
    umax23_1286 <= tmp21_1273 when (tmp22_1279(0) /=  '0') else type_cast_1284_wire_constant;
    -- flow-through select operator MUX_1488_inst
    umax_1489 <= tmp471_1221 when (tmp472_1227(0) /=  '0') else type_cast_1487_wire_constant;
    -- flow-through select operator MUX_789_inst
    umax31_790 <= tmp29_777 when (tmp30_783(0) /=  '0') else type_cast_788_wire_constant;
    -- flow-through select operator MUX_992_inst
    umax486_993 <= tmp484_742 when (tmp485_748(0) /=  '0') else type_cast_991_wire_constant;
    addr_of_1149_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1149_final_reg_req_0;
      addr_of_1149_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1149_final_reg_req_1;
      addr_of_1149_final_reg_ack_1<= rack(0);
      addr_of_1149_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1149_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1148_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx237_1150,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1302_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1302_final_reg_req_0;
      addr_of_1302_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1302_final_reg_req_1;
      addr_of_1302_final_reg_ack_1<= rack(0);
      addr_of_1302_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1302_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1301_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx337_1303,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1649_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1649_final_reg_req_0;
      addr_of_1649_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1649_final_reg_req_1;
      addr_of_1649_final_reg_ack_1<= rack(0);
      addr_of_1649_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1649_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1648_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx352_1650,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_806_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_806_final_reg_req_0;
      addr_of_806_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_806_final_reg_req_1;
      addr_of_806_final_reg_ack_1<= rack(0);
      addr_of_806_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_806_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_805_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_807,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1002_inst
    process(tmp487_999) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := tmp487_999(63 downto 0);
      type_cast_1002_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1007_inst
    process(ASHR_i64_i64_1006_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := ASHR_i64_i64_1006_wire(63 downto 0);
      phitmp_1008 <= tmp_var; -- 
    end process;
    type_cast_1014_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1014_inst_req_0;
      type_cast_1014_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1014_inst_req_1;
      type_cast_1014_inst_ack_1<= rack(0);
      type_cast_1014_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1014_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => phitmp_1008,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1014_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1058_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1058_inst_req_0;
      type_cast_1058_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1058_inst_req_1;
      type_cast_1058_inst_ack_1<= rack(0);
      type_cast_1058_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1058_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_82_1078,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1058_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1065_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1065_inst_req_0;
      type_cast_1065_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1065_inst_req_1;
      type_cast_1065_inst_ack_1<= rack(0);
      type_cast_1065_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1065_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shl11x_xi_1099,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1065_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1087_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1087_inst_req_0;
      type_cast_1087_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1087_inst_req_1;
      type_cast_1087_inst_ack_1<= rack(0);
      type_cast_1087_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1087_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => callx_xi_1081,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv8x_xi_1088,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1102_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1102_inst_req_0;
      type_cast_1102_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1102_inst_req_1;
      type_cast_1102_inst_ack_1<= rack(0);
      type_cast_1102_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1102_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp_1072,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => convx_xi_1103,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1119_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1119_inst_req_0;
      type_cast_1119_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1119_inst_req_1;
      type_cast_1119_inst_ack_1<= rack(0);
      type_cast_1119_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1119_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shl11x_xi_1099,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1119_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1159_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1159_inst_req_0;
      type_cast_1159_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1159_inst_req_1;
      type_cast_1159_inst_ack_1<= rack(0);
      type_cast_1159_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1159_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add45_529,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv239_1160,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1163_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1163_inst_req_0;
      type_cast_1163_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1163_inst_req_1;
      type_cast_1163_inst_ack_1<= rack(0);
      type_cast_1163_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1163_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add135_684,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv241_1164,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1167_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1167_inst_req_0;
      type_cast_1167_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1167_inst_req_1;
      type_cast_1167_inst_ack_1<= rack(0);
      type_cast_1167_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1167_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add117_653,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv244_1168,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1171_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1171_inst_req_0;
      type_cast_1171_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1171_inst_req_1;
      type_cast_1171_inst_ack_1<= rack(0);
      type_cast_1171_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1171_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add99_622,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv247_1172,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1196_inst
    process(sext_1193) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := sext_1193(63 downto 0);
      type_cast_1196_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1201_inst
    process(ASHR_i64_i64_1200_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := ASHR_i64_i64_1200_wire(63 downto 0);
      conv249_1202 <= tmp_var; -- 
    end process;
    type_cast_1230_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1230_inst_req_0;
      type_cast_1230_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1230_inst_req_1;
      type_cast_1230_inst_ack_1<= rack(0);
      type_cast_1230_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1230_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add99_622,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp12_1231,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1234_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1234_inst_req_0;
      type_cast_1234_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1234_inst_req_1;
      type_cast_1234_inst_ack_1<= rack(0);
      type_cast_1234_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1234_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add45_529,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp13_1235,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1243_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1243_inst_req_0;
      type_cast_1243_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1243_inst_req_1;
      type_cast_1243_inst_ack_1<= rack(0);
      type_cast_1243_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1243_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add117_653,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp15_1244,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1252_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1252_inst_req_0;
      type_cast_1252_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1252_inst_req_1;
      type_cast_1252_inst_ack_1<= rack(0);
      type_cast_1252_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1252_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add135_684,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp17_1253,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1261_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1261_inst_req_0;
      type_cast_1261_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1261_inst_req_1;
      type_cast_1261_inst_ack_1<= rack(0);
      type_cast_1261_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1261_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp18_1258,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp19_1262,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1266_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1266_inst_req_0;
      type_cast_1266_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1266_inst_req_1;
      type_cast_1266_inst_ack_1<= rack(0);
      type_cast_1266_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1266_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1265_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp20_1267,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1295_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1295_inst_req_0;
      type_cast_1295_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1295_inst_req_1;
      type_cast_1295_inst_ack_1<= rack(0);
      type_cast_1295_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1295_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext477_1470,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1295_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1312_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1312_inst_req_0;
      type_cast_1312_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1312_inst_req_1;
      type_cast_1312_inst_ack_1<= rack(0);
      type_cast_1312_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1312_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call260_1306,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv263_1313,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1328_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1328_inst_req_0;
      type_cast_1328_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1328_inst_req_1;
      type_cast_1328_inst_ack_1<= rack(0);
      type_cast_1328_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1328_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call268_1322,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv272_1329,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1349_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1349_inst_req_0;
      type_cast_1349_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1349_inst_req_1;
      type_cast_1349_inst_ack_1<= rack(0);
      type_cast_1349_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1349_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call278_1343,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv282_1350,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1370_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1370_inst_req_0;
      type_cast_1370_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1370_inst_req_1;
      type_cast_1370_inst_ack_1<= rack(0);
      type_cast_1370_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1370_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call288_1364,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv292_1371,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1391_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1391_inst_req_0;
      type_cast_1391_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1391_inst_req_1;
      type_cast_1391_inst_ack_1<= rack(0);
      type_cast_1391_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1391_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call298_1385,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv302_1392,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1412_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1412_inst_req_0;
      type_cast_1412_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1412_inst_req_1;
      type_cast_1412_inst_ack_1<= rack(0);
      type_cast_1412_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1412_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call308_1406,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv312_1413,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1433_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1433_inst_req_0;
      type_cast_1433_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1433_inst_req_1;
      type_cast_1433_inst_ack_1<= rack(0);
      type_cast_1433_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1433_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call318_1427,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv322_1434,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1454_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1454_inst_req_0;
      type_cast_1454_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1454_inst_req_1;
      type_cast_1454_inst_ack_1<= rack(0);
      type_cast_1454_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1454_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call328_1448,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv332_1455,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1498_inst
    process(tmp473_1495) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := tmp473_1495(63 downto 0);
      type_cast_1498_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1503_inst
    process(ASHR_i64_i64_1502_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := ASHR_i64_i64_1502_wire(63 downto 0);
      phitmp451_1504 <= tmp_var; -- 
    end process;
    type_cast_1510_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1510_inst_req_0;
      type_cast_1510_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1510_inst_req_1;
      type_cast_1510_inst_ack_1<= rack(0);
      type_cast_1510_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1510_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => phitmp451_1504,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1510_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1542_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1542_inst_req_0;
      type_cast_1542_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1542_inst_req_1;
      type_cast_1542_inst_ack_1<= rack(0);
      type_cast_1542_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1542_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_120_1539,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv2x_xi418_1543,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1558_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1558_inst_req_0;
      type_cast_1558_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1558_inst_req_1;
      type_cast_1558_inst_ack_1<= rack(0);
      type_cast_1558_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1558_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_128_1578,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1558_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1565_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1565_inst_req_0;
      type_cast_1565_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1565_inst_req_1;
      type_cast_1565_inst_ack_1<= rack(0);
      type_cast_1565_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1565_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shl11x_xi426_1599,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1565_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1587_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1587_inst_req_0;
      type_cast_1587_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1587_inst_req_1;
      type_cast_1587_inst_ack_1<= rack(0);
      type_cast_1587_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1587_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => callx_xi423_1581,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv8x_xi424_1588,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1602_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1602_inst_req_0;
      type_cast_1602_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1602_inst_req_1;
      type_cast_1602_inst_ack_1<= rack(0);
      type_cast_1602_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1602_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp452_1572,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => convx_xi427_1603,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1619_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1619_inst_req_0;
      type_cast_1619_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1619_inst_req_1;
      type_cast_1619_inst_ack_1<= rack(0);
      type_cast_1619_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1619_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shl11x_xi426_1599,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1619_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1698_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1698_inst_req_0;
      type_cast_1698_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1698_inst_req_1;
      type_cast_1698_inst_ack_1<= rack(0);
      type_cast_1698_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1698_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp453_1695,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp3_1699,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1708_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1708_inst_req_0;
      type_cast_1708_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1708_inst_req_1;
      type_cast_1708_inst_ack_1<= rack(0);
      type_cast_1708_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1708_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add117_653,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp6_1709,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1717_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1717_inst_req_0;
      type_cast_1717_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1717_inst_req_1;
      type_cast_1717_inst_ack_1<= rack(0);
      type_cast_1717_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1717_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp7_1714,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp8_1718,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1729_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1729_inst_req_0;
      type_cast_1729_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1729_inst_req_1;
      type_cast_1729_inst_ack_1<= rack(0);
      type_cast_1729_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1729_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1767,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1729_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1746_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1746_inst_req_0;
      type_cast_1746_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1746_inst_req_1;
      type_cast_1746_inst_ack_1<= rack(0);
      type_cast_1746_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1746_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => mul380_1738,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv381_1747,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1750_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1750_inst_req_0;
      type_cast_1750_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1750_inst_req_1;
      type_cast_1750_inst_ack_1<= rack(0);
      type_cast_1750_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1750_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => mul386_1743,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv387_1751,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1783_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1783_inst_req_0;
      type_cast_1783_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1783_inst_req_1;
      type_cast_1783_inst_ack_1<= rack(0);
      type_cast_1783_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1783_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1782_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv356_1784,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1791_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1791_inst_req_0;
      type_cast_1791_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1791_inst_req_1;
      type_cast_1791_inst_ack_1<= rack(0);
      type_cast_1791_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1791_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1790_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv411_1792,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_445_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_445_inst_req_0;
      type_cast_445_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_445_inst_req_1;
      type_cast_445_inst_ack_1<= rack(0);
      type_cast_445_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_445_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_439,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv3_446,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_461_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_461_inst_req_0;
      type_cast_461_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_461_inst_req_1;
      type_cast_461_inst_ack_1<= rack(0);
      type_cast_461_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_461_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call6_455,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv9_462,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_476_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_476_inst_req_0;
      type_cast_476_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_476_inst_req_1;
      type_cast_476_inst_ack_1<= rack(0);
      type_cast_476_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_476_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call14_470,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv19_477,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_492_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_492_inst_req_0;
      type_cast_492_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_492_inst_req_1;
      type_cast_492_inst_ack_1<= rack(0);
      type_cast_492_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_492_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call23_486,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv26_493,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_507_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_507_inst_req_0;
      type_cast_507_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_507_inst_req_1;
      type_cast_507_inst_ack_1<= rack(0);
      type_cast_507_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_507_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call32_501,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv37_508,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_523_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_523_inst_req_0;
      type_cast_523_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_523_inst_req_1;
      type_cast_523_inst_ack_1<= rack(0);
      type_cast_523_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_523_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call41_517,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv44_524,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_538_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_538_inst_req_0;
      type_cast_538_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_538_inst_req_1;
      type_cast_538_inst_ack_1<= rack(0);
      type_cast_538_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_538_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call50_532,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv55_539,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_554_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_554_inst_req_0;
      type_cast_554_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_554_inst_req_1;
      type_cast_554_inst_ack_1<= rack(0);
      type_cast_554_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_554_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call59_548,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv62_555,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_569_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_569_inst_req_0;
      type_cast_569_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_569_inst_req_1;
      type_cast_569_inst_ack_1<= rack(0);
      type_cast_569_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_569_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call68_563,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv73_570,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_585_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_585_inst_req_0;
      type_cast_585_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_585_inst_req_1;
      type_cast_585_inst_ack_1<= rack(0);
      type_cast_585_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_585_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call77_579,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv80_586,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_600_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_600_inst_req_0;
      type_cast_600_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_600_inst_req_1;
      type_cast_600_inst_ack_1<= rack(0);
      type_cast_600_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_600_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call86_594,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv91_601,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_616_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_616_inst_req_0;
      type_cast_616_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_616_inst_req_1;
      type_cast_616_inst_ack_1<= rack(0);
      type_cast_616_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_616_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call95_610,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv98_617,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_631_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_631_inst_req_0;
      type_cast_631_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_631_inst_req_1;
      type_cast_631_inst_ack_1<= rack(0);
      type_cast_631_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_631_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call104_625,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv109_632,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_647_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_647_inst_req_0;
      type_cast_647_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_647_inst_req_1;
      type_cast_647_inst_ack_1<= rack(0);
      type_cast_647_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_647_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call113_641,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv116_648,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_662_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_662_inst_req_0;
      type_cast_662_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_662_inst_req_1;
      type_cast_662_inst_ack_1<= rack(0);
      type_cast_662_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_662_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call122_656,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv127_663,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_678_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_678_inst_req_0;
      type_cast_678_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_678_inst_req_1;
      type_cast_678_inst_ack_1<= rack(0);
      type_cast_678_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_678_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call131_672,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv134_679,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_687_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_687_inst_req_0;
      type_cast_687_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_687_inst_req_1;
      type_cast_687_inst_ack_1<= rack(0);
      type_cast_687_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_687_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add27_498,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv141_688,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_691_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_691_inst_req_0;
      type_cast_691_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_691_inst_req_1;
      type_cast_691_inst_ack_1<= rack(0);
      type_cast_691_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_691_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add45_529,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv143_692,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_707_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_707_inst_req_0;
      type_cast_707_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_707_inst_req_1;
      type_cast_707_inst_ack_1<= rack(0);
      type_cast_707_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_707_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_706_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv145_708,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_735_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_735_inst_req_0;
      type_cast_735_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_735_inst_req_1;
      type_cast_735_inst_ack_1<= rack(0);
      type_cast_735_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_735_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_734_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp483_736,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_751_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_751_inst_req_0;
      type_cast_751_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_751_inst_req_1;
      type_cast_751_inst_ack_1<= rack(0);
      type_cast_751_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_751_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add27_498,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp24_752,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_760_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_760_inst_req_0;
      type_cast_760_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_760_inst_req_1;
      type_cast_760_inst_ack_1<= rack(0);
      type_cast_760_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_760_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add45_529,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp26_761,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_770_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_770_inst_req_0;
      type_cast_770_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_770_inst_req_1;
      type_cast_770_inst_ack_1<= rack(0);
      type_cast_770_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_770_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_769_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp28_771,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_799_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_799_inst_req_0;
      type_cast_799_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_799_inst_req_1;
      type_cast_799_inst_ack_1<= rack(0);
      type_cast_799_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_799_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext491_974,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_799_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_816_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_816_inst_req_0;
      type_cast_816_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_816_inst_req_1;
      type_cast_816_inst_ack_1<= rack(0);
      type_cast_816_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_816_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call153_810,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv156_817,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_832_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_832_inst_req_0;
      type_cast_832_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_832_inst_req_1;
      type_cast_832_inst_ack_1<= rack(0);
      type_cast_832_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_832_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call161_826,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv165_833,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_853_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_853_inst_req_0;
      type_cast_853_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_853_inst_req_1;
      type_cast_853_inst_ack_1<= rack(0);
      type_cast_853_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_853_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call171_847,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv175_854,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_874_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_874_inst_req_0;
      type_cast_874_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_874_inst_req_1;
      type_cast_874_inst_ack_1<= rack(0);
      type_cast_874_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_874_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call181_868,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv185_875,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_895_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_895_inst_req_0;
      type_cast_895_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_895_inst_req_1;
      type_cast_895_inst_ack_1<= rack(0);
      type_cast_895_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_895_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call191_889,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv195_896,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_916_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_916_inst_req_0;
      type_cast_916_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_916_inst_req_1;
      type_cast_916_inst_ack_1<= rack(0);
      type_cast_916_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_916_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call201_910,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv205_917,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_937_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_937_inst_req_0;
      type_cast_937_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_937_inst_req_1;
      type_cast_937_inst_ack_1<= rack(0);
      type_cast_937_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_937_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call211_931,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv215_938,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_958_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_958_inst_req_0;
      type_cast_958_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_958_inst_req_1;
      type_cast_958_inst_ack_1<= rack(0);
      type_cast_958_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_958_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call221_952,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv225_959,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1148_index_1_rename
    process(R_ix_x0x_xlcssa_1147_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_ix_x0x_xlcssa_1147_resized;
      ov(13 downto 0) := iv;
      R_ix_x0x_xlcssa_1147_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1148_index_1_resize
    process(ix_x0x_xlcssa_1011) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ix_x0x_xlcssa_1011;
      ov := iv(13 downto 0);
      R_ix_x0x_xlcssa_1147_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1148_root_address_inst
    process(array_obj_ref_1148_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1148_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1148_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1301_index_1_rename
    process(R_indvar476_1300_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar476_1300_resized;
      ov(13 downto 0) := iv;
      R_indvar476_1300_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1301_index_1_resize
    process(indvar476_1289) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar476_1289;
      ov := iv(13 downto 0);
      R_indvar476_1300_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1301_root_address_inst
    process(array_obj_ref_1301_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1301_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1301_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1648_index_1_rename
    process(R_ix_x1x_xlcssa_1647_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_ix_x1x_xlcssa_1647_resized;
      ov(13 downto 0) := iv;
      R_ix_x1x_xlcssa_1647_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1648_index_1_resize
    process(ix_x1x_xlcssa_1507) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ix_x1x_xlcssa_1507;
      ov := iv(13 downto 0);
      R_ix_x1x_xlcssa_1647_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1648_root_address_inst
    process(array_obj_ref_1648_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1648_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1648_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_805_index_1_rename
    process(R_indvar490_804_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar490_804_resized;
      ov(13 downto 0) := iv;
      R_indvar490_804_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_805_index_1_resize
    process(indvar490_793) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar490_793;
      ov := iv(13 downto 0);
      R_indvar490_804_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_805_root_address_inst
    process(array_obj_ref_805_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_805_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_805_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1152_addr_0
    process(ptr_deref_1152_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1152_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1152_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1152_base_resize
    process(arrayidx237_1150) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx237_1150;
      ov := iv(13 downto 0);
      ptr_deref_1152_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1152_gather_scatter
    process(shl17x_xi_1143) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := shl17x_xi_1143;
      ov(63 downto 0) := iv;
      ptr_deref_1152_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1152_root_address_inst
    process(ptr_deref_1152_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1152_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1152_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1462_addr_0
    process(ptr_deref_1462_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1462_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1462_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1462_base_resize
    process(arrayidx337_1303) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx337_1303;
      ov := iv(13 downto 0);
      ptr_deref_1462_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1462_gather_scatter
    process(add333_1460) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add333_1460;
      ov(63 downto 0) := iv;
      ptr_deref_1462_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1462_root_address_inst
    process(ptr_deref_1462_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1462_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1462_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1652_addr_0
    process(ptr_deref_1652_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1652_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1652_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1652_base_resize
    process(arrayidx352_1650) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx352_1650;
      ov := iv(13 downto 0);
      ptr_deref_1652_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1652_gather_scatter
    process(shl17x_xi436_1643) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := shl17x_xi436_1643;
      ov(63 downto 0) := iv;
      ptr_deref_1652_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1652_root_address_inst
    process(ptr_deref_1652_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1652_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1652_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_966_addr_0
    process(ptr_deref_966_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_966_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_966_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_966_base_resize
    process(arrayidx_807) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_807;
      ov := iv(13 downto 0);
      ptr_deref_966_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_966_gather_scatter
    process(add226_964) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add226_964;
      ov(63 downto 0) := iv;
      ptr_deref_966_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_966_root_address_inst
    process(ptr_deref_966_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_966_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_966_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1031_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tobool_1030;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1031_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1031_branch_req_0,
          ack0 => if_stmt_1031_branch_ack_0,
          ack1 => if_stmt_1031_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1109_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmpx_xi_1108;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1109_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1109_branch_req_0,
          ack0 => if_stmt_1109_branch_ack_0,
          ack1 => if_stmt_1109_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1209_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp255443_1208;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1209_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1209_branch_req_0,
          ack0 => if_stmt_1209_branch_ack_0,
          ack1 => if_stmt_1209_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1476_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond_1475;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1476_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1476_branch_req_0,
          ack0 => if_stmt_1476_branch_ack_0,
          ack1 => if_stmt_1476_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1527_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tobool344_1526;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1527_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1527_branch_req_0,
          ack0 => if_stmt_1527_branch_ack_0,
          ack1 => if_stmt_1527_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1609_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmpx_xi428_1608;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1609_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1609_branch_req_0,
          ack0 => if_stmt_1609_branch_ack_0,
          ack1 => if_stmt_1609_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1773_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond5_1772;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1773_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1773_branch_req_0,
          ack0 => if_stmt_1773_branch_ack_0,
          ack1 => if_stmt_1773_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_715_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp447_714;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_715_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_715_branch_req_0,
          ack0 => if_stmt_715_branch_ack_0,
          ack1 => if_stmt_715_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_980_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond32_979;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_980_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_980_branch_req_0,
          ack0 => if_stmt_980_branch_ack_0,
          ack1 => if_stmt_980_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1071_inst
    process(nx_x025x_xi_1052) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(nx_x025x_xi_1052, type_cast_1070_wire_constant, tmp_var);
      tmp_1072 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1077_inst
    process(nx_x025x_xi_1052) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(nx_x025x_xi_1052, type_cast_1076_wire_constant, tmp_var);
      iNsTr_82_1078 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1571_inst
    process(nx_x025x_xi421_1552) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(nx_x025x_xi421_1552, type_cast_1570_wire_constant, tmp_var);
      tmp452_1572 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1577_inst
    process(nx_x025x_xi421_1552) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(nx_x025x_xi421_1552, type_cast_1576_wire_constant, tmp_var);
      iNsTr_128_1578 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1682_inst
    process(add81_591) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add81_591, type_cast_1681_wire_constant, tmp_var);
      sub_1683 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1688_inst
    process(add117_653) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add117_653, type_cast_1687_wire_constant, tmp_var);
      sub395_1689 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1694_inst
    process(add99_622) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add99_622, type_cast_1693_wire_constant, tmp_var);
      tmp453_1695 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1704_inst
    process(tmp3_1699) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp3_1699, type_cast_1703_wire_constant, tmp_var);
      tmp4_1705 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1742_inst
    process(tmp9_1723, mul380_1738) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp9_1723, mul380_1738, tmp_var);
      mul386_1743 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1766_inst
    process(indvar_1726) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1726, type_cast_1765_wire_constant, tmp_var);
      indvarx_xnext_1767 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1469_inst
    process(indvar476_1289) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar476_1289, type_cast_1468_wire_constant, tmp_var);
      indvarx_xnext477_1470 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_973_inst
    process(indvar490_793) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar490_793, type_cast_972_wire_constant, tmp_var);
      indvarx_xnext491_974 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_1048_inst
    process(conv2x_xi_1043) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv2x_xi_1043, type_cast_1047_wire_constant, tmp_var);
      shlx_xi_1049 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_1548_inst
    process(conv2x_xi418_1543) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv2x_xi418_1543, type_cast_1547_wire_constant, tmp_var);
      shlx_xi419_1549 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_1023_inst
    process(conv145_708) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv145_708, type_cast_1022_wire_constant, tmp_var);
      and_1024 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_1131_inst
    process(Bx_xnot_1126) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(Bx_xnot_1126, type_cast_1130_wire_constant, tmp_var);
      add1519x_xi_1132 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_1519_inst
    process(conv249_1202) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv249_1202, type_cast_1518_wire_constant, tmp_var);
      and343_1520 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_1631_inst
    process(iNsTr_138_1626) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(iNsTr_138_1626, type_cast_1630_wire_constant, tmp_var);
      add1519x_xi434_1632 <= tmp_var; --
    end process;
    -- binary operator ASHR_i64_i64_1006_inst
    process(type_cast_1002_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1002_wire, type_cast_1005_wire_constant, tmp_var);
      ASHR_i64_i64_1006_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i64_i64_1200_inst
    process(type_cast_1196_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1196_wire, type_cast_1199_wire_constant, tmp_var);
      ASHR_i64_i64_1200_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i64_i64_1502_inst
    process(type_cast_1498_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1498_wire, type_cast_1501_wire_constant, tmp_var);
      ASHR_i64_i64_1502_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1771_inst
    process(indvarx_xnext_1767, tmp4_1705) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_1767, tmp4_1705, tmp_var);
      exitcond5_1772 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1029_inst
    process(and_1024) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(and_1024, type_cast_1028_wire_constant, tmp_var);
      tobool_1030 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1474_inst
    process(indvarx_xnext477_1470, umax23_1286) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext477_1470, umax23_1286, tmp_var);
      exitcond_1475 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1525_inst
    process(and343_1520) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(and343_1520, type_cast_1524_wire_constant, tmp_var);
      tobool344_1526 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_978_inst
    process(indvarx_xnext491_974, umax31_790) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext491_974, umax31_790, tmp_var);
      exitcond32_979 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1220_inst
    process(conv249_1202) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv249_1202, type_cast_1219_wire_constant, tmp_var);
      tmp471_1221 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1272_inst
    process(tmp20_1267) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp20_1267, type_cast_1271_wire_constant, tmp_var);
      tmp21_1273 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_741_inst
    process(tmp483_736) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp483_736, type_cast_740_wire_constant, tmp_var);
      tmp484_742 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_776_inst
    process(tmp28_771) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp28_771, type_cast_775_wire_constant, tmp_var);
      tmp29_777 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1664_inst
    process(add135_684, add45_529) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(add135_684, add45_529, tmp_var);
      mul362_1665 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1669_inst
    process(add81_591, add63_560) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(add81_591, add63_560, tmp_var);
      mul375_1670 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1713_inst
    process(add135_684, add45_529) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(add135_684, add45_529, tmp_var);
      tmp7_1714 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1722_inst
    process(tmp6_1709, tmp8_1718) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp6_1709, tmp8_1718, tmp_var);
      tmp9_1723 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1737_inst
    process(tmp9_1723, indvar_1726) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp9_1723, indvar_1726, tmp_var);
      mul380_1738 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_696_inst
    process(conv141_688, add_467) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv141_688, add_467, tmp_var);
      mul_697 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_701_inst
    process(mul_697, conv143_692) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_697, conv143_692, tmp_var);
      mul144_702 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_725_inst
    process(add_467, conv141_688) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add_467, conv141_688, tmp_var);
      tmp480_726 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_730_inst
    process(tmp480_726, conv143_692) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp480_726, conv143_692, tmp_var);
      tmp482_731 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_756_inst
    process(add_467, tmp24_752) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add_467, tmp24_752, tmp_var);
      tmp25_757 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_765_inst
    process(tmp25_757, tmp26_761) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp25_757, tmp26_761, tmp_var);
      tmp27_766 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1176_inst
    process(conv247_1172, conv239_1160) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv247_1172, conv239_1160, tmp_var);
      mul242_1177 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1181_inst
    process(mul242_1177, conv244_1168) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul242_1177, conv244_1168, tmp_var);
      mul245_1182 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1186_inst
    process(mul245_1182, conv241_1164) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul245_1182, conv241_1164, tmp_var);
      mul248_1187 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1239_inst
    process(tmp12_1231, tmp13_1235) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp12_1231, tmp13_1235, tmp_var);
      tmp14_1240 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1248_inst
    process(tmp14_1240, tmp15_1244) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp14_1240, tmp15_1244, tmp_var);
      tmp16_1249 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1257_inst
    process(tmp16_1249, tmp17_1253) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp16_1249, tmp17_1253, tmp_var);
      tmp18_1258 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_497_inst
    process(conv26_493, shl20_483) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv26_493, shl20_483, tmp_var);
      add27_498 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_528_inst
    process(conv44_524, shl38_514) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv44_524, shl38_514, tmp_var);
      add45_529 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_559_inst
    process(conv62_555, shl56_545) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv62_555, shl56_545, tmp_var);
      add63_560 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_590_inst
    process(conv80_586, shl74_576) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv80_586, shl74_576, tmp_var);
      add81_591 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_621_inst
    process(conv98_617, shl92_607) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv98_617, shl92_607, tmp_var);
      add99_622 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_652_inst
    process(conv116_648, shl110_638) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv116_648, shl110_638, tmp_var);
      add117_653 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_683_inst
    process(conv134_679, shl128_669) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv134_679, shl128_669, tmp_var);
      add135_684 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_466_inst
    process(conv9_462, shl_452) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv9_462, shl_452, tmp_var);
      add_467 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1092_inst
    process(conv8x_xi_1088, elementx_x024x_xi_1059) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv8x_xi_1088, elementx_x024x_xi_1059, tmp_var);
      addx_xi_1093 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1333_inst
    process(conv272_1329, shl265_1319) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv272_1329, shl265_1319, tmp_var);
      add273_1334 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1354_inst
    process(shl275_1340, conv282_1350) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl275_1340, conv282_1350, tmp_var);
      add283_1355 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1375_inst
    process(shl285_1361, conv292_1371) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl285_1361, conv292_1371, tmp_var);
      add293_1376 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1396_inst
    process(shl295_1382, conv302_1392) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl295_1382, conv302_1392, tmp_var);
      add303_1397 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1417_inst
    process(shl305_1403, conv312_1413) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl305_1403, conv312_1413, tmp_var);
      add313_1418 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1438_inst
    process(shl315_1424, conv322_1434) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl315_1424, conv322_1434, tmp_var);
      add323_1439 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1459_inst
    process(shl325_1445, conv332_1455) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl325_1445, conv332_1455, tmp_var);
      add333_1460 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1592_inst
    process(conv8x_xi424_1588, elementx_x024x_xi422_1559) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv8x_xi424_1588, elementx_x024x_xi422_1559, tmp_var);
      addx_xi425_1593 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_837_inst
    process(conv165_833, shl158_823) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv165_833, shl158_823, tmp_var);
      add166_838 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_858_inst
    process(shl168_844, conv175_854) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl168_844, conv175_854, tmp_var);
      add176_859 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_879_inst
    process(shl178_865, conv185_875) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl178_865, conv185_875, tmp_var);
      add186_880 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_900_inst
    process(shl188_886, conv195_896) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl188_886, conv195_896, tmp_var);
      add196_901 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_921_inst
    process(shl198_907, conv205_917) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl198_907, conv205_917, tmp_var);
      add206_922 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_942_inst
    process(shl208_928, conv215_938) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl208_928, conv215_938, tmp_var);
      add216_943 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_963_inst
    process(shl218_949, conv225_959) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl218_949, conv225_959, tmp_var);
      add226_964 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_482_inst
    process(conv19_477) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv19_477, type_cast_481_wire_constant, tmp_var);
      shl20_483 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_513_inst
    process(conv37_508) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv37_508, type_cast_512_wire_constant, tmp_var);
      shl38_514 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_544_inst
    process(conv55_539) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv55_539, type_cast_543_wire_constant, tmp_var);
      shl56_545 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_575_inst
    process(conv73_570) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv73_570, type_cast_574_wire_constant, tmp_var);
      shl74_576 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_606_inst
    process(conv91_601) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv91_601, type_cast_605_wire_constant, tmp_var);
      shl92_607 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_637_inst
    process(conv109_632) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv109_632, type_cast_636_wire_constant, tmp_var);
      shl110_638 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_668_inst
    process(conv127_663) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv127_663, type_cast_667_wire_constant, tmp_var);
      shl128_669 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1042_inst
    process(mul144_702) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul144_702, type_cast_1041_wire_constant, tmp_var);
      conv2x_xi_1043 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_451_inst
    process(conv3_446) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv3_446, type_cast_450_wire_constant, tmp_var);
      shl_452 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1098_inst
    process(addx_xi_1093) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(addx_xi_1093, type_cast_1097_wire_constant, tmp_var);
      shl11x_xi_1099 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1125_inst
    process(conv145_708) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv145_708, type_cast_1124_wire_constant, tmp_var);
      Bx_xnot_1126 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1142_inst
    process(shl11x_xix_xlcssa_1116, sh_promx_xi_1138) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(shl11x_xix_xlcssa_1116, sh_promx_xi_1138, tmp_var);
      shl17x_xi_1143 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1192_inst
    process(mul248_1187) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul248_1187, type_cast_1191_wire_constant, tmp_var);
      sext_1193 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1318_inst
    process(conv263_1313) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv263_1313, type_cast_1317_wire_constant, tmp_var);
      shl265_1319 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1339_inst
    process(add273_1334) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add273_1334, type_cast_1338_wire_constant, tmp_var);
      shl275_1340 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1360_inst
    process(add283_1355) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add283_1355, type_cast_1359_wire_constant, tmp_var);
      shl285_1361 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1381_inst
    process(add293_1376) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add293_1376, type_cast_1380_wire_constant, tmp_var);
      shl295_1382 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1402_inst
    process(add303_1397) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add303_1397, type_cast_1401_wire_constant, tmp_var);
      shl305_1403 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1423_inst
    process(add313_1418) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add313_1418, type_cast_1422_wire_constant, tmp_var);
      shl315_1424 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1444_inst
    process(add323_1439) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add323_1439, type_cast_1443_wire_constant, tmp_var);
      shl325_1445 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1494_inst
    process(umax_1489) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(umax_1489, type_cast_1493_wire_constant, tmp_var);
      tmp473_1495 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1538_inst
    process(mul248_1187) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul248_1187, type_cast_1537_wire_constant, tmp_var);
      iNsTr_120_1539 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1598_inst
    process(addx_xi425_1593) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(addx_xi425_1593, type_cast_1597_wire_constant, tmp_var);
      shl11x_xi426_1599 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1625_inst
    process(mul248_1187) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul248_1187, type_cast_1624_wire_constant, tmp_var);
      iNsTr_138_1626 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1642_inst
    process(shl11x_xi426x_xlcssa_1616, sh_promx_xi435_1638) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(shl11x_xi426x_xlcssa_1616, sh_promx_xi435_1638, tmp_var);
      shl17x_xi436_1643 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_822_inst
    process(conv156_817) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv156_817, type_cast_821_wire_constant, tmp_var);
      shl158_823 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_843_inst
    process(add166_838) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add166_838, type_cast_842_wire_constant, tmp_var);
      shl168_844 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_864_inst
    process(add176_859) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add176_859, type_cast_863_wire_constant, tmp_var);
      shl178_865 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_885_inst
    process(add186_880) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add186_880, type_cast_884_wire_constant, tmp_var);
      shl188_886 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_906_inst
    process(add196_901) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add196_901, type_cast_905_wire_constant, tmp_var);
      shl198_907 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_927_inst
    process(add206_922) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add206_922, type_cast_926_wire_constant, tmp_var);
      shl208_928 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_948_inst
    process(add216_943) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add216_943, type_cast_947_wire_constant, tmp_var);
      shl218_949 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_998_inst
    process(umax486_993) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(umax486_993, type_cast_997_wire_constant, tmp_var);
      tmp487_999 <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_1796_inst
    process(conv411_1792, conv356_1784) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv411_1792, conv356_1784, tmp_var);
      sub415_1797 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_713_inst
    process(mul144_702) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul144_702, type_cast_712_wire_constant, tmp_var);
      cmp447_714 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_1207_inst
    process(conv249_1202) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(conv249_1202, type_cast_1206_wire_constant, tmp_var);
      cmp255443_1208 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_1226_inst
    process(tmp471_1221) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp471_1221, type_cast_1225_wire_constant, tmp_var);
      tmp472_1227 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_1278_inst
    process(tmp21_1273) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp21_1273, type_cast_1277_wire_constant, tmp_var);
      tmp22_1279 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_747_inst
    process(tmp484_742) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp484_742, type_cast_746_wire_constant, tmp_var);
      tmp485_748 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_782_inst
    process(tmp29_777) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp29_777, type_cast_781_wire_constant, tmp_var);
      tmp30_783 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_1107_inst
    process(convx_xi_1103, shlx_xi_1049) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(convx_xi_1103, shlx_xi_1049, tmp_var);
      cmpx_xi_1108 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_1607_inst
    process(convx_xi427_1603, shlx_xi419_1549) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(convx_xi427_1603, shlx_xi419_1549, tmp_var);
      cmpx_xi428_1608 <= tmp_var; --
    end process;
    -- binary operator XOR_u64_u64_1137_inst
    process(add1519x_xi_1132) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntXor_proc(add1519x_xi_1132, type_cast_1136_wire_constant, tmp_var);
      sh_promx_xi_1138 <= tmp_var; --
    end process;
    -- binary operator XOR_u64_u64_1637_inst
    process(add1519x_xi434_1632) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntXor_proc(add1519x_xi434_1632, type_cast_1636_wire_constant, tmp_var);
      sh_promx_xi435_1638 <= tmp_var; --
    end process;
    -- shared split operator group (115) : array_obj_ref_1148_index_offset 
    ApIntAdd_group_115: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_ix_x0x_xlcssa_1147_scaled;
      array_obj_ref_1148_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1148_index_offset_req_0;
      array_obj_ref_1148_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1148_index_offset_req_1;
      array_obj_ref_1148_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_115_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_115_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_115",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 115
    -- shared split operator group (116) : array_obj_ref_1301_index_offset 
    ApIntAdd_group_116: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar476_1300_scaled;
      array_obj_ref_1301_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1301_index_offset_req_0;
      array_obj_ref_1301_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1301_index_offset_req_1;
      array_obj_ref_1301_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_116_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_116_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_116",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 116
    -- shared split operator group (117) : array_obj_ref_1648_index_offset 
    ApIntAdd_group_117: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_ix_x1x_xlcssa_1647_scaled;
      array_obj_ref_1648_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1648_index_offset_req_0;
      array_obj_ref_1648_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1648_index_offset_req_1;
      array_obj_ref_1648_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_117_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_117_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_117",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 117
    -- shared split operator group (118) : array_obj_ref_805_index_offset 
    ApIntAdd_group_118: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar490_804_scaled;
      array_obj_ref_805_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_805_index_offset_req_0;
      array_obj_ref_805_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_805_index_offset_req_1;
      array_obj_ref_805_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_118_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_118_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_118",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 118
    -- unary operator type_cast_1265_inst
    process(tmp19_1262) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", tmp19_1262, tmp_var);
      type_cast_1265_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1782_inst
    process(call355_1659) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call355_1659, tmp_var);
      type_cast_1782_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1790_inst
    process(call410_1787) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call410_1787, tmp_var);
      type_cast_1790_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_706_inst
    process(mul144_702) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", mul144_702, tmp_var);
      type_cast_706_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_734_inst
    process(tmp482_731) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", tmp482_731, tmp_var);
      type_cast_734_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_769_inst
    process(tmp27_766) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", tmp27_766, tmp_var);
      type_cast_769_wire <= tmp_var; -- 
    end process;
    -- shared store operator group (0) : ptr_deref_1152_store_0 ptr_deref_966_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(27 downto 0);
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1152_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_966_store_0_req_0;
      ptr_deref_1152_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_966_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1152_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_966_store_0_req_1;
      ptr_deref_1152_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_966_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup0_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1152_word_address_0 & ptr_deref_966_word_address_0;
      data_in <= ptr_deref_1152_data_0 & ptr_deref_966_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(13 downto 0),
          mdata => memory_space_1_sr_data(63 downto 0),
          mtag => memory_space_1_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : ptr_deref_1462_store_0 ptr_deref_1652_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(27 downto 0);
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1462_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1652_store_0_req_0;
      ptr_deref_1462_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1652_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1462_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1652_store_0_req_1;
      ptr_deref_1462_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1652_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup1_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup1_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup1_gI: SplitGuardInterface generic map(name => "StoreGroup1_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1462_word_address_0 & ptr_deref_1652_word_address_0;
      data_in <= ptr_deref_1462_data_0 & ptr_deref_1652_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup1 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(13 downto 0),
          mdata => memory_space_0_sr_data(63 downto 0),
          mtag => memory_space_0_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup1 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared inport operator group (0) : RPIPE_maxpool_input_pipe_1447_inst RPIPE_maxpool_input_pipe_1580_inst RPIPE_maxpool_input_pipe_1080_inst RPIPE_maxpool_input_pipe_1305_inst RPIPE_maxpool_input_pipe_1363_inst RPIPE_maxpool_input_pipe_1384_inst RPIPE_maxpool_input_pipe_1405_inst RPIPE_maxpool_input_pipe_1321_inst RPIPE_maxpool_input_pipe_438_inst RPIPE_maxpool_input_pipe_1426_inst RPIPE_maxpool_input_pipe_1342_inst RPIPE_maxpool_input_pipe_454_inst RPIPE_maxpool_input_pipe_469_inst RPIPE_maxpool_input_pipe_485_inst RPIPE_maxpool_input_pipe_500_inst RPIPE_maxpool_input_pipe_516_inst RPIPE_maxpool_input_pipe_531_inst RPIPE_maxpool_input_pipe_547_inst RPIPE_maxpool_input_pipe_562_inst RPIPE_maxpool_input_pipe_578_inst RPIPE_maxpool_input_pipe_593_inst RPIPE_maxpool_input_pipe_609_inst RPIPE_maxpool_input_pipe_624_inst RPIPE_maxpool_input_pipe_640_inst RPIPE_maxpool_input_pipe_655_inst RPIPE_maxpool_input_pipe_671_inst RPIPE_maxpool_input_pipe_809_inst RPIPE_maxpool_input_pipe_825_inst RPIPE_maxpool_input_pipe_846_inst RPIPE_maxpool_input_pipe_867_inst RPIPE_maxpool_input_pipe_888_inst RPIPE_maxpool_input_pipe_909_inst RPIPE_maxpool_input_pipe_930_inst RPIPE_maxpool_input_pipe_951_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(271 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 33 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 33 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 33 downto 0);
      signal guard_vector : std_logic_vector( 33 downto 0);
      constant outBUFs : IntegerArray(33 downto 0) := (33 => 1, 32 => 1, 31 => 1, 30 => 1, 29 => 1, 28 => 1, 27 => 1, 26 => 1, 25 => 1, 24 => 1, 23 => 1, 22 => 1, 21 => 1, 20 => 1, 19 => 1, 18 => 1, 17 => 1, 16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(33 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false, 17 => false, 18 => false, 19 => false, 20 => false, 21 => false, 22 => false, 23 => false, 24 => false, 25 => false, 26 => false, 27 => false, 28 => false, 29 => false, 30 => false, 31 => false, 32 => false, 33 => false);
      constant guardBuffering: IntegerArray(33 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2, 17 => 2, 18 => 2, 19 => 2, 20 => 2, 21 => 2, 22 => 2, 23 => 2, 24 => 2, 25 => 2, 26 => 2, 27 => 2, 28 => 2, 29 => 2, 30 => 2, 31 => 2, 32 => 2, 33 => 2);
      -- 
    begin -- 
      reqL_unguarded(33) <= RPIPE_maxpool_input_pipe_1447_inst_req_0;
      reqL_unguarded(32) <= RPIPE_maxpool_input_pipe_1580_inst_req_0;
      reqL_unguarded(31) <= RPIPE_maxpool_input_pipe_1080_inst_req_0;
      reqL_unguarded(30) <= RPIPE_maxpool_input_pipe_1305_inst_req_0;
      reqL_unguarded(29) <= RPIPE_maxpool_input_pipe_1363_inst_req_0;
      reqL_unguarded(28) <= RPIPE_maxpool_input_pipe_1384_inst_req_0;
      reqL_unguarded(27) <= RPIPE_maxpool_input_pipe_1405_inst_req_0;
      reqL_unguarded(26) <= RPIPE_maxpool_input_pipe_1321_inst_req_0;
      reqL_unguarded(25) <= RPIPE_maxpool_input_pipe_438_inst_req_0;
      reqL_unguarded(24) <= RPIPE_maxpool_input_pipe_1426_inst_req_0;
      reqL_unguarded(23) <= RPIPE_maxpool_input_pipe_1342_inst_req_0;
      reqL_unguarded(22) <= RPIPE_maxpool_input_pipe_454_inst_req_0;
      reqL_unguarded(21) <= RPIPE_maxpool_input_pipe_469_inst_req_0;
      reqL_unguarded(20) <= RPIPE_maxpool_input_pipe_485_inst_req_0;
      reqL_unguarded(19) <= RPIPE_maxpool_input_pipe_500_inst_req_0;
      reqL_unguarded(18) <= RPIPE_maxpool_input_pipe_516_inst_req_0;
      reqL_unguarded(17) <= RPIPE_maxpool_input_pipe_531_inst_req_0;
      reqL_unguarded(16) <= RPIPE_maxpool_input_pipe_547_inst_req_0;
      reqL_unguarded(15) <= RPIPE_maxpool_input_pipe_562_inst_req_0;
      reqL_unguarded(14) <= RPIPE_maxpool_input_pipe_578_inst_req_0;
      reqL_unguarded(13) <= RPIPE_maxpool_input_pipe_593_inst_req_0;
      reqL_unguarded(12) <= RPIPE_maxpool_input_pipe_609_inst_req_0;
      reqL_unguarded(11) <= RPIPE_maxpool_input_pipe_624_inst_req_0;
      reqL_unguarded(10) <= RPIPE_maxpool_input_pipe_640_inst_req_0;
      reqL_unguarded(9) <= RPIPE_maxpool_input_pipe_655_inst_req_0;
      reqL_unguarded(8) <= RPIPE_maxpool_input_pipe_671_inst_req_0;
      reqL_unguarded(7) <= RPIPE_maxpool_input_pipe_809_inst_req_0;
      reqL_unguarded(6) <= RPIPE_maxpool_input_pipe_825_inst_req_0;
      reqL_unguarded(5) <= RPIPE_maxpool_input_pipe_846_inst_req_0;
      reqL_unguarded(4) <= RPIPE_maxpool_input_pipe_867_inst_req_0;
      reqL_unguarded(3) <= RPIPE_maxpool_input_pipe_888_inst_req_0;
      reqL_unguarded(2) <= RPIPE_maxpool_input_pipe_909_inst_req_0;
      reqL_unguarded(1) <= RPIPE_maxpool_input_pipe_930_inst_req_0;
      reqL_unguarded(0) <= RPIPE_maxpool_input_pipe_951_inst_req_0;
      RPIPE_maxpool_input_pipe_1447_inst_ack_0 <= ackL_unguarded(33);
      RPIPE_maxpool_input_pipe_1580_inst_ack_0 <= ackL_unguarded(32);
      RPIPE_maxpool_input_pipe_1080_inst_ack_0 <= ackL_unguarded(31);
      RPIPE_maxpool_input_pipe_1305_inst_ack_0 <= ackL_unguarded(30);
      RPIPE_maxpool_input_pipe_1363_inst_ack_0 <= ackL_unguarded(29);
      RPIPE_maxpool_input_pipe_1384_inst_ack_0 <= ackL_unguarded(28);
      RPIPE_maxpool_input_pipe_1405_inst_ack_0 <= ackL_unguarded(27);
      RPIPE_maxpool_input_pipe_1321_inst_ack_0 <= ackL_unguarded(26);
      RPIPE_maxpool_input_pipe_438_inst_ack_0 <= ackL_unguarded(25);
      RPIPE_maxpool_input_pipe_1426_inst_ack_0 <= ackL_unguarded(24);
      RPIPE_maxpool_input_pipe_1342_inst_ack_0 <= ackL_unguarded(23);
      RPIPE_maxpool_input_pipe_454_inst_ack_0 <= ackL_unguarded(22);
      RPIPE_maxpool_input_pipe_469_inst_ack_0 <= ackL_unguarded(21);
      RPIPE_maxpool_input_pipe_485_inst_ack_0 <= ackL_unguarded(20);
      RPIPE_maxpool_input_pipe_500_inst_ack_0 <= ackL_unguarded(19);
      RPIPE_maxpool_input_pipe_516_inst_ack_0 <= ackL_unguarded(18);
      RPIPE_maxpool_input_pipe_531_inst_ack_0 <= ackL_unguarded(17);
      RPIPE_maxpool_input_pipe_547_inst_ack_0 <= ackL_unguarded(16);
      RPIPE_maxpool_input_pipe_562_inst_ack_0 <= ackL_unguarded(15);
      RPIPE_maxpool_input_pipe_578_inst_ack_0 <= ackL_unguarded(14);
      RPIPE_maxpool_input_pipe_593_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_maxpool_input_pipe_609_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_maxpool_input_pipe_624_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_maxpool_input_pipe_640_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_maxpool_input_pipe_655_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_maxpool_input_pipe_671_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_maxpool_input_pipe_809_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_maxpool_input_pipe_825_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_maxpool_input_pipe_846_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_maxpool_input_pipe_867_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_maxpool_input_pipe_888_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_maxpool_input_pipe_909_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_maxpool_input_pipe_930_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_maxpool_input_pipe_951_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(33) <= RPIPE_maxpool_input_pipe_1447_inst_req_1;
      reqR_unguarded(32) <= RPIPE_maxpool_input_pipe_1580_inst_req_1;
      reqR_unguarded(31) <= RPIPE_maxpool_input_pipe_1080_inst_req_1;
      reqR_unguarded(30) <= RPIPE_maxpool_input_pipe_1305_inst_req_1;
      reqR_unguarded(29) <= RPIPE_maxpool_input_pipe_1363_inst_req_1;
      reqR_unguarded(28) <= RPIPE_maxpool_input_pipe_1384_inst_req_1;
      reqR_unguarded(27) <= RPIPE_maxpool_input_pipe_1405_inst_req_1;
      reqR_unguarded(26) <= RPIPE_maxpool_input_pipe_1321_inst_req_1;
      reqR_unguarded(25) <= RPIPE_maxpool_input_pipe_438_inst_req_1;
      reqR_unguarded(24) <= RPIPE_maxpool_input_pipe_1426_inst_req_1;
      reqR_unguarded(23) <= RPIPE_maxpool_input_pipe_1342_inst_req_1;
      reqR_unguarded(22) <= RPIPE_maxpool_input_pipe_454_inst_req_1;
      reqR_unguarded(21) <= RPIPE_maxpool_input_pipe_469_inst_req_1;
      reqR_unguarded(20) <= RPIPE_maxpool_input_pipe_485_inst_req_1;
      reqR_unguarded(19) <= RPIPE_maxpool_input_pipe_500_inst_req_1;
      reqR_unguarded(18) <= RPIPE_maxpool_input_pipe_516_inst_req_1;
      reqR_unguarded(17) <= RPIPE_maxpool_input_pipe_531_inst_req_1;
      reqR_unguarded(16) <= RPIPE_maxpool_input_pipe_547_inst_req_1;
      reqR_unguarded(15) <= RPIPE_maxpool_input_pipe_562_inst_req_1;
      reqR_unguarded(14) <= RPIPE_maxpool_input_pipe_578_inst_req_1;
      reqR_unguarded(13) <= RPIPE_maxpool_input_pipe_593_inst_req_1;
      reqR_unguarded(12) <= RPIPE_maxpool_input_pipe_609_inst_req_1;
      reqR_unguarded(11) <= RPIPE_maxpool_input_pipe_624_inst_req_1;
      reqR_unguarded(10) <= RPIPE_maxpool_input_pipe_640_inst_req_1;
      reqR_unguarded(9) <= RPIPE_maxpool_input_pipe_655_inst_req_1;
      reqR_unguarded(8) <= RPIPE_maxpool_input_pipe_671_inst_req_1;
      reqR_unguarded(7) <= RPIPE_maxpool_input_pipe_809_inst_req_1;
      reqR_unguarded(6) <= RPIPE_maxpool_input_pipe_825_inst_req_1;
      reqR_unguarded(5) <= RPIPE_maxpool_input_pipe_846_inst_req_1;
      reqR_unguarded(4) <= RPIPE_maxpool_input_pipe_867_inst_req_1;
      reqR_unguarded(3) <= RPIPE_maxpool_input_pipe_888_inst_req_1;
      reqR_unguarded(2) <= RPIPE_maxpool_input_pipe_909_inst_req_1;
      reqR_unguarded(1) <= RPIPE_maxpool_input_pipe_930_inst_req_1;
      reqR_unguarded(0) <= RPIPE_maxpool_input_pipe_951_inst_req_1;
      RPIPE_maxpool_input_pipe_1447_inst_ack_1 <= ackR_unguarded(33);
      RPIPE_maxpool_input_pipe_1580_inst_ack_1 <= ackR_unguarded(32);
      RPIPE_maxpool_input_pipe_1080_inst_ack_1 <= ackR_unguarded(31);
      RPIPE_maxpool_input_pipe_1305_inst_ack_1 <= ackR_unguarded(30);
      RPIPE_maxpool_input_pipe_1363_inst_ack_1 <= ackR_unguarded(29);
      RPIPE_maxpool_input_pipe_1384_inst_ack_1 <= ackR_unguarded(28);
      RPIPE_maxpool_input_pipe_1405_inst_ack_1 <= ackR_unguarded(27);
      RPIPE_maxpool_input_pipe_1321_inst_ack_1 <= ackR_unguarded(26);
      RPIPE_maxpool_input_pipe_438_inst_ack_1 <= ackR_unguarded(25);
      RPIPE_maxpool_input_pipe_1426_inst_ack_1 <= ackR_unguarded(24);
      RPIPE_maxpool_input_pipe_1342_inst_ack_1 <= ackR_unguarded(23);
      RPIPE_maxpool_input_pipe_454_inst_ack_1 <= ackR_unguarded(22);
      RPIPE_maxpool_input_pipe_469_inst_ack_1 <= ackR_unguarded(21);
      RPIPE_maxpool_input_pipe_485_inst_ack_1 <= ackR_unguarded(20);
      RPIPE_maxpool_input_pipe_500_inst_ack_1 <= ackR_unguarded(19);
      RPIPE_maxpool_input_pipe_516_inst_ack_1 <= ackR_unguarded(18);
      RPIPE_maxpool_input_pipe_531_inst_ack_1 <= ackR_unguarded(17);
      RPIPE_maxpool_input_pipe_547_inst_ack_1 <= ackR_unguarded(16);
      RPIPE_maxpool_input_pipe_562_inst_ack_1 <= ackR_unguarded(15);
      RPIPE_maxpool_input_pipe_578_inst_ack_1 <= ackR_unguarded(14);
      RPIPE_maxpool_input_pipe_593_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_maxpool_input_pipe_609_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_maxpool_input_pipe_624_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_maxpool_input_pipe_640_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_maxpool_input_pipe_655_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_maxpool_input_pipe_671_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_maxpool_input_pipe_809_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_maxpool_input_pipe_825_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_maxpool_input_pipe_846_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_maxpool_input_pipe_867_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_maxpool_input_pipe_888_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_maxpool_input_pipe_909_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_maxpool_input_pipe_930_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_maxpool_input_pipe_951_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      guard_vector(18)  <=  '1';
      guard_vector(19)  <=  '1';
      guard_vector(20)  <=  '1';
      guard_vector(21)  <=  '1';
      guard_vector(22)  <=  '1';
      guard_vector(23)  <=  '1';
      guard_vector(24)  <=  '1';
      guard_vector(25)  <=  '1';
      guard_vector(26)  <=  '1';
      guard_vector(27)  <=  '1';
      guard_vector(28)  <=  '1';
      guard_vector(29)  <=  '1';
      guard_vector(30)  <=  '1';
      guard_vector(31)  <=  '1';
      guard_vector(32)  <=  '1';
      guard_vector(33)  <=  '1';
      call328_1448 <= data_out(271 downto 264);
      callx_xi423_1581 <= data_out(263 downto 256);
      callx_xi_1081 <= data_out(255 downto 248);
      call260_1306 <= data_out(247 downto 240);
      call288_1364 <= data_out(239 downto 232);
      call298_1385 <= data_out(231 downto 224);
      call308_1406 <= data_out(223 downto 216);
      call268_1322 <= data_out(215 downto 208);
      call_439 <= data_out(207 downto 200);
      call318_1427 <= data_out(199 downto 192);
      call278_1343 <= data_out(191 downto 184);
      call6_455 <= data_out(183 downto 176);
      call14_470 <= data_out(175 downto 168);
      call23_486 <= data_out(167 downto 160);
      call32_501 <= data_out(159 downto 152);
      call41_517 <= data_out(151 downto 144);
      call50_532 <= data_out(143 downto 136);
      call59_548 <= data_out(135 downto 128);
      call68_563 <= data_out(127 downto 120);
      call77_579 <= data_out(119 downto 112);
      call86_594 <= data_out(111 downto 104);
      call95_610 <= data_out(103 downto 96);
      call104_625 <= data_out(95 downto 88);
      call113_641 <= data_out(87 downto 80);
      call122_656 <= data_out(79 downto 72);
      call131_672 <= data_out(71 downto 64);
      call153_810 <= data_out(63 downto 56);
      call161_826 <= data_out(55 downto 48);
      call171_847 <= data_out(47 downto 40);
      call181_868 <= data_out(39 downto 32);
      call191_889 <= data_out(31 downto 24);
      call201_910 <= data_out(23 downto 16);
      call211_931 <= data_out(15 downto 8);
      call221_952 <= data_out(7 downto 0);
      maxpool_input_pipe_read_0_gI: SplitGuardInterface generic map(name => "maxpool_input_pipe_read_0_gI", nreqs => 34, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      maxpool_input_pipe_read_0: InputPortRevised -- 
        generic map ( name => "maxpool_input_pipe_read_0", data_width => 8,  num_reqs => 34,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => maxpool_input_pipe_pipe_read_req(0),
          oack => maxpool_input_pipe_pipe_read_ack(0),
          odata => maxpool_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_elapsed_time_pipe_1798_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_elapsed_time_pipe_1798_inst_req_0;
      WPIPE_elapsed_time_pipe_1798_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_elapsed_time_pipe_1798_inst_req_1;
      WPIPE_elapsed_time_pipe_1798_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= sub415_1797;
      elapsed_time_pipe_write_0_gI: SplitGuardInterface generic map(name => "elapsed_time_pipe_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      elapsed_time_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "elapsed_time_pipe", data_width => 64, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => elapsed_time_pipe_pipe_write_req(0),
          oack => elapsed_time_pipe_pipe_write_ack(0),
          odata => elapsed_time_pipe_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_maxpool_output_pipe_440_inst WPIPE_maxpool_output_pipe_1449_inst WPIPE_maxpool_output_pipe_1344_inst WPIPE_maxpool_output_pipe_1082_inst WPIPE_maxpool_output_pipe_1365_inst WPIPE_maxpool_output_pipe_1307_inst WPIPE_maxpool_output_pipe_1386_inst WPIPE_maxpool_output_pipe_1582_inst WPIPE_maxpool_output_pipe_1407_inst WPIPE_maxpool_output_pipe_1323_inst WPIPE_maxpool_output_pipe_1428_inst WPIPE_maxpool_output_pipe_456_inst WPIPE_maxpool_output_pipe_471_inst WPIPE_maxpool_output_pipe_487_inst WPIPE_maxpool_output_pipe_502_inst WPIPE_maxpool_output_pipe_518_inst WPIPE_maxpool_output_pipe_533_inst WPIPE_maxpool_output_pipe_549_inst WPIPE_maxpool_output_pipe_564_inst WPIPE_maxpool_output_pipe_580_inst WPIPE_maxpool_output_pipe_595_inst WPIPE_maxpool_output_pipe_611_inst WPIPE_maxpool_output_pipe_626_inst WPIPE_maxpool_output_pipe_642_inst WPIPE_maxpool_output_pipe_657_inst WPIPE_maxpool_output_pipe_673_inst WPIPE_maxpool_output_pipe_811_inst WPIPE_maxpool_output_pipe_827_inst WPIPE_maxpool_output_pipe_848_inst WPIPE_maxpool_output_pipe_869_inst WPIPE_maxpool_output_pipe_890_inst WPIPE_maxpool_output_pipe_911_inst WPIPE_maxpool_output_pipe_932_inst WPIPE_maxpool_output_pipe_953_inst WPIPE_maxpool_output_pipe_1674_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(279 downto 0);
      signal sample_req, sample_ack : BooleanArray( 34 downto 0);
      signal update_req, update_ack : BooleanArray( 34 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 34 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 34 downto 0);
      signal guard_vector : std_logic_vector( 34 downto 0);
      constant inBUFs : IntegerArray(34 downto 0) := (34 => 0, 33 => 0, 32 => 0, 31 => 0, 30 => 0, 29 => 0, 28 => 0, 27 => 0, 26 => 0, 25 => 0, 24 => 0, 23 => 0, 22 => 0, 21 => 0, 20 => 0, 19 => 0, 18 => 0, 17 => 0, 16 => 0, 15 => 0, 14 => 0, 13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(34 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false, 17 => false, 18 => false, 19 => false, 20 => false, 21 => false, 22 => false, 23 => false, 24 => false, 25 => false, 26 => false, 27 => false, 28 => false, 29 => false, 30 => false, 31 => false, 32 => false, 33 => false, 34 => false);
      constant guardBuffering: IntegerArray(34 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2, 17 => 2, 18 => 2, 19 => 2, 20 => 2, 21 => 2, 22 => 2, 23 => 2, 24 => 2, 25 => 2, 26 => 2, 27 => 2, 28 => 2, 29 => 2, 30 => 2, 31 => 2, 32 => 2, 33 => 2, 34 => 2);
      -- 
    begin -- 
      sample_req_unguarded(34) <= WPIPE_maxpool_output_pipe_440_inst_req_0;
      sample_req_unguarded(33) <= WPIPE_maxpool_output_pipe_1449_inst_req_0;
      sample_req_unguarded(32) <= WPIPE_maxpool_output_pipe_1344_inst_req_0;
      sample_req_unguarded(31) <= WPIPE_maxpool_output_pipe_1082_inst_req_0;
      sample_req_unguarded(30) <= WPIPE_maxpool_output_pipe_1365_inst_req_0;
      sample_req_unguarded(29) <= WPIPE_maxpool_output_pipe_1307_inst_req_0;
      sample_req_unguarded(28) <= WPIPE_maxpool_output_pipe_1386_inst_req_0;
      sample_req_unguarded(27) <= WPIPE_maxpool_output_pipe_1582_inst_req_0;
      sample_req_unguarded(26) <= WPIPE_maxpool_output_pipe_1407_inst_req_0;
      sample_req_unguarded(25) <= WPIPE_maxpool_output_pipe_1323_inst_req_0;
      sample_req_unguarded(24) <= WPIPE_maxpool_output_pipe_1428_inst_req_0;
      sample_req_unguarded(23) <= WPIPE_maxpool_output_pipe_456_inst_req_0;
      sample_req_unguarded(22) <= WPIPE_maxpool_output_pipe_471_inst_req_0;
      sample_req_unguarded(21) <= WPIPE_maxpool_output_pipe_487_inst_req_0;
      sample_req_unguarded(20) <= WPIPE_maxpool_output_pipe_502_inst_req_0;
      sample_req_unguarded(19) <= WPIPE_maxpool_output_pipe_518_inst_req_0;
      sample_req_unguarded(18) <= WPIPE_maxpool_output_pipe_533_inst_req_0;
      sample_req_unguarded(17) <= WPIPE_maxpool_output_pipe_549_inst_req_0;
      sample_req_unguarded(16) <= WPIPE_maxpool_output_pipe_564_inst_req_0;
      sample_req_unguarded(15) <= WPIPE_maxpool_output_pipe_580_inst_req_0;
      sample_req_unguarded(14) <= WPIPE_maxpool_output_pipe_595_inst_req_0;
      sample_req_unguarded(13) <= WPIPE_maxpool_output_pipe_611_inst_req_0;
      sample_req_unguarded(12) <= WPIPE_maxpool_output_pipe_626_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_maxpool_output_pipe_642_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_maxpool_output_pipe_657_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_maxpool_output_pipe_673_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_maxpool_output_pipe_811_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_maxpool_output_pipe_827_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_maxpool_output_pipe_848_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_maxpool_output_pipe_869_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_maxpool_output_pipe_890_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_maxpool_output_pipe_911_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_maxpool_output_pipe_932_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_maxpool_output_pipe_953_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_maxpool_output_pipe_1674_inst_req_0;
      WPIPE_maxpool_output_pipe_440_inst_ack_0 <= sample_ack_unguarded(34);
      WPIPE_maxpool_output_pipe_1449_inst_ack_0 <= sample_ack_unguarded(33);
      WPIPE_maxpool_output_pipe_1344_inst_ack_0 <= sample_ack_unguarded(32);
      WPIPE_maxpool_output_pipe_1082_inst_ack_0 <= sample_ack_unguarded(31);
      WPIPE_maxpool_output_pipe_1365_inst_ack_0 <= sample_ack_unguarded(30);
      WPIPE_maxpool_output_pipe_1307_inst_ack_0 <= sample_ack_unguarded(29);
      WPIPE_maxpool_output_pipe_1386_inst_ack_0 <= sample_ack_unguarded(28);
      WPIPE_maxpool_output_pipe_1582_inst_ack_0 <= sample_ack_unguarded(27);
      WPIPE_maxpool_output_pipe_1407_inst_ack_0 <= sample_ack_unguarded(26);
      WPIPE_maxpool_output_pipe_1323_inst_ack_0 <= sample_ack_unguarded(25);
      WPIPE_maxpool_output_pipe_1428_inst_ack_0 <= sample_ack_unguarded(24);
      WPIPE_maxpool_output_pipe_456_inst_ack_0 <= sample_ack_unguarded(23);
      WPIPE_maxpool_output_pipe_471_inst_ack_0 <= sample_ack_unguarded(22);
      WPIPE_maxpool_output_pipe_487_inst_ack_0 <= sample_ack_unguarded(21);
      WPIPE_maxpool_output_pipe_502_inst_ack_0 <= sample_ack_unguarded(20);
      WPIPE_maxpool_output_pipe_518_inst_ack_0 <= sample_ack_unguarded(19);
      WPIPE_maxpool_output_pipe_533_inst_ack_0 <= sample_ack_unguarded(18);
      WPIPE_maxpool_output_pipe_549_inst_ack_0 <= sample_ack_unguarded(17);
      WPIPE_maxpool_output_pipe_564_inst_ack_0 <= sample_ack_unguarded(16);
      WPIPE_maxpool_output_pipe_580_inst_ack_0 <= sample_ack_unguarded(15);
      WPIPE_maxpool_output_pipe_595_inst_ack_0 <= sample_ack_unguarded(14);
      WPIPE_maxpool_output_pipe_611_inst_ack_0 <= sample_ack_unguarded(13);
      WPIPE_maxpool_output_pipe_626_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_maxpool_output_pipe_642_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_maxpool_output_pipe_657_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_maxpool_output_pipe_673_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_maxpool_output_pipe_811_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_maxpool_output_pipe_827_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_maxpool_output_pipe_848_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_maxpool_output_pipe_869_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_maxpool_output_pipe_890_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_maxpool_output_pipe_911_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_maxpool_output_pipe_932_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_maxpool_output_pipe_953_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_maxpool_output_pipe_1674_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(34) <= WPIPE_maxpool_output_pipe_440_inst_req_1;
      update_req_unguarded(33) <= WPIPE_maxpool_output_pipe_1449_inst_req_1;
      update_req_unguarded(32) <= WPIPE_maxpool_output_pipe_1344_inst_req_1;
      update_req_unguarded(31) <= WPIPE_maxpool_output_pipe_1082_inst_req_1;
      update_req_unguarded(30) <= WPIPE_maxpool_output_pipe_1365_inst_req_1;
      update_req_unguarded(29) <= WPIPE_maxpool_output_pipe_1307_inst_req_1;
      update_req_unguarded(28) <= WPIPE_maxpool_output_pipe_1386_inst_req_1;
      update_req_unguarded(27) <= WPIPE_maxpool_output_pipe_1582_inst_req_1;
      update_req_unguarded(26) <= WPIPE_maxpool_output_pipe_1407_inst_req_1;
      update_req_unguarded(25) <= WPIPE_maxpool_output_pipe_1323_inst_req_1;
      update_req_unguarded(24) <= WPIPE_maxpool_output_pipe_1428_inst_req_1;
      update_req_unguarded(23) <= WPIPE_maxpool_output_pipe_456_inst_req_1;
      update_req_unguarded(22) <= WPIPE_maxpool_output_pipe_471_inst_req_1;
      update_req_unguarded(21) <= WPIPE_maxpool_output_pipe_487_inst_req_1;
      update_req_unguarded(20) <= WPIPE_maxpool_output_pipe_502_inst_req_1;
      update_req_unguarded(19) <= WPIPE_maxpool_output_pipe_518_inst_req_1;
      update_req_unguarded(18) <= WPIPE_maxpool_output_pipe_533_inst_req_1;
      update_req_unguarded(17) <= WPIPE_maxpool_output_pipe_549_inst_req_1;
      update_req_unguarded(16) <= WPIPE_maxpool_output_pipe_564_inst_req_1;
      update_req_unguarded(15) <= WPIPE_maxpool_output_pipe_580_inst_req_1;
      update_req_unguarded(14) <= WPIPE_maxpool_output_pipe_595_inst_req_1;
      update_req_unguarded(13) <= WPIPE_maxpool_output_pipe_611_inst_req_1;
      update_req_unguarded(12) <= WPIPE_maxpool_output_pipe_626_inst_req_1;
      update_req_unguarded(11) <= WPIPE_maxpool_output_pipe_642_inst_req_1;
      update_req_unguarded(10) <= WPIPE_maxpool_output_pipe_657_inst_req_1;
      update_req_unguarded(9) <= WPIPE_maxpool_output_pipe_673_inst_req_1;
      update_req_unguarded(8) <= WPIPE_maxpool_output_pipe_811_inst_req_1;
      update_req_unguarded(7) <= WPIPE_maxpool_output_pipe_827_inst_req_1;
      update_req_unguarded(6) <= WPIPE_maxpool_output_pipe_848_inst_req_1;
      update_req_unguarded(5) <= WPIPE_maxpool_output_pipe_869_inst_req_1;
      update_req_unguarded(4) <= WPIPE_maxpool_output_pipe_890_inst_req_1;
      update_req_unguarded(3) <= WPIPE_maxpool_output_pipe_911_inst_req_1;
      update_req_unguarded(2) <= WPIPE_maxpool_output_pipe_932_inst_req_1;
      update_req_unguarded(1) <= WPIPE_maxpool_output_pipe_953_inst_req_1;
      update_req_unguarded(0) <= WPIPE_maxpool_output_pipe_1674_inst_req_1;
      WPIPE_maxpool_output_pipe_440_inst_ack_1 <= update_ack_unguarded(34);
      WPIPE_maxpool_output_pipe_1449_inst_ack_1 <= update_ack_unguarded(33);
      WPIPE_maxpool_output_pipe_1344_inst_ack_1 <= update_ack_unguarded(32);
      WPIPE_maxpool_output_pipe_1082_inst_ack_1 <= update_ack_unguarded(31);
      WPIPE_maxpool_output_pipe_1365_inst_ack_1 <= update_ack_unguarded(30);
      WPIPE_maxpool_output_pipe_1307_inst_ack_1 <= update_ack_unguarded(29);
      WPIPE_maxpool_output_pipe_1386_inst_ack_1 <= update_ack_unguarded(28);
      WPIPE_maxpool_output_pipe_1582_inst_ack_1 <= update_ack_unguarded(27);
      WPIPE_maxpool_output_pipe_1407_inst_ack_1 <= update_ack_unguarded(26);
      WPIPE_maxpool_output_pipe_1323_inst_ack_1 <= update_ack_unguarded(25);
      WPIPE_maxpool_output_pipe_1428_inst_ack_1 <= update_ack_unguarded(24);
      WPIPE_maxpool_output_pipe_456_inst_ack_1 <= update_ack_unguarded(23);
      WPIPE_maxpool_output_pipe_471_inst_ack_1 <= update_ack_unguarded(22);
      WPIPE_maxpool_output_pipe_487_inst_ack_1 <= update_ack_unguarded(21);
      WPIPE_maxpool_output_pipe_502_inst_ack_1 <= update_ack_unguarded(20);
      WPIPE_maxpool_output_pipe_518_inst_ack_1 <= update_ack_unguarded(19);
      WPIPE_maxpool_output_pipe_533_inst_ack_1 <= update_ack_unguarded(18);
      WPIPE_maxpool_output_pipe_549_inst_ack_1 <= update_ack_unguarded(17);
      WPIPE_maxpool_output_pipe_564_inst_ack_1 <= update_ack_unguarded(16);
      WPIPE_maxpool_output_pipe_580_inst_ack_1 <= update_ack_unguarded(15);
      WPIPE_maxpool_output_pipe_595_inst_ack_1 <= update_ack_unguarded(14);
      WPIPE_maxpool_output_pipe_611_inst_ack_1 <= update_ack_unguarded(13);
      WPIPE_maxpool_output_pipe_626_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_maxpool_output_pipe_642_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_maxpool_output_pipe_657_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_maxpool_output_pipe_673_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_maxpool_output_pipe_811_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_maxpool_output_pipe_827_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_maxpool_output_pipe_848_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_maxpool_output_pipe_869_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_maxpool_output_pipe_890_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_maxpool_output_pipe_911_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_maxpool_output_pipe_932_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_maxpool_output_pipe_953_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_maxpool_output_pipe_1674_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      guard_vector(18)  <=  '1';
      guard_vector(19)  <=  '1';
      guard_vector(20)  <=  '1';
      guard_vector(21)  <=  '1';
      guard_vector(22)  <=  '1';
      guard_vector(23)  <=  '1';
      guard_vector(24)  <=  '1';
      guard_vector(25)  <=  '1';
      guard_vector(26)  <=  '1';
      guard_vector(27)  <=  '1';
      guard_vector(28)  <=  '1';
      guard_vector(29)  <=  '1';
      guard_vector(30)  <=  '1';
      guard_vector(31)  <=  '1';
      guard_vector(32)  <=  '1';
      guard_vector(33)  <=  '1';
      guard_vector(34)  <=  '1';
      data_in <= call_439 & call328_1448 & call278_1343 & callx_xi_1081 & call288_1364 & call260_1306 & call298_1385 & callx_xi423_1581 & call308_1406 & call268_1322 & call318_1427 & call6_455 & call14_470 & call23_486 & call32_501 & call41_517 & call50_532 & call59_548 & call68_563 & call77_579 & call86_594 & call95_610 & call104_625 & call113_641 & call122_656 & call131_672 & call153_810 & call161_826 & call171_847 & call181_868 & call191_889 & call201_910 & call211_931 & call221_952 & type_cast_1676_wire_constant;
      maxpool_output_pipe_write_1_gI: SplitGuardInterface generic map(name => "maxpool_output_pipe_write_1_gI", nreqs => 35, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      maxpool_output_pipe_write_1: OutputPortRevised -- 
        generic map ( name => "maxpool_output_pipe", data_width => 8, num_reqs => 35, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => maxpool_output_pipe_pipe_write_req(0),
          oack => maxpool_output_pipe_pipe_write_ack(0),
          odata => maxpool_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_num_out_pipe_1671_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_num_out_pipe_1671_inst_req_0;
      WPIPE_num_out_pipe_1671_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_num_out_pipe_1671_inst_req_1;
      WPIPE_num_out_pipe_1671_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= mul375_1670;
      num_out_pipe_write_2_gI: SplitGuardInterface generic map(name => "num_out_pipe_write_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      num_out_pipe_write_2: OutputPortRevised -- 
        generic map ( name => "num_out_pipe", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => num_out_pipe_pipe_write_req(0),
          oack => num_out_pipe_pipe_write_ack(0),
          odata => num_out_pipe_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared call operator group (0) : call_stmt_1659_call call_stmt_1787_call 
    timer_call_group_0: Block -- 
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_1659_call_req_0;
      reqL_unguarded(0) <= call_stmt_1787_call_req_0;
      call_stmt_1659_call_ack_0 <= ackL_unguarded(1);
      call_stmt_1787_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_1659_call_req_1;
      reqR_unguarded(0) <= call_stmt_1787_call_req_1;
      call_stmt_1659_call_ack_1 <= ackR_unguarded(1);
      call_stmt_1787_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      timer_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      timer_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      timer_call_group_0_gI: SplitGuardInterface generic map(name => "timer_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      call355_1659 <= data_out(127 downto 64);
      call410_1787 <= data_out(63 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 2,
        nreqs => 2,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => timer_call_reqs(0),
          ackR => timer_call_acks(0),
          tagR => timer_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => timer_return_acks(0), -- cross-over
          ackL => timer_return_reqs(0), -- cross-over
          dataL => timer_return_data(63 downto 0),
          tagL => timer_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_1754_call 
    loadKernelChannel_call_group_1: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1754_call_req_0;
      call_stmt_1754_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1754_call_req_1;
      call_stmt_1754_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      loadKernelChannel_call_group_1_gI: SplitGuardInterface generic map(name => "loadKernelChannel_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= conv381_1747 & conv387_1751;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 128,
        owidth => 128,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => loadKernelChannel_call_reqs(0),
          ackR => loadKernelChannel_call_acks(0),
          dataR => loadKernelChannel_call_data(127 downto 0),
          tagR => loadKernelChannel_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => loadKernelChannel_return_acks(0), -- cross-over
          ackL => loadKernelChannel_return_reqs(0), -- cross-over
          tagL => loadKernelChannel_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- shared call operator group (2) : call_stmt_1761_call 
    access_T_call_group_2: Block -- 
      signal data_in: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1761_call_req_0;
      call_stmt_1761_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1761_call_req_1;
      call_stmt_1761_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      access_T_call_group_2_gI: SplitGuardInterface generic map(name => "access_T_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= mul362_1665 & add63_560 & sub_1683 & sub395_1689 & add45_529 & add27_498;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 96,
        owidth => 96,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => access_T_call_reqs(0),
          ackR => access_T_call_acks(0),
          dataR => access_T_call_data(95 downto 0),
          tagR => access_T_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => access_T_return_acks(0), -- cross-over
          ackL => access_T_return_reqs(0), -- cross-over
          tagL => access_T_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- 
  end Block; -- data_path
  -- 
end convolution3D_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convolve is -- 
  generic (tag_length : integer); 
  port ( -- 
    input_pipe1_pipe_read_req : out  std_logic_vector(0 downto 0);
    input_pipe1_pipe_read_ack : in   std_logic_vector(0 downto 0);
    input_pipe1_pipe_read_data : in   std_logic_vector(15 downto 0);
    num_out_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    num_out_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    num_out_pipe_pipe_read_data : in   std_logic_vector(15 downto 0);
    size_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    size_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    size_pipe_pipe_read_data : in   std_logic_vector(31 downto 0);
    kernel_pipe1_pipe_read_req : out  std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_read_ack : in   std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_read_data : in   std_logic_vector(15 downto 0);
    input_done_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    input_done_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    input_done_pipe_pipe_write_data : out  std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    kernel_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convolve;
architecture convolve_arch of convolve is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convolve_CP_4290_start: Boolean;
  signal convolve_CP_4290_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_num_out_pipe_1809_inst_req_0 : boolean;
  signal phi_stmt_1825_req_1 : boolean;
  signal phi_stmt_1829_req_0 : boolean;
  signal nacc_1880_1831_buf_req_0 : boolean;
  signal RPIPE_kernel_pipe1_1847_inst_ack_0 : boolean;
  signal n_out_count_1909_1837_buf_req_1 : boolean;
  signal RPIPE_kernel_pipe1_1847_inst_req_0 : boolean;
  signal RPIPE_size_pipe_1812_inst_ack_1 : boolean;
  signal RPIPE_size_pipe_1812_inst_req_1 : boolean;
  signal WPIPE_input_done_pipe_1916_inst_ack_0 : boolean;
  signal phi_stmt_1825_ack_0 : boolean;
  signal n_out_count_1909_1837_buf_ack_1 : boolean;
  signal WPIPE_input_done_pipe_1916_inst_req_1 : boolean;
  signal WPIPE_input_done_pipe_1916_inst_ack_1 : boolean;
  signal slice_1925_inst_req_0 : boolean;
  signal slice_1925_inst_ack_0 : boolean;
  signal do_while_stmt_1823_branch_req_0 : boolean;
  signal RPIPE_input_pipe1_1840_inst_req_0 : boolean;
  signal SUB_u32_u32_1861_inst_req_0 : boolean;
  signal RPIPE_input_pipe1_1840_inst_ack_0 : boolean;
  signal RPIPE_num_out_pipe_1809_inst_ack_0 : boolean;
  signal WPIPE_kernel_pipe1_1895_inst_ack_1 : boolean;
  signal W_next_sum_1903_delayed_1_0_1927_inst_ack_1 : boolean;
  signal type_cast_1933_inst_req_0 : boolean;
  signal type_cast_1933_inst_ack_0 : boolean;
  signal SUB_u32_u32_1861_inst_ack_0 : boolean;
  signal slice_1925_inst_ack_1 : boolean;
  signal RPIPE_input_pipe1_1840_inst_req_1 : boolean;
  signal W_next_sum_1903_delayed_1_0_1927_inst_req_1 : boolean;
  signal slice_1921_inst_req_1 : boolean;
  signal phi_stmt_1829_req_1 : boolean;
  signal RPIPE_input_pipe1_1840_inst_ack_1 : boolean;
  signal nacc_1880_1831_buf_ack_0 : boolean;
  signal slice_1925_inst_req_1 : boolean;
  signal phi_stmt_1825_req_0 : boolean;
  signal W_next_sum_1903_delayed_1_0_1927_inst_req_0 : boolean;
  signal W_next_sum_1903_delayed_1_0_1927_inst_ack_0 : boolean;
  signal RPIPE_size_pipe_1812_inst_req_0 : boolean;
  signal nmycount_1888_1828_buf_req_0 : boolean;
  signal SUB_u32_u32_1861_inst_req_1 : boolean;
  signal RPIPE_num_out_pipe_1809_inst_req_1 : boolean;
  signal SUB_u32_u32_1861_inst_ack_1 : boolean;
  signal RPIPE_kernel_pipe1_1847_inst_req_1 : boolean;
  signal WPIPE_kernel_pipe1_1895_inst_req_0 : boolean;
  signal nmycount_1888_1828_buf_ack_0 : boolean;
  signal RPIPE_num_out_pipe_1809_inst_ack_1 : boolean;
  signal phi_stmt_1829_ack_0 : boolean;
  signal nmycount_1888_1828_buf_req_1 : boolean;
  signal slice_1921_inst_req_0 : boolean;
  signal WPIPE_kernel_pipe1_1895_inst_ack_0 : boolean;
  signal nmycount_1888_1828_buf_ack_1 : boolean;
  signal RPIPE_size_pipe_1812_inst_ack_0 : boolean;
  signal nacc_1880_1831_buf_req_1 : boolean;
  signal slice_1921_inst_ack_0 : boolean;
  signal nacc_1880_1831_buf_ack_1 : boolean;
  signal slice_1921_inst_ack_1 : boolean;
  signal WPIPE_kernel_pipe1_1895_inst_req_1 : boolean;
  signal n_out_count_1909_1837_buf_req_0 : boolean;
  signal WPIPE_input_done_pipe_1916_inst_req_0 : boolean;
  signal phi_stmt_1833_ack_0 : boolean;
  signal phi_stmt_1833_req_0 : boolean;
  signal phi_stmt_1833_req_1 : boolean;
  signal RPIPE_kernel_pipe1_1847_inst_ack_1 : boolean;
  signal n_out_count_1909_1837_buf_ack_0 : boolean;
  signal type_cast_1933_inst_req_1 : boolean;
  signal type_cast_1933_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1931_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1931_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1931_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1931_inst_ack_1 : boolean;
  signal W_next_sum_1908_delayed_1_0_1935_inst_req_0 : boolean;
  signal W_next_sum_1908_delayed_1_0_1935_inst_ack_0 : boolean;
  signal W_next_sum_1908_delayed_1_0_1935_inst_req_1 : boolean;
  signal W_next_sum_1908_delayed_1_0_1935_inst_ack_1 : boolean;
  signal type_cast_1941_inst_req_0 : boolean;
  signal type_cast_1941_inst_ack_0 : boolean;
  signal type_cast_1941_inst_req_1 : boolean;
  signal type_cast_1941_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1939_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1939_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1939_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1939_inst_ack_1 : boolean;
  signal do_while_stmt_1823_branch_ack_0 : boolean;
  signal do_while_stmt_1823_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convolve_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convolve_CP_4290_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convolve_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convolve_CP_4290_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convolve_CP_4290_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convolve_CP_4290_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convolve_CP_4290: Block -- control-path 
    signal convolve_CP_4290_elements: BooleanArray(127 downto 0);
    -- 
  begin -- 
    convolve_CP_4290_elements(0) <= convolve_CP_4290_start;
    convolve_CP_4290_symbol <= convolve_CP_4290_elements(1);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	4 
    -- CP-element group 0:  members (11) 
      -- CP-element group 0: 	 branch_block_stmt_1807/assign_stmt_1810_to_assign_stmt_1822/RPIPE_num_out_pipe_1809_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1807/assign_stmt_1810_to_assign_stmt_1822__entry__
      -- CP-element group 0: 	 branch_block_stmt_1807/assign_stmt_1810_to_assign_stmt_1822/RPIPE_num_out_pipe_1809_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_1807/assign_stmt_1810_to_assign_stmt_1822/RPIPE_num_out_pipe_1809_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1807/branch_block_stmt_1807__entry__
      -- CP-element group 0: 	 branch_block_stmt_1807/assign_stmt_1810_to_assign_stmt_1822/$entry
      -- CP-element group 0: 	 branch_block_stmt_1807/$entry
      -- CP-element group 0: 	 branch_block_stmt_1807/assign_stmt_1810_to_assign_stmt_1822/RPIPE_size_pipe_1812_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1807/assign_stmt_1810_to_assign_stmt_1822/RPIPE_size_pipe_1812_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_1807/assign_stmt_1810_to_assign_stmt_1822/RPIPE_size_pipe_1812_sample_start_
      -- CP-element group 0: 	 $entry
      -- 
    rr_4312_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4312_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4290_elements(0), ack => RPIPE_num_out_pipe_1809_inst_req_0); -- 
    rr_4326_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4326_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4290_elements(0), ack => RPIPE_size_pipe_1812_inst_req_0); -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	127 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 branch_block_stmt_1807/do_while_stmt_1823__exit__
      -- CP-element group 1: 	 branch_block_stmt_1807/branch_block_stmt_1807__exit__
      -- CP-element group 1: 	 branch_block_stmt_1807/$exit
      -- CP-element group 1: 	 $exit
      -- 
    convolve_CP_4290_elements(1) <= convolve_CP_4290_elements(127);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_1807/assign_stmt_1810_to_assign_stmt_1822/RPIPE_num_out_pipe_1809_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_1807/assign_stmt_1810_to_assign_stmt_1822/RPIPE_num_out_pipe_1809_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1807/assign_stmt_1810_to_assign_stmt_1822/RPIPE_num_out_pipe_1809_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_1807/assign_stmt_1810_to_assign_stmt_1822/RPIPE_num_out_pipe_1809_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_1807/assign_stmt_1810_to_assign_stmt_1822/RPIPE_num_out_pipe_1809_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1807/assign_stmt_1810_to_assign_stmt_1822/RPIPE_num_out_pipe_1809_Update/cr
      -- 
    ra_4313_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_num_out_pipe_1809_inst_ack_0, ack => convolve_CP_4290_elements(2)); -- 
    cr_4317_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4317_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4290_elements(2), ack => RPIPE_num_out_pipe_1809_inst_req_1); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	6 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_1807/assign_stmt_1810_to_assign_stmt_1822/RPIPE_num_out_pipe_1809_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_1807/assign_stmt_1810_to_assign_stmt_1822/RPIPE_num_out_pipe_1809_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_1807/assign_stmt_1810_to_assign_stmt_1822/RPIPE_num_out_pipe_1809_Update/ca
      -- 
    ca_4318_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_num_out_pipe_1809_inst_ack_1, ack => convolve_CP_4290_elements(3)); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_1807/assign_stmt_1810_to_assign_stmt_1822/RPIPE_size_pipe_1812_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_1807/assign_stmt_1810_to_assign_stmt_1822/RPIPE_size_pipe_1812_Update/cr
      -- CP-element group 4: 	 branch_block_stmt_1807/assign_stmt_1810_to_assign_stmt_1822/RPIPE_size_pipe_1812_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_1807/assign_stmt_1810_to_assign_stmt_1822/RPIPE_size_pipe_1812_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_1807/assign_stmt_1810_to_assign_stmt_1822/RPIPE_size_pipe_1812_update_start_
      -- CP-element group 4: 	 branch_block_stmt_1807/assign_stmt_1810_to_assign_stmt_1822/RPIPE_size_pipe_1812_Update/$entry
      -- 
    ra_4327_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_size_pipe_1812_inst_ack_0, ack => convolve_CP_4290_elements(4)); -- 
    cr_4331_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4331_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4290_elements(4), ack => RPIPE_size_pipe_1812_inst_req_1); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1807/assign_stmt_1810_to_assign_stmt_1822/RPIPE_size_pipe_1812_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_1807/assign_stmt_1810_to_assign_stmt_1822/RPIPE_size_pipe_1812_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_1807/assign_stmt_1810_to_assign_stmt_1822/RPIPE_size_pipe_1812_update_completed_
      -- 
    ca_4332_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_size_pipe_1812_inst_ack_1, ack => convolve_CP_4290_elements(5)); -- 
    -- CP-element group 6:  join  transition  place  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	3 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_1807/do_while_stmt_1823__entry__
      -- CP-element group 6: 	 branch_block_stmt_1807/assign_stmt_1810_to_assign_stmt_1822__exit__
      -- CP-element group 6: 	 branch_block_stmt_1807/assign_stmt_1810_to_assign_stmt_1822/$exit
      -- 
    convolve_cp_element_group_6: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "convolve_cp_element_group_6"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4290_elements(3) & convolve_CP_4290_elements(5);
      gj_convolve_cp_element_group_6 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4290_elements(6), clk => clk, reset => reset); --
    end block;
    -- CP-element group 7:  transition  place  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	13 
    -- CP-element group 7:  members (2) 
      -- CP-element group 7: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823__entry__
      -- CP-element group 7: 	 branch_block_stmt_1807/do_while_stmt_1823/$entry
      -- 
    convolve_CP_4290_elements(7) <= convolve_CP_4290_elements(6);
    -- CP-element group 8:  merge  place  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	127 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823__exit__
      -- 
    -- Element group convolve_CP_4290_elements(8) is bound as output of CP function.
    -- CP-element group 9:  merge  place  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	12 
    -- CP-element group 9:  members (1) 
      -- CP-element group 9: 	 branch_block_stmt_1807/do_while_stmt_1823/loop_back
      -- 
    -- Element group convolve_CP_4290_elements(9) is bound as output of CP function.
    -- CP-element group 10:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	15 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	125 
    -- CP-element group 10: 	126 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_1807/do_while_stmt_1823/condition_done
      -- CP-element group 10: 	 branch_block_stmt_1807/do_while_stmt_1823/loop_exit/$entry
      -- CP-element group 10: 	 branch_block_stmt_1807/do_while_stmt_1823/loop_taken/$entry
      -- 
    convolve_CP_4290_elements(10) <= convolve_CP_4290_elements(15);
    -- CP-element group 11:  branch  place  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	124 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (1) 
      -- CP-element group 11: 	 branch_block_stmt_1807/do_while_stmt_1823/loop_body_done
      -- 
    convolve_CP_4290_elements(11) <= convolve_CP_4290_elements(124);
    -- CP-element group 12:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	9 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	62 
    -- CP-element group 12: 	45 
    -- CP-element group 12: 	26 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/back_edge_to_loop_body
      -- 
    convolve_CP_4290_elements(12) <= convolve_CP_4290_elements(9);
    -- CP-element group 13:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	7 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	64 
    -- CP-element group 13: 	47 
    -- CP-element group 13: 	28 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/first_time_through_loop_body
      -- 
    convolve_CP_4290_elements(13) <= convolve_CP_4290_elements(7);
    -- CP-element group 14:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	58 
    -- CP-element group 14: 	59 
    -- CP-element group 14: 	39 
    -- CP-element group 14: 	40 
    -- CP-element group 14: 	123 
    -- CP-element group 14: 	20 
    -- CP-element group 14: 	21 
    -- CP-element group 14: 	75 
    -- CP-element group 14: 	79 
    -- CP-element group 14: 	83 
    -- CP-element group 14:  members (2) 
      -- CP-element group 14: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/$entry
      -- CP-element group 14: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/loop_body_start
      -- 
    -- Element group convolve_CP_4290_elements(14) is bound as output of CP function.
    -- CP-element group 15:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	123 
    -- CP-element group 15: 	19 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	10 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/condition_evaluated
      -- 
    condition_evaluated_4347_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_4347_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4290_elements(15), ack => do_while_stmt_1823_branch_req_0); -- 
    convolve_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4290_elements(123) & convolve_CP_4290_elements(19);
      gj_convolve_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4290_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	58 
    -- CP-element group 16: 	39 
    -- CP-element group 16: 	20 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	19 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	41 
    -- CP-element group 16: 	22 
    -- CP-element group 16:  members (2) 
      -- CP-element group 16: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/aggregated_phi_sample_req
      -- CP-element group 16: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/phi_stmt_1833_sample_start__ps
      -- 
    convolve_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4290_elements(58) & convolve_CP_4290_elements(39) & convolve_CP_4290_elements(20) & convolve_CP_4290_elements(19);
      gj_convolve_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4290_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	60 
    -- CP-element group 17: 	42 
    -- CP-element group 17: 	23 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	76 
    -- CP-element group 17: 	80 
    -- CP-element group 17: 	84 
    -- CP-element group 17: marked-successors 
    -- CP-element group 17: 	58 
    -- CP-element group 17: 	39 
    -- CP-element group 17: 	20 
    -- CP-element group 17:  members (4) 
      -- CP-element group 17: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/aggregated_phi_sample_ack
      -- CP-element group 17: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/phi_stmt_1829_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/phi_stmt_1825_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/phi_stmt_1833_sample_completed_
      -- 
    convolve_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4290_elements(60) & convolve_CP_4290_elements(42) & convolve_CP_4290_elements(23);
      gj_convolve_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4290_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	59 
    -- CP-element group 18: 	40 
    -- CP-element group 18: 	21 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	43 
    -- CP-element group 18: 	24 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/aggregated_phi_update_req
      -- CP-element group 18: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/phi_stmt_1833_update_start__ps
      -- 
    convolve_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4290_elements(59) & convolve_CP_4290_elements(40) & convolve_CP_4290_elements(21);
      gj_convolve_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4290_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	61 
    -- CP-element group 19: 	44 
    -- CP-element group 19: 	25 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	15 
    -- CP-element group 19: marked-successors 
    -- CP-element group 19: 	16 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/aggregated_phi_update_ack
      -- 
    convolve_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4290_elements(61) & convolve_CP_4290_elements(44) & convolve_CP_4290_elements(25);
      gj_convolve_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4290_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  join  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	14 
    -- CP-element group 20: marked-predecessors 
    -- CP-element group 20: 	17 
    -- CP-element group 20: 	86 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	16 
    -- CP-element group 20:  members (1) 
      -- CP-element group 20: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/phi_stmt_1825_sample_start_
      -- 
    convolve_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4290_elements(14) & convolve_CP_4290_elements(17) & convolve_CP_4290_elements(86);
      gj_convolve_cp_element_group_20 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4290_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  join  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	14 
    -- CP-element group 21: marked-predecessors 
    -- CP-element group 21: 	114 
    -- CP-element group 21: 	91 
    -- CP-element group 21: 	103 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	18 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/phi_stmt_1825_update_start_
      -- 
    convolve_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4290_elements(14) & convolve_CP_4290_elements(114) & convolve_CP_4290_elements(91) & convolve_CP_4290_elements(103);
      gj_convolve_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4290_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	16 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (1) 
      -- CP-element group 22: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/phi_stmt_1825_sample_start__ps
      -- 
    convolve_CP_4290_elements(22) <= convolve_CP_4290_elements(16);
    -- CP-element group 23:  join  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	17 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/phi_stmt_1825_sample_completed__ps
      -- 
    -- Element group convolve_CP_4290_elements(23) is bound as output of CP function.
    -- CP-element group 24:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	18 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/phi_stmt_1825_update_start__ps
      -- 
    convolve_CP_4290_elements(24) <= convolve_CP_4290_elements(18);
    -- CP-element group 25:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	112 
    -- CP-element group 25: 	19 
    -- CP-element group 25: 	90 
    -- CP-element group 25: 	101 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/phi_stmt_1825_update_completed__ps
      -- CP-element group 25: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/phi_stmt_1825_update_completed_
      -- 
    -- Element group convolve_CP_4290_elements(25) is bound as output of CP function.
    -- CP-element group 26:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	12 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/phi_stmt_1825_loopback_trigger
      -- 
    convolve_CP_4290_elements(26) <= convolve_CP_4290_elements(12);
    -- CP-element group 27:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (2) 
      -- CP-element group 27: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/phi_stmt_1825_loopback_sample_req
      -- CP-element group 27: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/phi_stmt_1825_loopback_sample_req_ps
      -- 
    phi_stmt_1825_loopback_sample_req_4362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1825_loopback_sample_req_4362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4290_elements(27), ack => phi_stmt_1825_req_1); -- 
    -- Element group convolve_CP_4290_elements(27) is bound as output of CP function.
    -- CP-element group 28:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	13 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/phi_stmt_1825_entry_trigger
      -- 
    convolve_CP_4290_elements(28) <= convolve_CP_4290_elements(13);
    -- CP-element group 29:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (2) 
      -- CP-element group 29: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/phi_stmt_1825_entry_sample_req
      -- CP-element group 29: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/phi_stmt_1825_entry_sample_req_ps
      -- 
    phi_stmt_1825_entry_sample_req_4365_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1825_entry_sample_req_4365_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4290_elements(29), ack => phi_stmt_1825_req_0); -- 
    -- Element group convolve_CP_4290_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (2) 
      -- CP-element group 30: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/phi_stmt_1825_phi_mux_ack_ps
      -- CP-element group 30: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/phi_stmt_1825_phi_mux_ack
      -- 
    phi_stmt_1825_phi_mux_ack_4368_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1825_ack_0, ack => convolve_CP_4290_elements(30)); -- 
    -- CP-element group 31:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/R_mcount_var_1827_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/R_mcount_var_1827_sample_completed_
      -- CP-element group 31: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/R_mcount_var_1827_sample_completed__ps
      -- CP-element group 31: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/R_mcount_var_1827_sample_start__ps
      -- 
    -- Element group convolve_CP_4290_elements(31) is bound as output of CP function.
    -- CP-element group 32:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	34 
    -- CP-element group 32:  members (2) 
      -- CP-element group 32: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/R_mcount_var_1827_update_start_
      -- CP-element group 32: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/R_mcount_var_1827_update_start__ps
      -- 
    -- Element group convolve_CP_4290_elements(32) is bound as output of CP function.
    -- CP-element group 33:  join  transition  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	34 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (1) 
      -- CP-element group 33: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/R_mcount_var_1827_update_completed__ps
      -- 
    convolve_CP_4290_elements(33) <= convolve_CP_4290_elements(34);
    -- CP-element group 34:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	32 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	33 
    -- CP-element group 34:  members (1) 
      -- CP-element group 34: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/R_mcount_var_1827_update_completed_
      -- 
    -- Element group convolve_CP_4290_elements(34) is a control-delay.
    cp_element_34_delay: control_delay_element  generic map(name => " 34_delay", delay_value => 1)  port map(req => convolve_CP_4290_elements(32), ack => convolve_CP_4290_elements(34), clk => clk, reset =>reset);
    -- CP-element group 35:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	37 
    -- CP-element group 35:  members (4) 
      -- CP-element group 35: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/R_nmycount_1828_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/R_nmycount_1828_sample_start__ps
      -- CP-element group 35: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/R_nmycount_1828_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/R_nmycount_1828_Sample/req
      -- 
    req_4389_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4389_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4290_elements(35), ack => nmycount_1888_1828_buf_req_0); -- 
    -- Element group convolve_CP_4290_elements(35) is bound as output of CP function.
    -- CP-element group 36:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	38 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/R_nmycount_1828_update_start_
      -- CP-element group 36: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/R_nmycount_1828_update_start__ps
      -- CP-element group 36: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/R_nmycount_1828_Update/$entry
      -- CP-element group 36: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/R_nmycount_1828_Update/req
      -- 
    req_4394_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4394_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4290_elements(36), ack => nmycount_1888_1828_buf_req_1); -- 
    -- Element group convolve_CP_4290_elements(36) is bound as output of CP function.
    -- CP-element group 37:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	35 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (4) 
      -- CP-element group 37: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/R_nmycount_1828_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/R_nmycount_1828_sample_completed__ps
      -- CP-element group 37: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/R_nmycount_1828_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/R_nmycount_1828_Sample/ack
      -- 
    ack_4390_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmycount_1888_1828_buf_ack_0, ack => convolve_CP_4290_elements(37)); -- 
    -- CP-element group 38:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	36 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (4) 
      -- CP-element group 38: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/R_nmycount_1828_update_completed__ps
      -- CP-element group 38: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/R_nmycount_1828_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/R_nmycount_1828_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/R_nmycount_1828_Update/ack
      -- 
    ack_4395_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmycount_1888_1828_buf_ack_1, ack => convolve_CP_4290_elements(38)); -- 
    -- CP-element group 39:  join  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	14 
    -- CP-element group 39: marked-predecessors 
    -- CP-element group 39: 	78 
    -- CP-element group 39: 	17 
    -- CP-element group 39: 	82 
    -- CP-element group 39: 	86 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	16 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/phi_stmt_1829_sample_start_
      -- 
    convolve_cp_element_group_39: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 1,3 => 0,4 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_39"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_4290_elements(14) & convolve_CP_4290_elements(78) & convolve_CP_4290_elements(17) & convolve_CP_4290_elements(82) & convolve_CP_4290_elements(86);
      gj_convolve_cp_element_group_39 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4290_elements(39), clk => clk, reset => reset); --
    end block;
    -- CP-element group 40:  join  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	14 
    -- CP-element group 40: marked-predecessors 
    -- CP-element group 40: 	95 
    -- CP-element group 40: 	99 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	18 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/phi_stmt_1829_update_start_
      -- 
    convolve_cp_element_group_40: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_40"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4290_elements(14) & convolve_CP_4290_elements(95) & convolve_CP_4290_elements(99);
      gj_convolve_cp_element_group_40 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4290_elements(40), clk => clk, reset => reset); --
    end block;
    -- CP-element group 41:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	16 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/phi_stmt_1829_sample_start__ps
      -- 
    convolve_CP_4290_elements(41) <= convolve_CP_4290_elements(16);
    -- CP-element group 42:  join  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	17 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/phi_stmt_1829_sample_completed__ps
      -- 
    -- Element group convolve_CP_4290_elements(42) is bound as output of CP function.
    -- CP-element group 43:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	18 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (1) 
      -- CP-element group 43: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/phi_stmt_1829_update_start__ps
      -- 
    convolve_CP_4290_elements(43) <= convolve_CP_4290_elements(18);
    -- CP-element group 44:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	93 
    -- CP-element group 44: 	97 
    -- CP-element group 44: 	19 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/phi_stmt_1829_update_completed__ps
      -- CP-element group 44: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/phi_stmt_1829_update_completed_
      -- 
    -- Element group convolve_CP_4290_elements(44) is bound as output of CP function.
    -- CP-element group 45:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	12 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/phi_stmt_1829_loopback_trigger
      -- 
    convolve_CP_4290_elements(45) <= convolve_CP_4290_elements(12);
    -- CP-element group 46:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/phi_stmt_1829_loopback_sample_req
      -- CP-element group 46: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/phi_stmt_1829_loopback_sample_req_ps
      -- 
    phi_stmt_1829_loopback_sample_req_4406_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1829_loopback_sample_req_4406_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4290_elements(46), ack => phi_stmt_1829_req_0); -- 
    -- Element group convolve_CP_4290_elements(46) is bound as output of CP function.
    -- CP-element group 47:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	13 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/phi_stmt_1829_entry_trigger
      -- 
    convolve_CP_4290_elements(47) <= convolve_CP_4290_elements(13);
    -- CP-element group 48:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (2) 
      -- CP-element group 48: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/phi_stmt_1829_entry_sample_req
      -- CP-element group 48: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/phi_stmt_1829_entry_sample_req_ps
      -- 
    phi_stmt_1829_entry_sample_req_4409_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1829_entry_sample_req_4409_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4290_elements(48), ack => phi_stmt_1829_req_1); -- 
    -- Element group convolve_CP_4290_elements(48) is bound as output of CP function.
    -- CP-element group 49:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (2) 
      -- CP-element group 49: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/phi_stmt_1829_phi_mux_ack
      -- CP-element group 49: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/phi_stmt_1829_phi_mux_ack_ps
      -- 
    phi_stmt_1829_phi_mux_ack_4412_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1829_ack_0, ack => convolve_CP_4290_elements(49)); -- 
    -- CP-element group 50:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (4) 
      -- CP-element group 50: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/R_nacc_1831_Sample/req
      -- CP-element group 50: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/R_nacc_1831_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/R_nacc_1831_sample_start__ps
      -- CP-element group 50: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/R_nacc_1831_Sample/$entry
      -- 
    req_4425_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4425_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4290_elements(50), ack => nacc_1880_1831_buf_req_0); -- 
    -- Element group convolve_CP_4290_elements(50) is bound as output of CP function.
    -- CP-element group 51:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	53 
    -- CP-element group 51:  members (4) 
      -- CP-element group 51: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/R_nacc_1831_update_start__ps
      -- CP-element group 51: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/R_nacc_1831_Update/$entry
      -- CP-element group 51: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/R_nacc_1831_update_start_
      -- CP-element group 51: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/R_nacc_1831_Update/req
      -- 
    req_4430_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4430_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4290_elements(51), ack => nacc_1880_1831_buf_req_1); -- 
    -- Element group convolve_CP_4290_elements(51) is bound as output of CP function.
    -- CP-element group 52:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (4) 
      -- CP-element group 52: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/R_nacc_1831_sample_completed__ps
      -- CP-element group 52: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/R_nacc_1831_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/R_nacc_1831_Sample/ack
      -- CP-element group 52: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/R_nacc_1831_sample_completed_
      -- 
    ack_4426_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nacc_1880_1831_buf_ack_0, ack => convolve_CP_4290_elements(52)); -- 
    -- CP-element group 53:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	51 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (4) 
      -- CP-element group 53: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/R_nacc_1831_update_completed__ps
      -- CP-element group 53: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/R_nacc_1831_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/R_nacc_1831_Update/ack
      -- CP-element group 53: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/R_nacc_1831_update_completed_
      -- 
    ack_4431_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nacc_1880_1831_buf_ack_1, ack => convolve_CP_4290_elements(53)); -- 
    -- CP-element group 54:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (4) 
      -- CP-element group 54: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/R_acc_var_1832_sample_start__ps
      -- CP-element group 54: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/R_acc_var_1832_sample_completed__ps
      -- CP-element group 54: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/R_acc_var_1832_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/R_acc_var_1832_sample_start_
      -- 
    -- Element group convolve_CP_4290_elements(54) is bound as output of CP function.
    -- CP-element group 55:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	57 
    -- CP-element group 55:  members (2) 
      -- CP-element group 55: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/R_acc_var_1832_update_start__ps
      -- CP-element group 55: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/R_acc_var_1832_update_start_
      -- 
    -- Element group convolve_CP_4290_elements(55) is bound as output of CP function.
    -- CP-element group 56:  join  transition  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	57 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (1) 
      -- CP-element group 56: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/R_acc_var_1832_update_completed__ps
      -- 
    convolve_CP_4290_elements(56) <= convolve_CP_4290_elements(57);
    -- CP-element group 57:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	55 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	56 
    -- CP-element group 57:  members (1) 
      -- CP-element group 57: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/R_acc_var_1832_update_completed_
      -- 
    -- Element group convolve_CP_4290_elements(57) is a control-delay.
    cp_element_57_delay: control_delay_element  generic map(name => " 57_delay", delay_value => 1)  port map(req => convolve_CP_4290_elements(55), ack => convolve_CP_4290_elements(57), clk => clk, reset =>reset);
    -- CP-element group 58:  join  transition  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	14 
    -- CP-element group 58: marked-predecessors 
    -- CP-element group 58: 	17 
    -- CP-element group 58: 	86 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	16 
    -- CP-element group 58:  members (1) 
      -- CP-element group 58: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/phi_stmt_1833_sample_start_
      -- 
    convolve_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4290_elements(14) & convolve_CP_4290_elements(17) & convolve_CP_4290_elements(86);
      gj_convolve_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4290_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  join  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	14 
    -- CP-element group 59: marked-predecessors 
    -- CP-element group 59: 	91 
    -- CP-element group 59: 	88 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	18 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/phi_stmt_1833_update_start_
      -- 
    convolve_cp_element_group_59: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_59"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4290_elements(14) & convolve_CP_4290_elements(91) & convolve_CP_4290_elements(88);
      gj_convolve_cp_element_group_59 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4290_elements(59), clk => clk, reset => reset); --
    end block;
    -- CP-element group 60:  join  transition  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	17 
    -- CP-element group 60:  members (1) 
      -- CP-element group 60: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/phi_stmt_1833_sample_completed__ps
      -- 
    -- Element group convolve_CP_4290_elements(60) is bound as output of CP function.
    -- CP-element group 61:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	19 
    -- CP-element group 61: 	87 
    -- CP-element group 61: 	90 
    -- CP-element group 61:  members (2) 
      -- CP-element group 61: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/phi_stmt_1833_update_completed__ps
      -- CP-element group 61: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/phi_stmt_1833_update_completed_
      -- 
    -- Element group convolve_CP_4290_elements(61) is bound as output of CP function.
    -- CP-element group 62:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	12 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (1) 
      -- CP-element group 62: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/phi_stmt_1833_loopback_trigger
      -- 
    convolve_CP_4290_elements(62) <= convolve_CP_4290_elements(12);
    -- CP-element group 63:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (2) 
      -- CP-element group 63: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/phi_stmt_1833_loopback_sample_req_ps
      -- CP-element group 63: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/phi_stmt_1833_loopback_sample_req
      -- 
    phi_stmt_1833_loopback_sample_req_4450_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1833_loopback_sample_req_4450_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4290_elements(63), ack => phi_stmt_1833_req_1); -- 
    -- Element group convolve_CP_4290_elements(63) is bound as output of CP function.
    -- CP-element group 64:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	13 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (1) 
      -- CP-element group 64: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/phi_stmt_1833_entry_trigger
      -- 
    convolve_CP_4290_elements(64) <= convolve_CP_4290_elements(13);
    -- CP-element group 65:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (2) 
      -- CP-element group 65: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/phi_stmt_1833_entry_sample_req_ps
      -- CP-element group 65: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/phi_stmt_1833_entry_sample_req
      -- 
    phi_stmt_1833_entry_sample_req_4453_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1833_entry_sample_req_4453_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4290_elements(65), ack => phi_stmt_1833_req_0); -- 
    -- Element group convolve_CP_4290_elements(65) is bound as output of CP function.
    -- CP-element group 66:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (2) 
      -- CP-element group 66: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/phi_stmt_1833_phi_mux_ack_ps
      -- CP-element group 66: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/phi_stmt_1833_phi_mux_ack
      -- 
    phi_stmt_1833_phi_mux_ack_4456_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1833_ack_0, ack => convolve_CP_4290_elements(66)); -- 
    -- CP-element group 67:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (4) 
      -- CP-element group 67: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/type_cast_1836_sample_start_
      -- CP-element group 67: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/type_cast_1836_sample_completed_
      -- CP-element group 67: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/type_cast_1836_sample_completed__ps
      -- CP-element group 67: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/type_cast_1836_sample_start__ps
      -- 
    -- Element group convolve_CP_4290_elements(67) is bound as output of CP function.
    -- CP-element group 68:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (2) 
      -- CP-element group 68: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/type_cast_1836_update_start_
      -- CP-element group 68: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/type_cast_1836_update_start__ps
      -- 
    -- Element group convolve_CP_4290_elements(68) is bound as output of CP function.
    -- CP-element group 69:  join  transition  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	70 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (1) 
      -- CP-element group 69: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/type_cast_1836_update_completed__ps
      -- 
    convolve_CP_4290_elements(69) <= convolve_CP_4290_elements(70);
    -- CP-element group 70:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	69 
    -- CP-element group 70:  members (1) 
      -- CP-element group 70: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/type_cast_1836_update_completed_
      -- 
    -- Element group convolve_CP_4290_elements(70) is a control-delay.
    cp_element_70_delay: control_delay_element  generic map(name => " 70_delay", delay_value => 1)  port map(req => convolve_CP_4290_elements(68), ack => convolve_CP_4290_elements(70), clk => clk, reset =>reset);
    -- CP-element group 71:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (4) 
      -- CP-element group 71: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/R_n_out_count_1837_sample_start_
      -- CP-element group 71: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/R_n_out_count_1837_sample_start__ps
      -- CP-element group 71: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/R_n_out_count_1837_Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/R_n_out_count_1837_Sample/req
      -- 
    req_4477_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4477_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4290_elements(71), ack => n_out_count_1909_1837_buf_req_0); -- 
    -- Element group convolve_CP_4290_elements(71) is bound as output of CP function.
    -- CP-element group 72:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	74 
    -- CP-element group 72:  members (4) 
      -- CP-element group 72: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/R_n_out_count_1837_Update/req
      -- CP-element group 72: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/R_n_out_count_1837_update_start__ps
      -- CP-element group 72: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/R_n_out_count_1837_update_start_
      -- CP-element group 72: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/R_n_out_count_1837_Update/$entry
      -- 
    req_4482_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4482_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4290_elements(72), ack => n_out_count_1909_1837_buf_req_1); -- 
    -- Element group convolve_CP_4290_elements(72) is bound as output of CP function.
    -- CP-element group 73:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (4) 
      -- CP-element group 73: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/R_n_out_count_1837_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/R_n_out_count_1837_sample_completed__ps
      -- CP-element group 73: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/R_n_out_count_1837_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/R_n_out_count_1837_Sample/ack
      -- 
    ack_4478_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_out_count_1909_1837_buf_ack_0, ack => convolve_CP_4290_elements(73)); -- 
    -- CP-element group 74:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	72 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (4) 
      -- CP-element group 74: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/R_n_out_count_1837_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/R_n_out_count_1837_Update/ack
      -- CP-element group 74: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/R_n_out_count_1837_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/R_n_out_count_1837_update_completed__ps
      -- 
    ack_4483_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_out_count_1909_1837_buf_ack_1, ack => convolve_CP_4290_elements(74)); -- 
    -- CP-element group 75:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	14 
    -- CP-element group 75: marked-predecessors 
    -- CP-element group 75: 	78 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/RPIPE_input_pipe1_1840_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/RPIPE_input_pipe1_1840_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/RPIPE_input_pipe1_1840_Sample/rr
      -- 
    rr_4492_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4492_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4290_elements(75), ack => RPIPE_input_pipe1_1840_inst_req_0); -- 
    convolve_cp_element_group_75: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_75"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4290_elements(14) & convolve_CP_4290_elements(78);
      gj_convolve_cp_element_group_75 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4290_elements(75), clk => clk, reset => reset); --
    end block;
    -- CP-element group 76:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	77 
    -- CP-element group 76: 	17 
    -- CP-element group 76: marked-predecessors 
    -- CP-element group 76: 	95 
    -- CP-element group 76: 	99 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	78 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/RPIPE_input_pipe1_1840_update_start_
      -- CP-element group 76: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/RPIPE_input_pipe1_1840_Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/RPIPE_input_pipe1_1840_Update/cr
      -- 
    cr_4497_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4497_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4290_elements(76), ack => RPIPE_input_pipe1_1840_inst_req_1); -- 
    convolve_cp_element_group_76: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 15,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_76"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4290_elements(77) & convolve_CP_4290_elements(17) & convolve_CP_4290_elements(95) & convolve_CP_4290_elements(99);
      gj_convolve_cp_element_group_76 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4290_elements(76), clk => clk, reset => reset); --
    end block;
    -- CP-element group 77:  transition  input  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	76 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/RPIPE_input_pipe1_1840_Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/RPIPE_input_pipe1_1840_sample_completed_
      -- CP-element group 77: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/RPIPE_input_pipe1_1840_Sample/ra
      -- 
    ra_4493_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_pipe1_1840_inst_ack_0, ack => convolve_CP_4290_elements(77)); -- 
    -- CP-element group 78:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	76 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	93 
    -- CP-element group 78: 	97 
    -- CP-element group 78: marked-successors 
    -- CP-element group 78: 	39 
    -- CP-element group 78: 	75 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/RPIPE_input_pipe1_1840_update_completed_
      -- CP-element group 78: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/RPIPE_input_pipe1_1840_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/RPIPE_input_pipe1_1840_Update/ca
      -- 
    ca_4498_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_pipe1_1840_inst_ack_1, ack => convolve_CP_4290_elements(78)); -- 
    -- CP-element group 79:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	14 
    -- CP-element group 79: marked-predecessors 
    -- CP-element group 79: 	82 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	81 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/RPIPE_kernel_pipe1_1847_Sample/rr
      -- CP-element group 79: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/RPIPE_kernel_pipe1_1847_Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/RPIPE_kernel_pipe1_1847_sample_start_
      -- 
    rr_4506_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4506_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4290_elements(79), ack => RPIPE_kernel_pipe1_1847_inst_req_0); -- 
    convolve_cp_element_group_79: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_79"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4290_elements(14) & convolve_CP_4290_elements(82);
      gj_convolve_cp_element_group_79 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4290_elements(79), clk => clk, reset => reset); --
    end block;
    -- CP-element group 80:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	17 
    -- CP-element group 80: 	81 
    -- CP-element group 80: marked-predecessors 
    -- CP-element group 80: 	95 
    -- CP-element group 80: 	99 
    -- CP-element group 80: 	88 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	82 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/RPIPE_kernel_pipe1_1847_Update/$entry
      -- CP-element group 80: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/RPIPE_kernel_pipe1_1847_Update/cr
      -- CP-element group 80: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/RPIPE_kernel_pipe1_1847_update_start_
      -- 
    cr_4511_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4511_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4290_elements(80), ack => RPIPE_kernel_pipe1_1847_inst_req_1); -- 
    convolve_cp_element_group_80: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_80"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_4290_elements(17) & convolve_CP_4290_elements(81) & convolve_CP_4290_elements(95) & convolve_CP_4290_elements(99) & convolve_CP_4290_elements(88);
      gj_convolve_cp_element_group_80 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4290_elements(80), clk => clk, reset => reset); --
    end block;
    -- CP-element group 81:  transition  input  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	79 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	80 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/RPIPE_kernel_pipe1_1847_Sample/$exit
      -- CP-element group 81: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/RPIPE_kernel_pipe1_1847_Sample/ra
      -- CP-element group 81: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/RPIPE_kernel_pipe1_1847_sample_completed_
      -- 
    ra_4507_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_kernel_pipe1_1847_inst_ack_0, ack => convolve_CP_4290_elements(81)); -- 
    -- CP-element group 82:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	80 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	93 
    -- CP-element group 82: 	97 
    -- CP-element group 82: 	87 
    -- CP-element group 82: marked-successors 
    -- CP-element group 82: 	39 
    -- CP-element group 82: 	79 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/RPIPE_kernel_pipe1_1847_Update/$exit
      -- CP-element group 82: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/RPIPE_kernel_pipe1_1847_update_completed_
      -- CP-element group 82: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/RPIPE_kernel_pipe1_1847_Update/ca
      -- 
    ca_4512_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_kernel_pipe1_1847_inst_ack_1, ack => convolve_CP_4290_elements(82)); -- 
    -- CP-element group 83:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	14 
    -- CP-element group 83: marked-predecessors 
    -- CP-element group 83: 	85 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	85 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/SUB_u32_u32_1861_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/SUB_u32_u32_1861_Sample/rr
      -- CP-element group 83: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/SUB_u32_u32_1861_Sample/$entry
      -- 
    rr_4520_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4520_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4290_elements(83), ack => SUB_u32_u32_1861_inst_req_0); -- 
    convolve_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4290_elements(14) & convolve_CP_4290_elements(85);
      gj_convolve_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4290_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	17 
    -- CP-element group 84: marked-predecessors 
    -- CP-element group 84: 	114 
    -- CP-element group 84: 	91 
    -- CP-element group 84: 	103 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/SUB_u32_u32_1861_Update/$entry
      -- CP-element group 84: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/SUB_u32_u32_1861_Update/cr
      -- CP-element group 84: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/SUB_u32_u32_1861_update_start_
      -- 
    cr_4525_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4525_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4290_elements(84), ack => SUB_u32_u32_1861_inst_req_1); -- 
    convolve_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4290_elements(17) & convolve_CP_4290_elements(114) & convolve_CP_4290_elements(91) & convolve_CP_4290_elements(103);
      gj_convolve_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4290_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	83 
    -- CP-element group 85: successors 
    -- CP-element group 85: marked-successors 
    -- CP-element group 85: 	83 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/SUB_u32_u32_1861_sample_completed_
      -- CP-element group 85: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/SUB_u32_u32_1861_Sample/ra
      -- CP-element group 85: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/SUB_u32_u32_1861_Sample/$exit
      -- 
    ra_4521_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u32_u32_1861_inst_ack_0, ack => convolve_CP_4290_elements(85)); -- 
    -- CP-element group 86:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	112 
    -- CP-element group 86: 	90 
    -- CP-element group 86: 	101 
    -- CP-element group 86: marked-successors 
    -- CP-element group 86: 	58 
    -- CP-element group 86: 	39 
    -- CP-element group 86: 	20 
    -- CP-element group 86:  members (3) 
      -- CP-element group 86: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/SUB_u32_u32_1861_update_completed_
      -- CP-element group 86: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/SUB_u32_u32_1861_Update/$exit
      -- CP-element group 86: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/SUB_u32_u32_1861_Update/ca
      -- 
    ca_4526_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u32_u32_1861_inst_ack_1, ack => convolve_CP_4290_elements(86)); -- 
    -- CP-element group 87:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	61 
    -- CP-element group 87: 	82 
    -- CP-element group 87: marked-predecessors 
    -- CP-element group 87: 	89 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (3) 
      -- CP-element group 87: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/WPIPE_kernel_pipe1_1895_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/WPIPE_kernel_pipe1_1895_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/WPIPE_kernel_pipe1_1895_Sample/req
      -- 
    req_4534_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4534_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4290_elements(87), ack => WPIPE_kernel_pipe1_1895_inst_req_0); -- 
    convolve_cp_element_group_87: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_87"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4290_elements(61) & convolve_CP_4290_elements(82) & convolve_CP_4290_elements(89);
      gj_convolve_cp_element_group_87 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4290_elements(87), clk => clk, reset => reset); --
    end block;
    -- CP-element group 88:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	89 
    -- CP-element group 88: marked-successors 
    -- CP-element group 88: 	59 
    -- CP-element group 88: 	80 
    -- CP-element group 88:  members (6) 
      -- CP-element group 88: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/WPIPE_kernel_pipe1_1895_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/WPIPE_kernel_pipe1_1895_Sample/$exit
      -- CP-element group 88: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/WPIPE_kernel_pipe1_1895_Sample/ack
      -- CP-element group 88: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/WPIPE_kernel_pipe1_1895_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/WPIPE_kernel_pipe1_1895_Update/req
      -- CP-element group 88: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/WPIPE_kernel_pipe1_1895_sample_completed_
      -- 
    ack_4535_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe1_1895_inst_ack_0, ack => convolve_CP_4290_elements(88)); -- 
    req_4539_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4539_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4290_elements(88), ack => WPIPE_kernel_pipe1_1895_inst_req_1); -- 
    -- CP-element group 89:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	88 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	124 
    -- CP-element group 89: marked-successors 
    -- CP-element group 89: 	87 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/WPIPE_kernel_pipe1_1895_Update/ack
      -- CP-element group 89: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/WPIPE_kernel_pipe1_1895_Update/$exit
      -- CP-element group 89: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/WPIPE_kernel_pipe1_1895_update_completed_
      -- 
    ack_4540_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe1_1895_inst_ack_1, ack => convolve_CP_4290_elements(89)); -- 
    -- CP-element group 90:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	61 
    -- CP-element group 90: 	25 
    -- CP-element group 90: 	86 
    -- CP-element group 90: marked-predecessors 
    -- CP-element group 90: 	92 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (3) 
      -- CP-element group 90: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/WPIPE_input_done_pipe_1916_Sample/$entry
      -- CP-element group 90: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/WPIPE_input_done_pipe_1916_sample_start_
      -- CP-element group 90: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/WPIPE_input_done_pipe_1916_Sample/req
      -- 
    req_4548_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4548_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4290_elements(90), ack => WPIPE_input_done_pipe_1916_inst_req_0); -- 
    convolve_cp_element_group_90: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_90"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4290_elements(61) & convolve_CP_4290_elements(25) & convolve_CP_4290_elements(86) & convolve_CP_4290_elements(92);
      gj_convolve_cp_element_group_90 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4290_elements(90), clk => clk, reset => reset); --
    end block;
    -- CP-element group 91:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91: marked-successors 
    -- CP-element group 91: 	59 
    -- CP-element group 91: 	21 
    -- CP-element group 91: 	84 
    -- CP-element group 91:  members (6) 
      -- CP-element group 91: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/WPIPE_input_done_pipe_1916_Sample/$exit
      -- CP-element group 91: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/WPIPE_input_done_pipe_1916_Sample/ack
      -- CP-element group 91: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/WPIPE_input_done_pipe_1916_Update/req
      -- CP-element group 91: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/WPIPE_input_done_pipe_1916_sample_completed_
      -- CP-element group 91: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/WPIPE_input_done_pipe_1916_update_start_
      -- CP-element group 91: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/WPIPE_input_done_pipe_1916_Update/$entry
      -- 
    ack_4549_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_done_pipe_1916_inst_ack_0, ack => convolve_CP_4290_elements(91)); -- 
    req_4553_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4553_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4290_elements(91), ack => WPIPE_input_done_pipe_1916_inst_req_1); -- 
    -- CP-element group 92:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	124 
    -- CP-element group 92: marked-successors 
    -- CP-element group 92: 	90 
    -- CP-element group 92:  members (3) 
      -- CP-element group 92: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/WPIPE_input_done_pipe_1916_Update/ack
      -- CP-element group 92: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/WPIPE_input_done_pipe_1916_update_completed_
      -- CP-element group 92: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/WPIPE_input_done_pipe_1916_Update/$exit
      -- 
    ack_4554_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_done_pipe_1916_inst_ack_1, ack => convolve_CP_4290_elements(92)); -- 
    -- CP-element group 93:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	44 
    -- CP-element group 93: 	78 
    -- CP-element group 93: 	82 
    -- CP-element group 93: marked-predecessors 
    -- CP-element group 93: 	95 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/slice_1921_Sample/$entry
      -- CP-element group 93: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/slice_1921_Sample/rr
      -- CP-element group 93: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/slice_1921_sample_start_
      -- 
    rr_4562_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4562_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4290_elements(93), ack => slice_1921_inst_req_0); -- 
    convolve_cp_element_group_93: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_93"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4290_elements(44) & convolve_CP_4290_elements(78) & convolve_CP_4290_elements(82) & convolve_CP_4290_elements(95);
      gj_convolve_cp_element_group_93 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4290_elements(93), clk => clk, reset => reset); --
    end block;
    -- CP-element group 94:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: marked-predecessors 
    -- CP-element group 94: 	107 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	96 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/slice_1921_Update/cr
      -- CP-element group 94: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/slice_1921_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/slice_1921_update_start_
      -- 
    cr_4567_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4567_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4290_elements(94), ack => slice_1921_inst_req_1); -- 
    convolve_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= convolve_CP_4290_elements(107);
      gj_convolve_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4290_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: successors 
    -- CP-element group 95: marked-successors 
    -- CP-element group 95: 	40 
    -- CP-element group 95: 	93 
    -- CP-element group 95: 	76 
    -- CP-element group 95: 	80 
    -- CP-element group 95:  members (3) 
      -- CP-element group 95: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/slice_1921_sample_completed_
      -- CP-element group 95: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/slice_1921_Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/slice_1921_Sample/ra
      -- 
    ra_4563_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_1921_inst_ack_0, ack => convolve_CP_4290_elements(95)); -- 
    -- CP-element group 96:  transition  input  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	94 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	105 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/slice_1921_Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/slice_1921_update_completed_
      -- CP-element group 96: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/slice_1921_Update/ca
      -- 
    ca_4568_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_1921_inst_ack_1, ack => convolve_CP_4290_elements(96)); -- 
    -- CP-element group 97:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	44 
    -- CP-element group 97: 	78 
    -- CP-element group 97: 	82 
    -- CP-element group 97: marked-predecessors 
    -- CP-element group 97: 	99 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	99 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/slice_1925_Sample/$entry
      -- CP-element group 97: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/slice_1925_Sample/rr
      -- CP-element group 97: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/slice_1925_sample_start_
      -- 
    rr_4576_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4576_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4290_elements(97), ack => slice_1925_inst_req_0); -- 
    convolve_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4290_elements(44) & convolve_CP_4290_elements(78) & convolve_CP_4290_elements(82) & convolve_CP_4290_elements(99);
      gj_convolve_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4290_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: marked-predecessors 
    -- CP-element group 98: 	118 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	100 
    -- CP-element group 98:  members (3) 
      -- CP-element group 98: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/slice_1925_update_start_
      -- CP-element group 98: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/slice_1925_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/slice_1925_Update/cr
      -- 
    cr_4581_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4581_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4290_elements(98), ack => slice_1925_inst_req_1); -- 
    convolve_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= convolve_CP_4290_elements(118);
      gj_convolve_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4290_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	97 
    -- CP-element group 99: successors 
    -- CP-element group 99: marked-successors 
    -- CP-element group 99: 	40 
    -- CP-element group 99: 	97 
    -- CP-element group 99: 	76 
    -- CP-element group 99: 	80 
    -- CP-element group 99:  members (3) 
      -- CP-element group 99: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/slice_1925_Sample/$exit
      -- CP-element group 99: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/slice_1925_Sample/ra
      -- CP-element group 99: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/slice_1925_sample_completed_
      -- 
    ra_4577_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_1925_inst_ack_0, ack => convolve_CP_4290_elements(99)); -- 
    -- CP-element group 100:  transition  input  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	98 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	116 
    -- CP-element group 100:  members (3) 
      -- CP-element group 100: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/slice_1925_Update/ca
      -- CP-element group 100: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/slice_1925_Update/$exit
      -- CP-element group 100: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/slice_1925_update_completed_
      -- 
    ca_4582_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_1925_inst_ack_1, ack => convolve_CP_4290_elements(100)); -- 
    -- CP-element group 101:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	25 
    -- CP-element group 101: 	86 
    -- CP-element group 101: marked-predecessors 
    -- CP-element group 101: 	103 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	103 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/assign_stmt_1929_Sample/$entry
      -- CP-element group 101: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/assign_stmt_1929_sample_start_
      -- CP-element group 101: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/assign_stmt_1929_Sample/req
      -- 
    req_4590_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4590_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4290_elements(101), ack => W_next_sum_1903_delayed_1_0_1927_inst_req_0); -- 
    convolve_cp_element_group_101: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_101"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4290_elements(25) & convolve_CP_4290_elements(86) & convolve_CP_4290_elements(103);
      gj_convolve_cp_element_group_101 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4290_elements(101), clk => clk, reset => reset); --
    end block;
    -- CP-element group 102:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: marked-predecessors 
    -- CP-element group 102: 	107 
    -- CP-element group 102: 	110 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	104 
    -- CP-element group 102:  members (3) 
      -- CP-element group 102: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/assign_stmt_1929_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/assign_stmt_1929_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/assign_stmt_1929_Update/req
      -- 
    req_4595_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4595_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4290_elements(102), ack => W_next_sum_1903_delayed_1_0_1927_inst_req_1); -- 
    convolve_cp_element_group_102: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_102"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4290_elements(107) & convolve_CP_4290_elements(110);
      gj_convolve_cp_element_group_102 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4290_elements(102), clk => clk, reset => reset); --
    end block;
    -- CP-element group 103:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	101 
    -- CP-element group 103: successors 
    -- CP-element group 103: marked-successors 
    -- CP-element group 103: 	21 
    -- CP-element group 103: 	84 
    -- CP-element group 103: 	101 
    -- CP-element group 103:  members (3) 
      -- CP-element group 103: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/assign_stmt_1929_Sample/$exit
      -- CP-element group 103: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/assign_stmt_1929_sample_completed_
      -- CP-element group 103: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/assign_stmt_1929_Sample/ack
      -- 
    ack_4591_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_next_sum_1903_delayed_1_0_1927_inst_ack_0, ack => convolve_CP_4290_elements(103)); -- 
    -- CP-element group 104:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	102 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	105 
    -- CP-element group 104: 	109 
    -- CP-element group 104:  members (3) 
      -- CP-element group 104: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/assign_stmt_1929_update_completed_
      -- CP-element group 104: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/assign_stmt_1929_Update/ack
      -- CP-element group 104: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/assign_stmt_1929_Update/$exit
      -- 
    ack_4596_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_next_sum_1903_delayed_1_0_1927_inst_ack_1, ack => convolve_CP_4290_elements(104)); -- 
    -- CP-element group 105:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	96 
    -- CP-element group 105: 	104 
    -- CP-element group 105: marked-predecessors 
    -- CP-element group 105: 	107 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	107 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/type_cast_1933_Sample/rr
      -- CP-element group 105: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/type_cast_1933_Sample/$entry
      -- CP-element group 105: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/type_cast_1933_sample_start_
      -- 
    rr_4604_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4604_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4290_elements(105), ack => type_cast_1933_inst_req_0); -- 
    convolve_cp_element_group_105: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_105"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4290_elements(96) & convolve_CP_4290_elements(104) & convolve_CP_4290_elements(107);
      gj_convolve_cp_element_group_105 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4290_elements(105), clk => clk, reset => reset); --
    end block;
    -- CP-element group 106:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: marked-predecessors 
    -- CP-element group 106: 	110 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	108 
    -- CP-element group 106:  members (3) 
      -- CP-element group 106: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/type_cast_1933_update_start_
      -- CP-element group 106: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/type_cast_1933_Update/$entry
      -- CP-element group 106: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/type_cast_1933_Update/cr
      -- 
    cr_4609_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4609_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4290_elements(106), ack => type_cast_1933_inst_req_1); -- 
    convolve_cp_element_group_106: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_106"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= convolve_CP_4290_elements(110);
      gj_convolve_cp_element_group_106 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4290_elements(106), clk => clk, reset => reset); --
    end block;
    -- CP-element group 107:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	105 
    -- CP-element group 107: successors 
    -- CP-element group 107: marked-successors 
    -- CP-element group 107: 	94 
    -- CP-element group 107: 	102 
    -- CP-element group 107: 	105 
    -- CP-element group 107:  members (3) 
      -- CP-element group 107: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/type_cast_1933_Sample/$exit
      -- CP-element group 107: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/type_cast_1933_Sample/ra
      -- CP-element group 107: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/type_cast_1933_sample_completed_
      -- 
    ra_4605_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1933_inst_ack_0, ack => convolve_CP_4290_elements(107)); -- 
    -- CP-element group 108:  transition  input  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	106 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	109 
    -- CP-element group 108:  members (3) 
      -- CP-element group 108: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/type_cast_1933_update_completed_
      -- CP-element group 108: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/type_cast_1933_Update/$exit
      -- CP-element group 108: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/type_cast_1933_Update/ca
      -- 
    ca_4610_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1933_inst_ack_1, ack => convolve_CP_4290_elements(108)); -- 
    -- CP-element group 109:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	104 
    -- CP-element group 109: 	108 
    -- CP-element group 109: marked-predecessors 
    -- CP-element group 109: 	122 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	110 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/WPIPE_maxpool_output_pipe_1931_sample_start_
      -- CP-element group 109: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/WPIPE_maxpool_output_pipe_1931_Sample/$entry
      -- CP-element group 109: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/WPIPE_maxpool_output_pipe_1931_Sample/req
      -- 
    req_4618_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4618_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4290_elements(109), ack => WPIPE_maxpool_output_pipe_1931_inst_req_0); -- 
    convolve_cp_element_group_109: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_109"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4290_elements(104) & convolve_CP_4290_elements(108) & convolve_CP_4290_elements(122);
      gj_convolve_cp_element_group_109 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4290_elements(109), clk => clk, reset => reset); --
    end block;
    -- CP-element group 110:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	109 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110: marked-successors 
    -- CP-element group 110: 	102 
    -- CP-element group 110: 	106 
    -- CP-element group 110:  members (6) 
      -- CP-element group 110: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/WPIPE_maxpool_output_pipe_1931_sample_completed_
      -- CP-element group 110: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/WPIPE_maxpool_output_pipe_1931_update_start_
      -- CP-element group 110: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/WPIPE_maxpool_output_pipe_1931_Sample/$exit
      -- CP-element group 110: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/WPIPE_maxpool_output_pipe_1931_Sample/ack
      -- CP-element group 110: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/WPIPE_maxpool_output_pipe_1931_Update/$entry
      -- CP-element group 110: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/WPIPE_maxpool_output_pipe_1931_Update/req
      -- 
    ack_4619_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1931_inst_ack_0, ack => convolve_CP_4290_elements(110)); -- 
    req_4623_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4623_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4290_elements(110), ack => WPIPE_maxpool_output_pipe_1931_inst_req_1); -- 
    -- CP-element group 111:  transition  input  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	120 
    -- CP-element group 111:  members (3) 
      -- CP-element group 111: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/WPIPE_maxpool_output_pipe_1931_update_completed_
      -- CP-element group 111: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/WPIPE_maxpool_output_pipe_1931_Update/$exit
      -- CP-element group 111: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/WPIPE_maxpool_output_pipe_1931_Update/ack
      -- 
    ack_4624_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1931_inst_ack_1, ack => convolve_CP_4290_elements(111)); -- 
    -- CP-element group 112:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	25 
    -- CP-element group 112: 	86 
    -- CP-element group 112: marked-predecessors 
    -- CP-element group 112: 	114 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	114 
    -- CP-element group 112:  members (3) 
      -- CP-element group 112: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/assign_stmt_1937_sample_start_
      -- CP-element group 112: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/assign_stmt_1937_Sample/$entry
      -- CP-element group 112: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/assign_stmt_1937_Sample/req
      -- 
    req_4632_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4632_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4290_elements(112), ack => W_next_sum_1908_delayed_1_0_1935_inst_req_0); -- 
    convolve_cp_element_group_112: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_112"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4290_elements(25) & convolve_CP_4290_elements(86) & convolve_CP_4290_elements(114);
      gj_convolve_cp_element_group_112 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4290_elements(112), clk => clk, reset => reset); --
    end block;
    -- CP-element group 113:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: marked-predecessors 
    -- CP-element group 113: 	118 
    -- CP-element group 113: 	121 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/assign_stmt_1937_update_start_
      -- CP-element group 113: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/assign_stmt_1937_Update/$entry
      -- CP-element group 113: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/assign_stmt_1937_Update/req
      -- 
    req_4637_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4637_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4290_elements(113), ack => W_next_sum_1908_delayed_1_0_1935_inst_req_1); -- 
    convolve_cp_element_group_113: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_113"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4290_elements(118) & convolve_CP_4290_elements(121);
      gj_convolve_cp_element_group_113 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4290_elements(113), clk => clk, reset => reset); --
    end block;
    -- CP-element group 114:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	112 
    -- CP-element group 114: successors 
    -- CP-element group 114: marked-successors 
    -- CP-element group 114: 	112 
    -- CP-element group 114: 	21 
    -- CP-element group 114: 	84 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/assign_stmt_1937_sample_completed_
      -- CP-element group 114: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/assign_stmt_1937_Sample/$exit
      -- CP-element group 114: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/assign_stmt_1937_Sample/ack
      -- 
    ack_4633_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_next_sum_1908_delayed_1_0_1935_inst_ack_0, ack => convolve_CP_4290_elements(114)); -- 
    -- CP-element group 115:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	116 
    -- CP-element group 115: 	120 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/assign_stmt_1937_update_completed_
      -- CP-element group 115: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/assign_stmt_1937_Update/$exit
      -- CP-element group 115: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/assign_stmt_1937_Update/ack
      -- 
    ack_4638_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_next_sum_1908_delayed_1_0_1935_inst_ack_1, ack => convolve_CP_4290_elements(115)); -- 
    -- CP-element group 116:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	115 
    -- CP-element group 116: 	100 
    -- CP-element group 116: marked-predecessors 
    -- CP-element group 116: 	118 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	118 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/type_cast_1941_sample_start_
      -- CP-element group 116: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/type_cast_1941_Sample/$entry
      -- CP-element group 116: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/type_cast_1941_Sample/rr
      -- 
    rr_4646_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4646_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4290_elements(116), ack => type_cast_1941_inst_req_0); -- 
    convolve_cp_element_group_116: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_116"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4290_elements(115) & convolve_CP_4290_elements(100) & convolve_CP_4290_elements(118);
      gj_convolve_cp_element_group_116 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4290_elements(116), clk => clk, reset => reset); --
    end block;
    -- CP-element group 117:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: marked-predecessors 
    -- CP-element group 117: 	121 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	119 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/type_cast_1941_update_start_
      -- CP-element group 117: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/type_cast_1941_Update/$entry
      -- CP-element group 117: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/type_cast_1941_Update/cr
      -- 
    cr_4651_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4651_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4290_elements(117), ack => type_cast_1941_inst_req_1); -- 
    convolve_cp_element_group_117: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_117"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= convolve_CP_4290_elements(121);
      gj_convolve_cp_element_group_117 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4290_elements(117), clk => clk, reset => reset); --
    end block;
    -- CP-element group 118:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	116 
    -- CP-element group 118: successors 
    -- CP-element group 118: marked-successors 
    -- CP-element group 118: 	113 
    -- CP-element group 118: 	116 
    -- CP-element group 118: 	98 
    -- CP-element group 118:  members (3) 
      -- CP-element group 118: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/type_cast_1941_sample_completed_
      -- CP-element group 118: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/type_cast_1941_Sample/$exit
      -- CP-element group 118: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/type_cast_1941_Sample/ra
      -- 
    ra_4647_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1941_inst_ack_0, ack => convolve_CP_4290_elements(118)); -- 
    -- CP-element group 119:  transition  input  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	117 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	120 
    -- CP-element group 119:  members (3) 
      -- CP-element group 119: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/type_cast_1941_update_completed_
      -- CP-element group 119: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/type_cast_1941_Update/$exit
      -- CP-element group 119: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/type_cast_1941_Update/ca
      -- 
    ca_4652_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1941_inst_ack_1, ack => convolve_CP_4290_elements(119)); -- 
    -- CP-element group 120:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	111 
    -- CP-element group 120: 	115 
    -- CP-element group 120: 	119 
    -- CP-element group 120: marked-predecessors 
    -- CP-element group 120: 	122 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120:  members (3) 
      -- CP-element group 120: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/WPIPE_maxpool_output_pipe_1939_sample_start_
      -- CP-element group 120: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/WPIPE_maxpool_output_pipe_1939_Sample/$entry
      -- CP-element group 120: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/WPIPE_maxpool_output_pipe_1939_Sample/req
      -- 
    req_4660_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4660_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4290_elements(120), ack => WPIPE_maxpool_output_pipe_1939_inst_req_0); -- 
    convolve_cp_element_group_120: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_120"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4290_elements(111) & convolve_CP_4290_elements(115) & convolve_CP_4290_elements(119) & convolve_CP_4290_elements(122);
      gj_convolve_cp_element_group_120 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4290_elements(120), clk => clk, reset => reset); --
    end block;
    -- CP-element group 121:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121: marked-successors 
    -- CP-element group 121: 	113 
    -- CP-element group 121: 	117 
    -- CP-element group 121:  members (6) 
      -- CP-element group 121: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/WPIPE_maxpool_output_pipe_1939_sample_completed_
      -- CP-element group 121: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/WPIPE_maxpool_output_pipe_1939_update_start_
      -- CP-element group 121: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/WPIPE_maxpool_output_pipe_1939_Sample/$exit
      -- CP-element group 121: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/WPIPE_maxpool_output_pipe_1939_Sample/ack
      -- CP-element group 121: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/WPIPE_maxpool_output_pipe_1939_Update/$entry
      -- CP-element group 121: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/WPIPE_maxpool_output_pipe_1939_Update/req
      -- 
    ack_4661_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1939_inst_ack_0, ack => convolve_CP_4290_elements(121)); -- 
    req_4665_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4665_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4290_elements(121), ack => WPIPE_maxpool_output_pipe_1939_inst_req_1); -- 
    -- CP-element group 122:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	124 
    -- CP-element group 122: marked-successors 
    -- CP-element group 122: 	120 
    -- CP-element group 122: 	109 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/WPIPE_maxpool_output_pipe_1939_update_completed_
      -- CP-element group 122: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/WPIPE_maxpool_output_pipe_1939_Update/$exit
      -- CP-element group 122: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/WPIPE_maxpool_output_pipe_1939_Update/ack
      -- 
    ack_4666_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1939_inst_ack_1, ack => convolve_CP_4290_elements(122)); -- 
    -- CP-element group 123:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	14 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	15 
    -- CP-element group 123:  members (1) 
      -- CP-element group 123: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group convolve_CP_4290_elements(123) is a control-delay.
    cp_element_123_delay: control_delay_element  generic map(name => " 123_delay", delay_value => 1)  port map(req => convolve_CP_4290_elements(14), ack => convolve_CP_4290_elements(123), clk => clk, reset =>reset);
    -- CP-element group 124:  join  transition  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	122 
    -- CP-element group 124: 	92 
    -- CP-element group 124: 	89 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	11 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_1807/do_while_stmt_1823/do_while_stmt_1823_loop_body/$exit
      -- 
    convolve_cp_element_group_124: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_124"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4290_elements(122) & convolve_CP_4290_elements(92) & convolve_CP_4290_elements(89);
      gj_convolve_cp_element_group_124 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4290_elements(124), clk => clk, reset => reset); --
    end block;
    -- CP-element group 125:  transition  input  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	10 
    -- CP-element group 125: successors 
    -- CP-element group 125:  members (2) 
      -- CP-element group 125: 	 branch_block_stmt_1807/do_while_stmt_1823/loop_exit/$exit
      -- CP-element group 125: 	 branch_block_stmt_1807/do_while_stmt_1823/loop_exit/ack
      -- 
    ack_4671_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1823_branch_ack_0, ack => convolve_CP_4290_elements(125)); -- 
    -- CP-element group 126:  transition  input  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	10 
    -- CP-element group 126: successors 
    -- CP-element group 126:  members (2) 
      -- CP-element group 126: 	 branch_block_stmt_1807/do_while_stmt_1823/loop_taken/$exit
      -- CP-element group 126: 	 branch_block_stmt_1807/do_while_stmt_1823/loop_taken/ack
      -- 
    ack_4675_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1823_branch_ack_1, ack => convolve_CP_4290_elements(126)); -- 
    -- CP-element group 127:  transition  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	8 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	1 
    -- CP-element group 127:  members (1) 
      -- CP-element group 127: 	 branch_block_stmt_1807/do_while_stmt_1823/$exit
      -- 
    convolve_CP_4290_elements(127) <= convolve_CP_4290_elements(8);
    convolve_do_while_stmt_1823_terminator_4676: loop_terminator -- 
      generic map (name => " convolve_do_while_stmt_1823_terminator_4676", max_iterations_in_flight =>15) 
      port map(loop_body_exit => convolve_CP_4290_elements(11),loop_continue => convolve_CP_4290_elements(126),loop_terminate => convolve_CP_4290_elements(125),loop_back => convolve_CP_4290_elements(9),loop_exit => convolve_CP_4290_elements(8),clk => clk, reset => reset); -- 
    phi_stmt_1825_phi_seq_4396_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convolve_CP_4290_elements(28);
      convolve_CP_4290_elements(31)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convolve_CP_4290_elements(31);
      convolve_CP_4290_elements(32)<= src_update_reqs(0);
      src_update_acks(0)  <= convolve_CP_4290_elements(33);
      convolve_CP_4290_elements(29) <= phi_mux_reqs(0);
      triggers(1)  <= convolve_CP_4290_elements(26);
      convolve_CP_4290_elements(35)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convolve_CP_4290_elements(37);
      convolve_CP_4290_elements(36)<= src_update_reqs(1);
      src_update_acks(1)  <= convolve_CP_4290_elements(38);
      convolve_CP_4290_elements(27) <= phi_mux_reqs(1);
      phi_stmt_1825_phi_seq_4396 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1825_phi_seq_4396") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convolve_CP_4290_elements(22), 
          phi_sample_ack => convolve_CP_4290_elements(23), 
          phi_update_req => convolve_CP_4290_elements(24), 
          phi_update_ack => convolve_CP_4290_elements(25), 
          phi_mux_ack => convolve_CP_4290_elements(30), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1829_phi_seq_4440_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convolve_CP_4290_elements(45);
      convolve_CP_4290_elements(50)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convolve_CP_4290_elements(52);
      convolve_CP_4290_elements(51)<= src_update_reqs(0);
      src_update_acks(0)  <= convolve_CP_4290_elements(53);
      convolve_CP_4290_elements(46) <= phi_mux_reqs(0);
      triggers(1)  <= convolve_CP_4290_elements(47);
      convolve_CP_4290_elements(54)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convolve_CP_4290_elements(54);
      convolve_CP_4290_elements(55)<= src_update_reqs(1);
      src_update_acks(1)  <= convolve_CP_4290_elements(56);
      convolve_CP_4290_elements(48) <= phi_mux_reqs(1);
      phi_stmt_1829_phi_seq_4440 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1829_phi_seq_4440") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convolve_CP_4290_elements(41), 
          phi_sample_ack => convolve_CP_4290_elements(42), 
          phi_update_req => convolve_CP_4290_elements(43), 
          phi_update_ack => convolve_CP_4290_elements(44), 
          phi_mux_ack => convolve_CP_4290_elements(49), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1833_phi_seq_4484_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convolve_CP_4290_elements(64);
      convolve_CP_4290_elements(67)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convolve_CP_4290_elements(67);
      convolve_CP_4290_elements(68)<= src_update_reqs(0);
      src_update_acks(0)  <= convolve_CP_4290_elements(69);
      convolve_CP_4290_elements(65) <= phi_mux_reqs(0);
      triggers(1)  <= convolve_CP_4290_elements(62);
      convolve_CP_4290_elements(71)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convolve_CP_4290_elements(73);
      convolve_CP_4290_elements(72)<= src_update_reqs(1);
      src_update_acks(1)  <= convolve_CP_4290_elements(74);
      convolve_CP_4290_elements(63) <= phi_mux_reqs(1);
      phi_stmt_1833_phi_seq_4484 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1833_phi_seq_4484") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convolve_CP_4290_elements(16), 
          phi_sample_ack => convolve_CP_4290_elements(60), 
          phi_update_req => convolve_CP_4290_elements(18), 
          phi_update_ack => convolve_CP_4290_elements(61), 
          phi_mux_ack => convolve_CP_4290_elements(66), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_4348_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= convolve_CP_4290_elements(12);
        preds(1)  <= convolve_CP_4290_elements(13);
        entry_tmerge_4348 : transition_merge -- 
          generic map(name => " entry_tmerge_4348")
          port map (preds => preds, symbol_out => convolve_CP_4290_elements(14));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u16_u16_1905_wire : std_logic_vector(15 downto 0);
    signal ADD_u32_u32_1886_wire : std_logic_vector(31 downto 0);
    signal MUX_1906_wire : std_logic_vector(15 downto 0);
    signal SUB_u32_u32_1841_1841_delayed_1_0_1862 : std_logic_vector(31 downto 0);
    signal acc_1829 : std_logic_vector(15 downto 0);
    signal acc_val_1874 : std_logic_vector(15 downto 0);
    signal acc_val_dn_1926 : std_logic_vector(7 downto 0);
    signal acc_val_up_1922 : std_logic_vector(7 downto 0);
    signal acc_var_1822 : std_logic_vector(15 downto 0);
    signal all_done_flag_1914 : std_logic_vector(0 downto 0);
    signal iread_1841 : std_logic_vector(15 downto 0);
    signal ival_1845 : std_logic_vector(15 downto 0);
    signal konst_1860_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1877_wire_constant : std_logic_vector(15 downto 0);
    signal konst_1883_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1885_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1904_wire_constant : std_logic_vector(15 downto 0);
    signal konst_1917_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1944_wire_constant : std_logic_vector(0 downto 0);
    signal kread_1848 : std_logic_vector(15 downto 0);
    signal kval_1852 : std_logic_vector(15 downto 0);
    signal mcount_var_1817 : std_logic_vector(31 downto 0);
    signal mul_val_1857 : std_logic_vector(15 downto 0);
    signal mycount_1825 : std_logic_vector(31 downto 0);
    signal n_out_count_1909 : std_logic_vector(15 downto 0);
    signal n_out_count_1909_1837_buffered : std_logic_vector(15 downto 0);
    signal nacc_1880 : std_logic_vector(15 downto 0);
    signal nacc_1880_1831_buffered : std_logic_vector(15 downto 0);
    signal next_sum_1867 : std_logic_vector(0 downto 0);
    signal next_sum_1903_delayed_1_0_1929 : std_logic_vector(0 downto 0);
    signal next_sum_1908_delayed_1_0_1937 : std_logic_vector(0 downto 0);
    signal nmycount_1888 : std_logic_vector(31 downto 0);
    signal nmycount_1888_1828_buffered : std_logic_vector(31 downto 0);
    signal num_out_1810 : std_logic_vector(15 downto 0);
    signal out_count_1833 : std_logic_vector(15 downto 0);
    signal out_done_flag_1893 : std_logic_vector(0 downto 0);
    signal size_1813 : std_logic_vector(31 downto 0);
    signal type_cast_1836_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1870_wire : std_logic_vector(15 downto 0);
    signal type_cast_1872_wire : std_logic_vector(15 downto 0);
    signal type_cast_1902_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1933_wire : std_logic_vector(7 downto 0);
    signal type_cast_1941_wire : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    acc_var_1822 <= "0000000000000000";
    konst_1860_wire_constant <= "00000000000000000000000000000001";
    konst_1877_wire_constant <= "0000000000000000";
    konst_1883_wire_constant <= "00000000000000000000000000000000";
    konst_1885_wire_constant <= "00000000000000000000000000000001";
    konst_1904_wire_constant <= "0000000000000001";
    konst_1917_wire_constant <= "1";
    konst_1944_wire_constant <= "1";
    mcount_var_1817 <= "00000000000000000000000000000000";
    type_cast_1836_wire_constant <= "0000000000000001";
    type_cast_1902_wire_constant <= "0000000000000001";
    phi_stmt_1825: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= mcount_var_1817 & nmycount_1888_1828_buffered;
      req <= phi_stmt_1825_req_0 & phi_stmt_1825_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1825",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1825_ack_0,
          idata => idata,
          odata => mycount_1825,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1825
    phi_stmt_1829: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= nacc_1880_1831_buffered & acc_var_1822;
      req <= phi_stmt_1829_req_0 & phi_stmt_1829_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1829",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1829_ack_0,
          idata => idata,
          odata => acc_1829,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1829
    phi_stmt_1833: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1836_wire_constant & n_out_count_1909_1837_buffered;
      req <= phi_stmt_1833_req_0 & phi_stmt_1833_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1833",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1833_ack_0,
          idata => idata,
          odata => out_count_1833,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1833
    -- flow-through select operator MUX_1879_inst
    nacc_1880 <= konst_1877_wire_constant when (next_sum_1867(0) /=  '0') else acc_val_1874;
    -- flow-through select operator MUX_1887_inst
    nmycount_1888 <= konst_1883_wire_constant when (next_sum_1867(0) /=  '0') else ADD_u32_u32_1886_wire;
    -- flow-through select operator MUX_1906_inst
    MUX_1906_wire <= type_cast_1902_wire_constant when (out_done_flag_1893(0) /=  '0') else ADD_u16_u16_1905_wire;
    -- flow-through select operator MUX_1908_inst
    n_out_count_1909 <= MUX_1906_wire when (next_sum_1867(0) /=  '0') else out_count_1833;
    slice_1921_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_1921_inst_req_0;
      slice_1921_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_1921_inst_req_1;
      slice_1921_inst_ack_1<= update_ack(0);
      slice_1921_inst: SliceSplitProtocol generic map(name => "slice_1921_inst", in_data_width => 16, high_index => 15, low_index => 8, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => acc_val_1874, dout => acc_val_up_1922, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_1925_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_1925_inst_req_0;
      slice_1925_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_1925_inst_req_1;
      slice_1925_inst_ack_1<= update_ack(0);
      slice_1925_inst: SliceSplitProtocol generic map(name => "slice_1925_inst", in_data_width => 16, high_index => 7, low_index => 0, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => acc_val_1874, dout => acc_val_dn_1926, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    W_next_sum_1903_delayed_1_0_1927_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_next_sum_1903_delayed_1_0_1927_inst_req_0;
      W_next_sum_1903_delayed_1_0_1927_inst_ack_0<= wack(0);
      rreq(0) <= W_next_sum_1903_delayed_1_0_1927_inst_req_1;
      W_next_sum_1903_delayed_1_0_1927_inst_ack_1<= rack(0);
      W_next_sum_1903_delayed_1_0_1927_inst : InterlockBuffer generic map ( -- 
        name => "W_next_sum_1903_delayed_1_0_1927_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_sum_1867,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_sum_1903_delayed_1_0_1929,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_next_sum_1908_delayed_1_0_1935_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_next_sum_1908_delayed_1_0_1935_inst_req_0;
      W_next_sum_1908_delayed_1_0_1935_inst_ack_0<= wack(0);
      rreq(0) <= W_next_sum_1908_delayed_1_0_1935_inst_req_1;
      W_next_sum_1908_delayed_1_0_1935_inst_ack_1<= rack(0);
      W_next_sum_1908_delayed_1_0_1935_inst : InterlockBuffer generic map ( -- 
        name => "W_next_sum_1908_delayed_1_0_1935_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_sum_1867,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_sum_1908_delayed_1_0_1937,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_out_count_1909_1837_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_out_count_1909_1837_buf_req_0;
      n_out_count_1909_1837_buf_ack_0<= wack(0);
      rreq(0) <= n_out_count_1909_1837_buf_req_1;
      n_out_count_1909_1837_buf_ack_1<= rack(0);
      n_out_count_1909_1837_buf : InterlockBuffer generic map ( -- 
        name => "n_out_count_1909_1837_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_out_count_1909,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_out_count_1909_1837_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nacc_1880_1831_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nacc_1880_1831_buf_req_0;
      nacc_1880_1831_buf_ack_0<= wack(0);
      rreq(0) <= nacc_1880_1831_buf_req_1;
      nacc_1880_1831_buf_ack_1<= rack(0);
      nacc_1880_1831_buf : InterlockBuffer generic map ( -- 
        name => "nacc_1880_1831_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nacc_1880,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nacc_1880_1831_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nmycount_1888_1828_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nmycount_1888_1828_buf_req_0;
      nmycount_1888_1828_buf_ack_0<= wack(0);
      rreq(0) <= nmycount_1888_1828_buf_req_1;
      nmycount_1888_1828_buf_ack_1<= rack(0);
      nmycount_1888_1828_buf : InterlockBuffer generic map ( -- 
        name => "nmycount_1888_1828_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nmycount_1888,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nmycount_1888_1828_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1844_inst
    process(iread_1841) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := iread_1841(15 downto 0);
      ival_1845 <= tmp_var; -- 
    end process;
    -- interlock type_cast_1851_inst
    process(kread_1848) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := kread_1848(15 downto 0);
      kval_1852 <= tmp_var; -- 
    end process;
    -- interlock type_cast_1870_inst
    process(acc_1829) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := acc_1829(15 downto 0);
      type_cast_1870_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1872_inst
    process(mul_val_1857) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := mul_val_1857(15 downto 0);
      type_cast_1872_wire <= tmp_var; -- 
    end process;
    type_cast_1933_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_1933_inst_req_0;
      type_cast_1933_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_1933_inst_req_1;
      type_cast_1933_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  next_sum_1903_delayed_1_0_1929(0);
      type_cast_1933_inst_gI: SplitGuardInterface generic map(name => "type_cast_1933_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_1933_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1933_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => acc_val_up_1922,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1933_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1941_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_1941_inst_req_0;
      type_cast_1941_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_1941_inst_req_1;
      type_cast_1941_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  next_sum_1908_delayed_1_0_1937(0);
      type_cast_1941_inst_gI: SplitGuardInterface generic map(name => "type_cast_1941_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_1941_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1941_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => acc_val_dn_1926,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1941_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    do_while_stmt_1823_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_1944_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1823_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1823_branch_req_0,
          ack0 => do_while_stmt_1823_branch_ack_0,
          ack1 => do_while_stmt_1823_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_i16_i16_1873_inst
    process(type_cast_1870_wire, type_cast_1872_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(type_cast_1870_wire, type_cast_1872_wire, tmp_var);
      acc_val_1874 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1905_inst
    process(out_count_1833) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(out_count_1833, konst_1904_wire_constant, tmp_var);
      ADD_u16_u16_1905_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1886_inst
    process(mycount_1825) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mycount_1825, konst_1885_wire_constant, tmp_var);
      ADD_u32_u32_1886_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1913_inst
    process(out_done_flag_1893, next_sum_1867) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(out_done_flag_1893, next_sum_1867, tmp_var);
      all_done_flag_1914 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_1892_inst
    process(out_count_1833, num_out_1810) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(out_count_1833, num_out_1810, tmp_var);
      out_done_flag_1893 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1866_inst
    process(mycount_1825, SUB_u32_u32_1841_1841_delayed_1_0_1862) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(mycount_1825, SUB_u32_u32_1841_1841_delayed_1_0_1862, tmp_var);
      next_sum_1867 <= tmp_var; --
    end process;
    -- binary operator MUL_i16_i16_1856_inst
    process(kval_1852, ival_1845) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval_1852, ival_1845, tmp_var);
      mul_val_1857 <= tmp_var; --
    end process;
    -- shared split operator group (7) : SUB_u32_u32_1861_inst 
    ApIntSub_group_7: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= size_1813;
      SUB_u32_u32_1841_1841_delayed_1_0_1862 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u32_u32_1861_inst_req_0;
      SUB_u32_u32_1861_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u32_u32_1861_inst_req_1;
      SUB_u32_u32_1861_inst_ack_1 <= ackR_unguarded(0);
      ApIntSub_group_7_gI: SplitGuardInterface generic map(name => "ApIntSub_group_7_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_7",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- shared inport operator group (0) : RPIPE_input_pipe1_1840_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_input_pipe1_1840_inst_req_0;
      RPIPE_input_pipe1_1840_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_input_pipe1_1840_inst_req_1;
      RPIPE_input_pipe1_1840_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      iread_1841 <= data_out(15 downto 0);
      input_pipe1_read_0_gI: SplitGuardInterface generic map(name => "input_pipe1_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      input_pipe1_read_0: InputPortRevised -- 
        generic map ( name => "input_pipe1_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => input_pipe1_pipe_read_req(0),
          oack => input_pipe1_pipe_read_ack(0),
          odata => input_pipe1_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_kernel_pipe1_1847_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_kernel_pipe1_1847_inst_req_0;
      RPIPE_kernel_pipe1_1847_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_kernel_pipe1_1847_inst_req_1;
      RPIPE_kernel_pipe1_1847_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      kread_1848 <= data_out(15 downto 0);
      kernel_pipe1_read_1_gI: SplitGuardInterface generic map(name => "kernel_pipe1_read_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      kernel_pipe1_read_1: InputPortRevised -- 
        generic map ( name => "kernel_pipe1_read_1", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => kernel_pipe1_pipe_read_req(0),
          oack => kernel_pipe1_pipe_read_ack(0),
          odata => kernel_pipe1_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : RPIPE_num_out_pipe_1809_inst 
    InportGroup_2: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_num_out_pipe_1809_inst_req_0;
      RPIPE_num_out_pipe_1809_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_num_out_pipe_1809_inst_req_1;
      RPIPE_num_out_pipe_1809_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      num_out_1810 <= data_out(15 downto 0);
      num_out_pipe_read_2_gI: SplitGuardInterface generic map(name => "num_out_pipe_read_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      num_out_pipe_read_2: InputPortRevised -- 
        generic map ( name => "num_out_pipe_read_2", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => num_out_pipe_pipe_read_req(0),
          oack => num_out_pipe_pipe_read_ack(0),
          odata => num_out_pipe_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : RPIPE_size_pipe_1812_inst 
    InportGroup_3: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_size_pipe_1812_inst_req_0;
      RPIPE_size_pipe_1812_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_size_pipe_1812_inst_req_1;
      RPIPE_size_pipe_1812_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      size_1813 <= data_out(31 downto 0);
      size_pipe_read_3_gI: SplitGuardInterface generic map(name => "size_pipe_read_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      size_pipe_read_3: InputPortRevised -- 
        generic map ( name => "size_pipe_read_3", data_width => 32,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => size_pipe_pipe_read_req(0),
          oack => size_pipe_pipe_read_ack(0),
          odata => size_pipe_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- shared outport operator group (0) : WPIPE_input_done_pipe_1916_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_input_done_pipe_1916_inst_req_0;
      WPIPE_input_done_pipe_1916_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_input_done_pipe_1916_inst_req_1;
      WPIPE_input_done_pipe_1916_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= all_done_flag_1914(0);
      data_in <= konst_1917_wire_constant;
      input_done_pipe_write_0_gI: SplitGuardInterface generic map(name => "input_done_pipe_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      input_done_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "input_done_pipe", data_width => 1, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => input_done_pipe_pipe_write_req(0),
          oack => input_done_pipe_pipe_write_ack(0),
          odata => input_done_pipe_pipe_write_data(0 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_kernel_pipe1_1895_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_kernel_pipe1_1895_inst_req_0;
      WPIPE_kernel_pipe1_1895_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_kernel_pipe1_1895_inst_req_1;
      WPIPE_kernel_pipe1_1895_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  not out_done_flag_1893(0);
      data_in <= kread_1848;
      kernel_pipe1_write_1_gI: SplitGuardInterface generic map(name => "kernel_pipe1_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      kernel_pipe1_write_1: OutputPortRevised -- 
        generic map ( name => "kernel_pipe1", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => kernel_pipe1_pipe_write_req(0),
          oack => kernel_pipe1_pipe_write_ack(0),
          odata => kernel_pipe1_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_maxpool_output_pipe_1931_inst WPIPE_maxpool_output_pipe_1939_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 1 downto 0);
      signal update_req, update_ack : BooleanArray( 1 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 1 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => true, 1 => true);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      sample_req_unguarded(1) <= WPIPE_maxpool_output_pipe_1931_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_maxpool_output_pipe_1939_inst_req_0;
      WPIPE_maxpool_output_pipe_1931_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_maxpool_output_pipe_1939_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(1) <= WPIPE_maxpool_output_pipe_1931_inst_req_1;
      update_req_unguarded(0) <= WPIPE_maxpool_output_pipe_1939_inst_req_1;
      WPIPE_maxpool_output_pipe_1931_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_maxpool_output_pipe_1939_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= next_sum_1908_delayed_1_0_1937(0);
      guard_vector(1)  <= next_sum_1903_delayed_1_0_1929(0);
      data_in <= type_cast_1933_wire & type_cast_1941_wire;
      maxpool_output_pipe_write_2_gI: SplitGuardInterface generic map(name => "maxpool_output_pipe_write_2_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      maxpool_output_pipe_write_2: OutputPortRevised -- 
        generic map ( name => "maxpool_output_pipe", data_width => 8, num_reqs => 2, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => maxpool_output_pipe_pipe_write_req(0),
          oack => maxpool_output_pipe_pipe_write_ack(0),
          odata => maxpool_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- 
  end Block; -- data_path
  -- 
end convolve_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity loadKernelChannel is -- 
  generic (tag_length : integer); 
  port ( -- 
    start_add : in  std_logic_vector(63 downto 0);
    end_add : in  std_logic_vector(63 downto 0);
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
    input_done_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    input_done_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    input_done_pipe_pipe_read_data : in   std_logic_vector(0 downto 0);
    size_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    size_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    size_pipe_pipe_write_data : out  std_logic_vector(31 downto 0);
    kernel_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity loadKernelChannel;
architecture loadKernelChannel_arch of loadKernelChannel is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 128)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal start_add_buffer :  std_logic_vector(63 downto 0);
  signal start_add_update_enable: Boolean;
  signal end_add_buffer :  std_logic_vector(63 downto 0);
  signal end_add_update_enable: Boolean;
  -- output port buffer signals
  signal loadKernelChannel_CP_676_start: Boolean;
  signal loadKernelChannel_CP_676_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal nfetch_val_419_358_buf_req_1 : boolean;
  signal addr_of_398_final_reg_ack_0 : boolean;
  signal do_while_stmt_350_branch_ack_0 : boolean;
  signal nfetch_val_419_358_buf_ack_1 : boolean;
  signal my_fetch_339_359_buf_ack_0 : boolean;
  signal type_cast_432_inst_ack_1 : boolean;
  signal array_obj_ref_397_index_offset_ack_0 : boolean;
  signal addr_of_398_final_reg_req_1 : boolean;
  signal ptr_deref_406_load_0_req_0 : boolean;
  signal addr_of_398_final_reg_ack_1 : boolean;
  signal W_fn_394_delayed_13_0_408_inst_req_0 : boolean;
  signal phi_stmt_356_ack_0 : boolean;
  signal W_fn_394_delayed_13_0_408_inst_ack_0 : boolean;
  signal phi_stmt_356_req_1 : boolean;
  signal array_obj_ref_397_index_offset_req_1 : boolean;
  signal ptr_deref_406_load_0_req_1 : boolean;
  signal WPIPE_size_pipe_428_inst_req_0 : boolean;
  signal ptr_deref_406_load_0_ack_0 : boolean;
  signal array_obj_ref_397_index_offset_req_0 : boolean;
  signal W_fn_394_delayed_13_0_408_inst_req_1 : boolean;
  signal W_fn_394_delayed_13_0_408_inst_ack_1 : boolean;
  signal W_fn_388_delayed_7_0_400_inst_req_0 : boolean;
  signal WPIPE_size_pipe_428_inst_ack_0 : boolean;
  signal W_fn_388_delayed_7_0_400_inst_ack_0 : boolean;
  signal array_obj_ref_397_index_offset_ack_1 : boolean;
  signal my_fetch_339_359_buf_req_0 : boolean;
  signal WPIPE_kernel_pipe1_381_inst_ack_0 : boolean;
  signal WPIPE_kernel_pipe1_381_inst_ack_1 : boolean;
  signal W_fn_388_delayed_7_0_400_inst_req_1 : boolean;
  signal W_fetch_val_396_delayed_13_0_411_inst_ack_0 : boolean;
  signal W_fetch_val_396_delayed_13_0_411_inst_req_0 : boolean;
  signal W_fn_388_delayed_7_0_400_inst_ack_1 : boolean;
  signal do_while_stmt_350_branch_ack_1 : boolean;
  signal addr_of_398_final_reg_req_0 : boolean;
  signal WPIPE_kernel_pipe1_381_inst_req_1 : boolean;
  signal phi_stmt_356_req_0 : boolean;
  signal type_cast_432_inst_ack_0 : boolean;
  signal type_cast_432_inst_req_0 : boolean;
  signal my_fetch_339_359_buf_req_1 : boolean;
  signal type_cast_432_inst_req_1 : boolean;
  signal ptr_deref_406_load_0_ack_1 : boolean;
  signal WPIPE_size_pipe_428_inst_req_1 : boolean;
  signal WPIPE_kernel_pipe1_381_inst_req_0 : boolean;
  signal my_fetch_339_359_buf_ack_1 : boolean;
  signal WPIPE_size_pipe_428_inst_ack_1 : boolean;
  signal nfetch_val_419_358_buf_req_0 : boolean;
  signal array_obj_ref_333_index_offset_req_0 : boolean;
  signal array_obj_ref_333_index_offset_ack_0 : boolean;
  signal array_obj_ref_333_index_offset_req_1 : boolean;
  signal array_obj_ref_333_index_offset_ack_1 : boolean;
  signal W_fetch_val_396_delayed_13_0_411_inst_ack_1 : boolean;
  signal addr_of_334_final_reg_req_0 : boolean;
  signal W_fetch_val_396_delayed_13_0_411_inst_req_1 : boolean;
  signal addr_of_334_final_reg_ack_0 : boolean;
  signal addr_of_334_final_reg_req_1 : boolean;
  signal addr_of_334_final_reg_ack_1 : boolean;
  signal ptr_deref_338_load_0_req_0 : boolean;
  signal ptr_deref_338_load_0_ack_0 : boolean;
  signal start_add_355_buf_ack_1 : boolean;
  signal nfetch_val_419_358_buf_ack_0 : boolean;
  signal ptr_deref_338_load_0_req_1 : boolean;
  signal ptr_deref_338_load_0_ack_1 : boolean;
  signal RPIPE_input_done_pipe_347_inst_req_0 : boolean;
  signal RPIPE_input_done_pipe_347_inst_ack_0 : boolean;
  signal RPIPE_input_done_pipe_347_inst_req_1 : boolean;
  signal RPIPE_input_done_pipe_347_inst_ack_1 : boolean;
  signal do_while_stmt_350_branch_req_0 : boolean;
  signal phi_stmt_352_req_0 : boolean;
  signal phi_stmt_352_req_1 : boolean;
  signal phi_stmt_352_ack_0 : boolean;
  signal nmycount_374_354_buf_req_0 : boolean;
  signal nmycount_374_354_buf_ack_0 : boolean;
  signal nmycount_374_354_buf_req_1 : boolean;
  signal nmycount_374_354_buf_ack_1 : boolean;
  signal start_add_355_buf_req_0 : boolean;
  signal start_add_355_buf_ack_0 : boolean;
  signal start_add_355_buf_req_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "loadKernelChannel_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 128) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(63 downto 0) <= start_add;
  start_add_buffer <= in_buffer_data_out(63 downto 0);
  in_buffer_data_in(127 downto 64) <= end_add;
  end_add_buffer <= in_buffer_data_out(127 downto 64);
  in_buffer_data_in(tag_length + 127 downto 128) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 127 downto 128);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  loadKernelChannel_CP_676_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "loadKernelChannel_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= loadKernelChannel_CP_676_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= loadKernelChannel_CP_676_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= loadKernelChannel_CP_676_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  loadKernelChannel_CP_676: Block -- control-path 
    signal loadKernelChannel_CP_676_elements: BooleanArray(94 downto 0);
    -- 
  begin -- 
    loadKernelChannel_CP_676_elements(0) <= loadKernelChannel_CP_676_start;
    loadKernelChannel_CP_676_symbol <= loadKernelChannel_CP_676_elements(94);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	7 
    -- CP-element group 0: 	6 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (29) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/$entry
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/addr_of_334_update_start_
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_index_resized_1
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_index_scaled_1
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_index_computed_1
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_index_resize_1/$entry
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_index_resize_1/$exit
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_index_resize_1/index_resize_req
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_index_resize_1/index_resize_ack
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_index_scale_1/$entry
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_index_scale_1/$exit
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_index_scale_1/scale_rename_req
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_index_scale_1/scale_rename_ack
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_final_index_sum_regn_update_start
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_final_index_sum_regn_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_final_index_sum_regn_Sample/req
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_final_index_sum_regn_Update/$entry
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_final_index_sum_regn_Update/req
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/addr_of_334_complete/$entry
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/addr_of_334_complete/req
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_update_start_
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Update/$entry
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/RPIPE_input_done_pipe_347_sample_start_
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/RPIPE_input_done_pipe_347_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_328_to_assign_stmt_348/RPIPE_input_done_pipe_347_Sample/rr
      -- 
    req_726_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_726_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(0), ack => addr_of_334_final_reg_req_1); -- 
    req_706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(0), ack => array_obj_ref_333_index_offset_req_0); -- 
    req_711_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_711_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(0), ack => array_obj_ref_333_index_offset_req_1); -- 
    rr_785_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_785_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(0), ack => RPIPE_input_done_pipe_347_inst_req_0); -- 
    cr_771_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_771_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(0), ack => ptr_deref_338_load_0_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	9 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_final_index_sum_regn_sample_complete
      -- CP-element group 1: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_final_index_sum_regn_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_final_index_sum_regn_Sample/ack
      -- 
    ack_707_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_333_index_offset_ack_0, ack => loadKernelChannel_CP_676_elements(1)); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (11) 
      -- CP-element group 2: 	 assign_stmt_328_to_assign_stmt_348/addr_of_334_sample_start_
      -- CP-element group 2: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_root_address_calculated
      -- CP-element group 2: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_offset_calculated
      -- CP-element group 2: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_final_index_sum_regn_Update/$exit
      -- CP-element group 2: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_final_index_sum_regn_Update/ack
      -- CP-element group 2: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_base_plus_offset/$entry
      -- CP-element group 2: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_base_plus_offset/$exit
      -- CP-element group 2: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 assign_stmt_328_to_assign_stmt_348/array_obj_ref_333_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 assign_stmt_328_to_assign_stmt_348/addr_of_334_request/$entry
      -- CP-element group 2: 	 assign_stmt_328_to_assign_stmt_348/addr_of_334_request/req
      -- 
    ack_712_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_333_index_offset_ack_1, ack => loadKernelChannel_CP_676_elements(2)); -- 
    req_721_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_721_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(2), ack => addr_of_334_final_reg_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 assign_stmt_328_to_assign_stmt_348/addr_of_334_sample_completed_
      -- CP-element group 3: 	 assign_stmt_328_to_assign_stmt_348/addr_of_334_request/$exit
      -- CP-element group 3: 	 assign_stmt_328_to_assign_stmt_348/addr_of_334_request/ack
      -- 
    ack_722_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_334_final_reg_ack_0, ack => loadKernelChannel_CP_676_elements(3)); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (24) 
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/addr_of_334_update_completed_
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/addr_of_334_complete/$exit
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/addr_of_334_complete/ack
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_sample_start_
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_base_address_calculated
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_word_address_calculated
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_root_address_calculated
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_base_address_resized
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_base_addr_resize/$entry
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_base_addr_resize/$exit
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_base_addr_resize/base_resize_req
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_base_addr_resize/base_resize_ack
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_base_plus_offset/$entry
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_base_plus_offset/$exit
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_base_plus_offset/sum_rename_req
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_base_plus_offset/sum_rename_ack
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_word_addrgen/$entry
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_word_addrgen/$exit
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_word_addrgen/root_register_req
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_word_addrgen/root_register_ack
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Sample/$entry
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Sample/word_access_start/$entry
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Sample/word_access_start/word_0/$entry
      -- CP-element group 4: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Sample/word_access_start/word_0/rr
      -- 
    ack_727_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_334_final_reg_ack_1, ack => loadKernelChannel_CP_676_elements(4)); -- 
    rr_760_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_760_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(4), ack => ptr_deref_338_load_0_req_0); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (5) 
      -- CP-element group 5: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_sample_completed_
      -- CP-element group 5: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Sample/$exit
      -- CP-element group 5: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Sample/word_access_start/$exit
      -- CP-element group 5: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Sample/word_access_start/word_0/$exit
      -- CP-element group 5: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Sample/word_access_start/word_0/ra
      -- 
    ra_761_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_338_load_0_ack_0, ack => loadKernelChannel_CP_676_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	0 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	9 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_update_completed_
      -- CP-element group 6: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Update/$exit
      -- CP-element group 6: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Update/word_access_complete/$exit
      -- CP-element group 6: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Update/word_access_complete/word_0/$exit
      -- CP-element group 6: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Update/word_access_complete/word_0/ca
      -- CP-element group 6: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Update/ptr_deref_338_Merge/$entry
      -- CP-element group 6: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Update/ptr_deref_338_Merge/$exit
      -- CP-element group 6: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Update/ptr_deref_338_Merge/merge_req
      -- CP-element group 6: 	 assign_stmt_328_to_assign_stmt_348/ptr_deref_338_Update/ptr_deref_338_Merge/merge_ack
      -- 
    ca_772_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_338_load_0_ack_1, ack => loadKernelChannel_CP_676_elements(6)); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	0 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 assign_stmt_328_to_assign_stmt_348/RPIPE_input_done_pipe_347_sample_completed_
      -- CP-element group 7: 	 assign_stmt_328_to_assign_stmt_348/RPIPE_input_done_pipe_347_update_start_
      -- CP-element group 7: 	 assign_stmt_328_to_assign_stmt_348/RPIPE_input_done_pipe_347_Sample/$exit
      -- CP-element group 7: 	 assign_stmt_328_to_assign_stmt_348/RPIPE_input_done_pipe_347_Sample/ra
      -- CP-element group 7: 	 assign_stmt_328_to_assign_stmt_348/RPIPE_input_done_pipe_347_Update/$entry
      -- CP-element group 7: 	 assign_stmt_328_to_assign_stmt_348/RPIPE_input_done_pipe_347_Update/cr
      -- 
    ra_786_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_done_pipe_347_inst_ack_0, ack => loadKernelChannel_CP_676_elements(7)); -- 
    cr_790_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_790_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(7), ack => RPIPE_input_done_pipe_347_inst_req_1); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 assign_stmt_328_to_assign_stmt_348/RPIPE_input_done_pipe_347_update_completed_
      -- CP-element group 8: 	 assign_stmt_328_to_assign_stmt_348/RPIPE_input_done_pipe_347_Update/$exit
      -- CP-element group 8: 	 assign_stmt_328_to_assign_stmt_348/RPIPE_input_done_pipe_347_Update/ca
      -- 
    ca_791_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_done_pipe_347_inst_ack_1, ack => loadKernelChannel_CP_676_elements(8)); -- 
    -- CP-element group 9:  join  transition  place  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	1 
    -- CP-element group 9: 	8 
    -- CP-element group 9: 	6 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9:  members (4) 
      -- CP-element group 9: 	 assign_stmt_328_to_assign_stmt_348/$exit
      -- CP-element group 9: 	 branch_block_stmt_349/$entry
      -- CP-element group 9: 	 branch_block_stmt_349/branch_block_stmt_349__entry__
      -- CP-element group 9: 	 branch_block_stmt_349/do_while_stmt_350__entry__
      -- 
    loadKernelChannel_cp_element_group_9: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 36) := "loadKernelChannel_cp_element_group_9"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(1) & loadKernelChannel_CP_676_elements(8) & loadKernelChannel_CP_676_elements(6);
      gj_loadKernelChannel_cp_element_group_9 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(9), clk => clk, reset => reset); --
    end block;
    -- CP-element group 10:  fork  transition  place  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	90 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	92 
    -- CP-element group 10: 	91 
    -- CP-element group 10:  members (10) 
      -- CP-element group 10: 	 assign_stmt_433/$entry
      -- CP-element group 10: 	 assign_stmt_433/type_cast_432_sample_start_
      -- CP-element group 10: 	 assign_stmt_433/type_cast_432_update_start_
      -- CP-element group 10: 	 assign_stmt_433/type_cast_432_Sample/rr
      -- CP-element group 10: 	 assign_stmt_433/type_cast_432_Update/cr
      -- CP-element group 10: 	 assign_stmt_433/type_cast_432_Sample/$entry
      -- CP-element group 10: 	 assign_stmt_433/type_cast_432_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_349/$exit
      -- CP-element group 10: 	 branch_block_stmt_349/branch_block_stmt_349__exit__
      -- CP-element group 10: 	 branch_block_stmt_349/do_while_stmt_350__exit__
      -- 
    rr_1099_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1099_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(10), ack => type_cast_432_inst_req_0); -- 
    cr_1104_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1104_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(10), ack => type_cast_432_inst_req_1); -- 
    loadKernelChannel_CP_676_elements(10) <= loadKernelChannel_CP_676_elements(90);
    -- CP-element group 11:  transition  place  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	17 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_349/do_while_stmt_350/$entry
      -- CP-element group 11: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350__entry__
      -- 
    loadKernelChannel_CP_676_elements(11) <= loadKernelChannel_CP_676_elements(9);
    -- CP-element group 12:  merge  place  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	90 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350__exit__
      -- 
    -- Element group loadKernelChannel_CP_676_elements(12) is bound as output of CP function.
    -- CP-element group 13:  merge  place  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	16 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 branch_block_stmt_349/do_while_stmt_350/loop_back
      -- 
    -- Element group loadKernelChannel_CP_676_elements(13) is bound as output of CP function.
    -- CP-element group 14:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	19 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	88 
    -- CP-element group 14: 	89 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_349/do_while_stmt_350/loop_taken/$entry
      -- CP-element group 14: 	 branch_block_stmt_349/do_while_stmt_350/loop_exit/$entry
      -- CP-element group 14: 	 branch_block_stmt_349/do_while_stmt_350/condition_done
      -- 
    loadKernelChannel_CP_676_elements(14) <= loadKernelChannel_CP_676_elements(19);
    -- CP-element group 15:  branch  place  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	87 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_349/do_while_stmt_350/loop_body_done
      -- 
    loadKernelChannel_CP_676_elements(15) <= loadKernelChannel_CP_676_elements(87);
    -- CP-element group 16:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	13 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	47 
    -- CP-element group 16: 	30 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/back_edge_to_loop_body
      -- 
    loadKernelChannel_CP_676_elements(16) <= loadKernelChannel_CP_676_elements(13);
    -- CP-element group 17:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	11 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	32 
    -- CP-element group 17: 	49 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/first_time_through_loop_body
      -- 
    loadKernelChannel_CP_676_elements(17) <= loadKernelChannel_CP_676_elements(11);
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	43 
    -- CP-element group 18: 	44 
    -- CP-element group 18: 	86 
    -- CP-element group 18: 	64 
    -- CP-element group 18: 	65 
    -- CP-element group 18: 	24 
    -- CP-element group 18: 	25 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/$entry
      -- CP-element group 18: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/loop_body_start
      -- 
    -- Element group loadKernelChannel_CP_676_elements(18) is bound as output of CP function.
    -- CP-element group 19:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	86 
    -- CP-element group 19: 	29 
    -- CP-element group 19: 	23 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	14 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/condition_evaluated
      -- 
    condition_evaluated_813_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_813_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(19), ack => do_while_stmt_350_branch_req_0); -- 
    loadKernelChannel_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(86) & loadKernelChannel_CP_676_elements(29) & loadKernelChannel_CP_676_elements(23);
      gj_loadKernelChannel_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	43 
    -- CP-element group 20: 	24 
    -- CP-element group 20: marked-predecessors 
    -- CP-element group 20: 	23 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	26 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_356_sample_start__ps
      -- CP-element group 20: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/aggregated_phi_sample_req
      -- 
    loadKernelChannel_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(43) & loadKernelChannel_CP_676_elements(24) & loadKernelChannel_CP_676_elements(23);
      gj_loadKernelChannel_cp_element_group_20 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	45 
    -- CP-element group 21: 	27 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	83 
    -- CP-element group 21: 	79 
    -- CP-element group 21: 	75 
    -- CP-element group 21: 	87 
    -- CP-element group 21: marked-successors 
    -- CP-element group 21: 	43 
    -- CP-element group 21: 	24 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_356_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/aggregated_phi_sample_ack
      -- CP-element group 21: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_352_sample_completed_
      -- 
    loadKernelChannel_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(45) & loadKernelChannel_CP_676_elements(27);
      gj_loadKernelChannel_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	44 
    -- CP-element group 22: 	25 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	28 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_356_update_start__ps
      -- CP-element group 22: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/aggregated_phi_update_req
      -- 
    loadKernelChannel_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(44) & loadKernelChannel_CP_676_elements(25);
      gj_loadKernelChannel_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	46 
    -- CP-element group 23: 	29 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	19 
    -- CP-element group 23: marked-successors 
    -- CP-element group 23: 	20 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/aggregated_phi_update_ack
      -- 
    loadKernelChannel_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(46) & loadKernelChannel_CP_676_elements(29);
      gj_loadKernelChannel_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  join  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	18 
    -- CP-element group 24: marked-predecessors 
    -- CP-element group 24: 	21 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	20 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_352_sample_start_
      -- 
    loadKernelChannel_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(18) & loadKernelChannel_CP_676_elements(21);
      gj_loadKernelChannel_cp_element_group_24 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(24), clk => clk, reset => reset); --
    end block;
    -- CP-element group 25:  join  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	18 
    -- CP-element group 25: marked-predecessors 
    -- CP-element group 25: 	61 
    -- CP-element group 25: 	80 
    -- CP-element group 25: 	29 
    -- CP-element group 25: 	72 
    -- CP-element group 25: 	66 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	22 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_352_update_start_
      -- 
    loadKernelChannel_cp_element_group_25: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_25"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(18) & loadKernelChannel_CP_676_elements(61) & loadKernelChannel_CP_676_elements(80) & loadKernelChannel_CP_676_elements(29) & loadKernelChannel_CP_676_elements(72) & loadKernelChannel_CP_676_elements(66);
      gj_loadKernelChannel_cp_element_group_25 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(25), clk => clk, reset => reset); --
    end block;
    -- CP-element group 26:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	20 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_352_sample_start__ps
      -- 
    loadKernelChannel_CP_676_elements(26) <= loadKernelChannel_CP_676_elements(20);
    -- CP-element group 27:  join  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	21 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_352_sample_completed__ps
      -- 
    -- Element group loadKernelChannel_CP_676_elements(27) is bound as output of CP function.
    -- CP-element group 28:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	22 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_352_update_start__ps
      -- 
    loadKernelChannel_CP_676_elements(28) <= loadKernelChannel_CP_676_elements(22);
    -- CP-element group 29:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	60 
    -- CP-element group 29: 	78 
    -- CP-element group 29: 	70 
    -- CP-element group 29: 	66 
    -- CP-element group 29: 	19 
    -- CP-element group 29: 	23 
    -- CP-element group 29: marked-successors 
    -- CP-element group 29: 	25 
    -- CP-element group 29:  members (15) 
      -- CP-element group 29: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_index_resize_1/index_resize_req
      -- CP-element group 29: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_index_scale_1/scale_rename_ack
      -- CP-element group 29: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_index_scale_1/$exit
      -- CP-element group 29: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_index_resize_1/index_resize_ack
      -- CP-element group 29: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_final_index_sum_regn_Sample/req
      -- CP-element group 29: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_index_scale_1/scale_rename_req
      -- CP-element group 29: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_index_scale_1/$entry
      -- CP-element group 29: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_final_index_sum_regn_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_index_resize_1/$exit
      -- CP-element group 29: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_index_resize_1/$entry
      -- CP-element group 29: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_index_computed_1
      -- CP-element group 29: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_index_scaled_1
      -- CP-element group 29: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_index_resized_1
      -- CP-element group 29: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_352_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_352_update_completed__ps
      -- 
    req_965_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_965_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(29), ack => array_obj_ref_397_index_offset_req_0); -- 
    -- Element group loadKernelChannel_CP_676_elements(29) is bound as output of CP function.
    -- CP-element group 30:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	16 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_352_loopback_trigger
      -- 
    loadKernelChannel_CP_676_elements(30) <= loadKernelChannel_CP_676_elements(16);
    -- CP-element group 31:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (2) 
      -- CP-element group 31: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_352_loopback_sample_req
      -- CP-element group 31: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_352_loopback_sample_req_ps
      -- 
    phi_stmt_352_loopback_sample_req_828_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_352_loopback_sample_req_828_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(31), ack => phi_stmt_352_req_0); -- 
    -- Element group loadKernelChannel_CP_676_elements(31) is bound as output of CP function.
    -- CP-element group 32:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	17 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_352_entry_trigger
      -- 
    loadKernelChannel_CP_676_elements(32) <= loadKernelChannel_CP_676_elements(17);
    -- CP-element group 33:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (2) 
      -- CP-element group 33: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_352_entry_sample_req
      -- CP-element group 33: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_352_entry_sample_req_ps
      -- 
    phi_stmt_352_entry_sample_req_831_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_352_entry_sample_req_831_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(33), ack => phi_stmt_352_req_1); -- 
    -- Element group loadKernelChannel_CP_676_elements(33) is bound as output of CP function.
    -- CP-element group 34:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (2) 
      -- CP-element group 34: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_352_phi_mux_ack
      -- CP-element group 34: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_352_phi_mux_ack_ps
      -- 
    phi_stmt_352_phi_mux_ack_834_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_352_ack_0, ack => loadKernelChannel_CP_676_elements(34)); -- 
    -- CP-element group 35:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	37 
    -- CP-element group 35:  members (4) 
      -- CP-element group 35: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nmycount_354_sample_start__ps
      -- CP-element group 35: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nmycount_354_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nmycount_354_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nmycount_354_Sample/req
      -- 
    req_847_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_847_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(35), ack => nmycount_374_354_buf_req_0); -- 
    -- Element group loadKernelChannel_CP_676_elements(35) is bound as output of CP function.
    -- CP-element group 36:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	38 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nmycount_354_update_start__ps
      -- CP-element group 36: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nmycount_354_update_start_
      -- CP-element group 36: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nmycount_354_Update/$entry
      -- CP-element group 36: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nmycount_354_Update/req
      -- 
    req_852_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_852_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(36), ack => nmycount_374_354_buf_req_1); -- 
    -- Element group loadKernelChannel_CP_676_elements(36) is bound as output of CP function.
    -- CP-element group 37:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	35 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (4) 
      -- CP-element group 37: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nmycount_354_sample_completed__ps
      -- CP-element group 37: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nmycount_354_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nmycount_354_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nmycount_354_Sample/ack
      -- 
    ack_848_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmycount_374_354_buf_ack_0, ack => loadKernelChannel_CP_676_elements(37)); -- 
    -- CP-element group 38:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	36 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (4) 
      -- CP-element group 38: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nmycount_354_update_completed__ps
      -- CP-element group 38: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nmycount_354_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nmycount_354_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nmycount_354_Update/ack
      -- 
    ack_853_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmycount_374_354_buf_ack_1, ack => loadKernelChannel_CP_676_elements(38)); -- 
    -- CP-element group 39:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	41 
    -- CP-element group 39:  members (4) 
      -- CP-element group 39: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_start_add_355_sample_start__ps
      -- CP-element group 39: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_start_add_355_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_start_add_355_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_start_add_355_Sample/req
      -- 
    req_865_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_865_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(39), ack => start_add_355_buf_req_0); -- 
    -- Element group loadKernelChannel_CP_676_elements(39) is bound as output of CP function.
    -- CP-element group 40:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	42 
    -- CP-element group 40:  members (4) 
      -- CP-element group 40: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_start_add_355_update_start__ps
      -- CP-element group 40: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_start_add_355_update_start_
      -- CP-element group 40: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_start_add_355_Update/$entry
      -- CP-element group 40: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_start_add_355_Update/req
      -- 
    req_870_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_870_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(40), ack => start_add_355_buf_req_1); -- 
    -- Element group loadKernelChannel_CP_676_elements(40) is bound as output of CP function.
    -- CP-element group 41:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	39 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (4) 
      -- CP-element group 41: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_start_add_355_sample_completed__ps
      -- CP-element group 41: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_start_add_355_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_start_add_355_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_start_add_355_Sample/ack
      -- 
    ack_866_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => start_add_355_buf_ack_0, ack => loadKernelChannel_CP_676_elements(41)); -- 
    -- CP-element group 42:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	40 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (4) 
      -- CP-element group 42: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_start_add_355_Update/ack
      -- CP-element group 42: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_start_add_355_update_completed__ps
      -- CP-element group 42: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_start_add_355_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_start_add_355_Update/$exit
      -- 
    ack_871_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => start_add_355_buf_ack_1, ack => loadKernelChannel_CP_676_elements(42)); -- 
    -- CP-element group 43:  join  transition  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	18 
    -- CP-element group 43: marked-predecessors 
    -- CP-element group 43: 	81 
    -- CP-element group 43: 	85 
    -- CP-element group 43: 	77 
    -- CP-element group 43: 	21 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	20 
    -- CP-element group 43:  members (1) 
      -- CP-element group 43: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_356_sample_start_
      -- 
    loadKernelChannel_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(18) & loadKernelChannel_CP_676_elements(81) & loadKernelChannel_CP_676_elements(85) & loadKernelChannel_CP_676_elements(77) & loadKernelChannel_CP_676_elements(21);
      gj_loadKernelChannel_cp_element_group_43 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  join  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	18 
    -- CP-element group 44: marked-predecessors 
    -- CP-element group 44: 	61 
    -- CP-element group 44: 	46 
    -- CP-element group 44: 	84 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	22 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_356_update_start_
      -- 
    loadKernelChannel_cp_element_group_44: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_44"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(18) & loadKernelChannel_CP_676_elements(61) & loadKernelChannel_CP_676_elements(46) & loadKernelChannel_CP_676_elements(84);
      gj_loadKernelChannel_cp_element_group_44 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(44), clk => clk, reset => reset); --
    end block;
    -- CP-element group 45:  join  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	21 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_356_sample_completed__ps
      -- 
    -- Element group loadKernelChannel_CP_676_elements(45) is bound as output of CP function.
    -- CP-element group 46:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	60 
    -- CP-element group 46: 	82 
    -- CP-element group 46: 	23 
    -- CP-element group 46: marked-successors 
    -- CP-element group 46: 	44 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_356_update_completed__ps
      -- CP-element group 46: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_356_update_completed_
      -- 
    -- Element group loadKernelChannel_CP_676_elements(46) is bound as output of CP function.
    -- CP-element group 47:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	16 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_356_loopback_trigger
      -- 
    loadKernelChannel_CP_676_elements(47) <= loadKernelChannel_CP_676_elements(16);
    -- CP-element group 48:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (2) 
      -- CP-element group 48: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_356_loopback_sample_req_ps
      -- CP-element group 48: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_356_loopback_sample_req
      -- 
    phi_stmt_356_loopback_sample_req_882_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_356_loopback_sample_req_882_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(48), ack => phi_stmt_356_req_0); -- 
    -- Element group loadKernelChannel_CP_676_elements(48) is bound as output of CP function.
    -- CP-element group 49:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	17 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_356_entry_trigger
      -- 
    loadKernelChannel_CP_676_elements(49) <= loadKernelChannel_CP_676_elements(17);
    -- CP-element group 50:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (2) 
      -- CP-element group 50: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_356_entry_sample_req
      -- CP-element group 50: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_356_entry_sample_req_ps
      -- 
    phi_stmt_356_entry_sample_req_885_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_356_entry_sample_req_885_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(50), ack => phi_stmt_356_req_1); -- 
    -- Element group loadKernelChannel_CP_676_elements(50) is bound as output of CP function.
    -- CP-element group 51:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (2) 
      -- CP-element group 51: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_356_phi_mux_ack
      -- CP-element group 51: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/phi_stmt_356_phi_mux_ack_ps
      -- 
    phi_stmt_356_phi_mux_ack_888_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_356_ack_0, ack => loadKernelChannel_CP_676_elements(51)); -- 
    -- CP-element group 52:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (4) 
      -- CP-element group 52: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nfetch_val_358_sample_start__ps
      -- CP-element group 52: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nfetch_val_358_sample_start_
      -- CP-element group 52: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nfetch_val_358_Sample/$entry
      -- CP-element group 52: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nfetch_val_358_Sample/req
      -- 
    req_901_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_901_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(52), ack => nfetch_val_419_358_buf_req_0); -- 
    -- Element group loadKernelChannel_CP_676_elements(52) is bound as output of CP function.
    -- CP-element group 53:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (4) 
      -- CP-element group 53: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nfetch_val_358_Update/req
      -- CP-element group 53: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nfetch_val_358_update_start__ps
      -- CP-element group 53: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nfetch_val_358_update_start_
      -- CP-element group 53: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nfetch_val_358_Update/$entry
      -- 
    req_906_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_906_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(53), ack => nfetch_val_419_358_buf_req_1); -- 
    -- Element group loadKernelChannel_CP_676_elements(53) is bound as output of CP function.
    -- CP-element group 54:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (4) 
      -- CP-element group 54: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nfetch_val_358_sample_completed__ps
      -- CP-element group 54: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nfetch_val_358_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nfetch_val_358_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nfetch_val_358_Sample/ack
      -- 
    ack_902_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nfetch_val_419_358_buf_ack_0, ack => loadKernelChannel_CP_676_elements(54)); -- 
    -- CP-element group 55:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (4) 
      -- CP-element group 55: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nfetch_val_358_Update/ack
      -- CP-element group 55: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nfetch_val_358_update_completed__ps
      -- CP-element group 55: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nfetch_val_358_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_nfetch_val_358_Update/$exit
      -- 
    ack_907_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nfetch_val_419_358_buf_ack_1, ack => loadKernelChannel_CP_676_elements(55)); -- 
    -- CP-element group 56:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	58 
    -- CP-element group 56:  members (4) 
      -- CP-element group 56: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_my_fetch_359_sample_start__ps
      -- CP-element group 56: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_my_fetch_359_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_my_fetch_359_Sample/req
      -- CP-element group 56: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_my_fetch_359_sample_start_
      -- 
    req_919_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_919_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(56), ack => my_fetch_339_359_buf_req_0); -- 
    -- Element group loadKernelChannel_CP_676_elements(56) is bound as output of CP function.
    -- CP-element group 57:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	59 
    -- CP-element group 57:  members (4) 
      -- CP-element group 57: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_my_fetch_359_update_start_
      -- CP-element group 57: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_my_fetch_359_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_my_fetch_359_Update/req
      -- CP-element group 57: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_my_fetch_359_update_start__ps
      -- 
    req_924_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_924_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(57), ack => my_fetch_339_359_buf_req_1); -- 
    -- Element group loadKernelChannel_CP_676_elements(57) is bound as output of CP function.
    -- CP-element group 58:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	56 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (4) 
      -- CP-element group 58: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_my_fetch_359_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_my_fetch_359_Sample/ack
      -- CP-element group 58: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_my_fetch_359_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_my_fetch_359_sample_completed__ps
      -- 
    ack_920_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_fetch_339_359_buf_ack_0, ack => loadKernelChannel_CP_676_elements(58)); -- 
    -- CP-element group 59:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	57 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (4) 
      -- CP-element group 59: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_my_fetch_359_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_my_fetch_359_update_completed__ps
      -- CP-element group 59: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_my_fetch_359_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/R_my_fetch_359_Update/ack
      -- 
    ack_925_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_fetch_339_359_buf_ack_1, ack => loadKernelChannel_CP_676_elements(59)); -- 
    -- CP-element group 60:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	46 
    -- CP-element group 60: 	29 
    -- CP-element group 60: marked-predecessors 
    -- CP-element group 60: 	62 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/WPIPE_kernel_pipe1_381_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/WPIPE_kernel_pipe1_381_Sample/req
      -- CP-element group 60: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/WPIPE_kernel_pipe1_381_sample_start_
      -- 
    req_934_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_934_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(60), ack => WPIPE_kernel_pipe1_381_inst_req_0); -- 
    loadKernelChannel_cp_element_group_60: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_60"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(46) & loadKernelChannel_CP_676_elements(29) & loadKernelChannel_CP_676_elements(62);
      gj_loadKernelChannel_cp_element_group_60 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(60), clk => clk, reset => reset); --
    end block;
    -- CP-element group 61:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61: marked-successors 
    -- CP-element group 61: 	44 
    -- CP-element group 61: 	25 
    -- CP-element group 61:  members (6) 
      -- CP-element group 61: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/WPIPE_kernel_pipe1_381_Update/$entry
      -- CP-element group 61: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/WPIPE_kernel_pipe1_381_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/WPIPE_kernel_pipe1_381_update_start_
      -- CP-element group 61: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/WPIPE_kernel_pipe1_381_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/WPIPE_kernel_pipe1_381_Sample/ack
      -- CP-element group 61: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/WPIPE_kernel_pipe1_381_Update/req
      -- 
    ack_935_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe1_381_inst_ack_0, ack => loadKernelChannel_CP_676_elements(61)); -- 
    req_939_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_939_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(61), ack => WPIPE_kernel_pipe1_381_inst_req_1); -- 
    -- CP-element group 62:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	87 
    -- CP-element group 62: marked-successors 
    -- CP-element group 62: 	60 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/WPIPE_kernel_pipe1_381_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/WPIPE_kernel_pipe1_381_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/WPIPE_kernel_pipe1_381_Update/ack
      -- 
    ack_940_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe1_381_inst_ack_1, ack => loadKernelChannel_CP_676_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	67 
    -- CP-element group 63: marked-predecessors 
    -- CP-element group 63: 	68 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	68 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/addr_of_398_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/addr_of_398_request/req
      -- CP-element group 63: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/addr_of_398_request/$entry
      -- 
    req_980_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_980_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(63), ack => addr_of_398_final_reg_req_0); -- 
    loadKernelChannel_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(67) & loadKernelChannel_CP_676_elements(68);
      gj_loadKernelChannel_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	18 
    -- CP-element group 64: marked-predecessors 
    -- CP-element group 64: 	76 
    -- CP-element group 64: 	69 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	69 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/addr_of_398_complete/$entry
      -- CP-element group 64: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/addr_of_398_complete/req
      -- CP-element group 64: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/addr_of_398_update_start_
      -- 
    req_985_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_985_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(64), ack => addr_of_398_final_reg_req_1); -- 
    loadKernelChannel_cp_element_group_64: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_64"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(18) & loadKernelChannel_CP_676_elements(76) & loadKernelChannel_CP_676_elements(69);
      gj_loadKernelChannel_cp_element_group_64 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(64), clk => clk, reset => reset); --
    end block;
    -- CP-element group 65:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	18 
    -- CP-element group 65: marked-predecessors 
    -- CP-element group 65: 	67 
    -- CP-element group 65: 	68 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	67 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_final_index_sum_regn_Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_final_index_sum_regn_Update/req
      -- CP-element group 65: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_final_index_sum_regn_update_start
      -- 
    req_970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(65), ack => array_obj_ref_397_index_offset_req_1); -- 
    loadKernelChannel_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(18) & loadKernelChannel_CP_676_elements(67) & loadKernelChannel_CP_676_elements(68);
      gj_loadKernelChannel_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	29 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	87 
    -- CP-element group 66: marked-successors 
    -- CP-element group 66: 	25 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_final_index_sum_regn_Sample/ack
      -- CP-element group 66: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_final_index_sum_regn_sample_complete
      -- CP-element group 66: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_final_index_sum_regn_Sample/$exit
      -- 
    ack_966_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_397_index_offset_ack_0, ack => loadKernelChannel_CP_676_elements(66)); -- 
    -- CP-element group 67:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	65 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	63 
    -- CP-element group 67: marked-successors 
    -- CP-element group 67: 	65 
    -- CP-element group 67:  members (8) 
      -- CP-element group 67: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_final_index_sum_regn_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_base_plus_offset/sum_rename_ack
      -- CP-element group 67: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_final_index_sum_regn_Update/ack
      -- CP-element group 67: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_base_plus_offset/$entry
      -- CP-element group 67: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_base_plus_offset/$exit
      -- CP-element group 67: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_base_plus_offset/sum_rename_req
      -- CP-element group 67: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_offset_calculated
      -- CP-element group 67: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/array_obj_ref_397_root_address_calculated
      -- 
    ack_971_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_397_index_offset_ack_1, ack => loadKernelChannel_CP_676_elements(67)); -- 
    -- CP-element group 68:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	63 
    -- CP-element group 68: successors 
    -- CP-element group 68: marked-successors 
    -- CP-element group 68: 	63 
    -- CP-element group 68: 	65 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/addr_of_398_request/ack
      -- CP-element group 68: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/addr_of_398_request/$exit
      -- CP-element group 68: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/addr_of_398_sample_completed_
      -- 
    ack_981_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_398_final_reg_ack_0, ack => loadKernelChannel_CP_676_elements(68)); -- 
    -- CP-element group 69:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	64 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	74 
    -- CP-element group 69: marked-successors 
    -- CP-element group 69: 	64 
    -- CP-element group 69:  members (19) 
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_base_plus_offset/$entry
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/addr_of_398_complete/$exit
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_word_addrgen/$exit
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/addr_of_398_complete/ack
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_base_plus_offset/$exit
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_word_addrgen/root_register_req
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_word_addrgen/$entry
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_base_plus_offset/sum_rename_req
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_base_addr_resize/$exit
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_base_address_calculated
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_base_plus_offset/sum_rename_ack
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_word_addrgen/root_register_ack
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_base_addr_resize/base_resize_req
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_base_addr_resize/base_resize_ack
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_base_addr_resize/$entry
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_base_address_resized
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/addr_of_398_update_completed_
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_root_address_calculated
      -- CP-element group 69: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_word_address_calculated
      -- 
    ack_986_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_398_final_reg_ack_1, ack => loadKernelChannel_CP_676_elements(69)); -- 
    -- CP-element group 70:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	29 
    -- CP-element group 70: marked-predecessors 
    -- CP-element group 70: 	72 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_402_Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_402_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_402_Sample/req
      -- 
    req_994_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_994_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(70), ack => W_fn_388_delayed_7_0_400_inst_req_0); -- 
    loadKernelChannel_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(29) & loadKernelChannel_CP_676_elements(72);
      gj_loadKernelChannel_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: marked-predecessors 
    -- CP-element group 71: 	76 
    -- CP-element group 71: 	73 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_402_update_start_
      -- CP-element group 71: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_402_Update/$entry
      -- CP-element group 71: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_402_Update/req
      -- 
    req_999_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_999_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(71), ack => W_fn_388_delayed_7_0_400_inst_req_1); -- 
    loadKernelChannel_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(76) & loadKernelChannel_CP_676_elements(73);
      gj_loadKernelChannel_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: marked-successors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: 	25 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_402_sample_completed_
      -- CP-element group 72: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_402_Sample/$exit
      -- CP-element group 72: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_402_Sample/ack
      -- 
    ack_995_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn_388_delayed_7_0_400_inst_ack_0, ack => loadKernelChannel_CP_676_elements(72)); -- 
    -- CP-element group 73:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73: marked-successors 
    -- CP-element group 73: 	71 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_402_update_completed_
      -- CP-element group 73: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_402_Update/$exit
      -- CP-element group 73: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_402_Update/ack
      -- 
    ack_1000_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn_388_delayed_7_0_400_inst_ack_1, ack => loadKernelChannel_CP_676_elements(73)); -- 
    -- CP-element group 74:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	69 
    -- CP-element group 74: 	73 
    -- CP-element group 74: marked-predecessors 
    -- CP-element group 74: 	76 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (5) 
      -- CP-element group 74: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Sample/$entry
      -- CP-element group 74: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Sample/word_access_start/word_0/$entry
      -- CP-element group 74: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Sample/word_access_start/$entry
      -- CP-element group 74: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Sample/word_access_start/word_0/rr
      -- CP-element group 74: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_sample_start_
      -- 
    rr_1033_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1033_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(74), ack => ptr_deref_406_load_0_req_0); -- 
    loadKernelChannel_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(69) & loadKernelChannel_CP_676_elements(73) & loadKernelChannel_CP_676_elements(76);
      gj_loadKernelChannel_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	21 
    -- CP-element group 75: marked-predecessors 
    -- CP-element group 75: 	77 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (5) 
      -- CP-element group 75: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Update/word_access_complete/word_0/cr
      -- CP-element group 75: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Update/word_access_complete/$entry
      -- CP-element group 75: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_update_start_
      -- CP-element group 75: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Update/word_access_complete/word_0/$entry
      -- 
    cr_1044_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1044_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(75), ack => ptr_deref_406_load_0_req_1); -- 
    loadKernelChannel_cp_element_group_75: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_75"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(21) & loadKernelChannel_CP_676_elements(77);
      gj_loadKernelChannel_cp_element_group_75 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(75), clk => clk, reset => reset); --
    end block;
    -- CP-element group 76:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: marked-successors 
    -- CP-element group 76: 	64 
    -- CP-element group 76: 	71 
    -- CP-element group 76: 	74 
    -- CP-element group 76:  members (5) 
      -- CP-element group 76: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Sample/$exit
      -- CP-element group 76: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Sample/word_access_start/word_0/$exit
      -- CP-element group 76: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Sample/word_access_start/word_0/ra
      -- CP-element group 76: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_sample_completed_
      -- CP-element group 76: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Sample/word_access_start/$exit
      -- 
    ra_1034_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_406_load_0_ack_0, ack => loadKernelChannel_CP_676_elements(76)); -- 
    -- CP-element group 77:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	87 
    -- CP-element group 77: marked-successors 
    -- CP-element group 77: 	43 
    -- CP-element group 77: 	75 
    -- CP-element group 77:  members (9) 
      -- CP-element group 77: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Update/$exit
      -- CP-element group 77: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Update/word_access_complete/$exit
      -- CP-element group 77: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Update/word_access_complete/word_0/ca
      -- CP-element group 77: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_update_completed_
      -- CP-element group 77: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Update/word_access_complete/word_0/$exit
      -- CP-element group 77: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Update/ptr_deref_406_Merge/merge_ack
      -- CP-element group 77: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Update/ptr_deref_406_Merge/merge_req
      -- CP-element group 77: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Update/ptr_deref_406_Merge/$exit
      -- CP-element group 77: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/ptr_deref_406_Update/ptr_deref_406_Merge/$entry
      -- 
    ca_1045_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_406_load_0_ack_1, ack => loadKernelChannel_CP_676_elements(77)); -- 
    -- CP-element group 78:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	29 
    -- CP-element group 78: marked-predecessors 
    -- CP-element group 78: 	80 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	80 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_410_Sample/$entry
      -- CP-element group 78: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_410_Sample/req
      -- CP-element group 78: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_410_sample_start_
      -- 
    req_1058_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1058_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(78), ack => W_fn_394_delayed_13_0_408_inst_req_0); -- 
    loadKernelChannel_cp_element_group_78: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_78"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(29) & loadKernelChannel_CP_676_elements(80);
      gj_loadKernelChannel_cp_element_group_78 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(78), clk => clk, reset => reset); --
    end block;
    -- CP-element group 79:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	21 
    -- CP-element group 79: marked-predecessors 
    -- CP-element group 79: 	81 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	81 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_410_update_start_
      -- CP-element group 79: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_410_Update/$entry
      -- CP-element group 79: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_410_Update/req
      -- 
    req_1063_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1063_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(79), ack => W_fn_394_delayed_13_0_408_inst_req_1); -- 
    loadKernelChannel_cp_element_group_79: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_79"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(21) & loadKernelChannel_CP_676_elements(81);
      gj_loadKernelChannel_cp_element_group_79 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(79), clk => clk, reset => reset); --
    end block;
    -- CP-element group 80:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: successors 
    -- CP-element group 80: marked-successors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: 	25 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_410_Sample/$exit
      -- CP-element group 80: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_410_Sample/ack
      -- CP-element group 80: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_410_sample_completed_
      -- 
    ack_1059_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn_394_delayed_13_0_408_inst_ack_0, ack => loadKernelChannel_CP_676_elements(80)); -- 
    -- CP-element group 81:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	79 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	87 
    -- CP-element group 81: marked-successors 
    -- CP-element group 81: 	43 
    -- CP-element group 81: 	79 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_410_update_completed_
      -- CP-element group 81: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_410_Update/$exit
      -- CP-element group 81: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_410_Update/ack
      -- 
    ack_1064_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn_394_delayed_13_0_408_inst_ack_1, ack => loadKernelChannel_CP_676_elements(81)); -- 
    -- CP-element group 82:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	46 
    -- CP-element group 82: marked-predecessors 
    -- CP-element group 82: 	84 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	84 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_413_Sample/$entry
      -- CP-element group 82: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_413_sample_start_
      -- CP-element group 82: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_413_Sample/req
      -- 
    req_1072_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1072_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(82), ack => W_fetch_val_396_delayed_13_0_411_inst_req_0); -- 
    loadKernelChannel_cp_element_group_82: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_82"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(46) & loadKernelChannel_CP_676_elements(84);
      gj_loadKernelChannel_cp_element_group_82 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(82), clk => clk, reset => reset); --
    end block;
    -- CP-element group 83:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	21 
    -- CP-element group 83: marked-predecessors 
    -- CP-element group 83: 	85 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	85 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_413_update_start_
      -- CP-element group 83: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_413_Update/req
      -- CP-element group 83: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_413_Update/$entry
      -- 
    req_1077_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1077_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(83), ack => W_fetch_val_396_delayed_13_0_411_inst_req_1); -- 
    loadKernelChannel_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(21) & loadKernelChannel_CP_676_elements(85);
      gj_loadKernelChannel_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: successors 
    -- CP-element group 84: marked-successors 
    -- CP-element group 84: 	44 
    -- CP-element group 84: 	82 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_413_sample_completed_
      -- CP-element group 84: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_413_Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_413_Sample/ack
      -- 
    ack_1073_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_val_396_delayed_13_0_411_inst_ack_0, ack => loadKernelChannel_CP_676_elements(84)); -- 
    -- CP-element group 85:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	83 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85: marked-successors 
    -- CP-element group 85: 	43 
    -- CP-element group 85: 	83 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_413_update_completed_
      -- CP-element group 85: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_413_Update/ack
      -- CP-element group 85: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/assign_stmt_413_Update/$exit
      -- 
    ack_1078_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_val_396_delayed_13_0_411_inst_ack_1, ack => loadKernelChannel_CP_676_elements(85)); -- 
    -- CP-element group 86:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	18 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	19 
    -- CP-element group 86:  members (1) 
      -- CP-element group 86: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group loadKernelChannel_CP_676_elements(86) is a control-delay.
    cp_element_86_delay: control_delay_element  generic map(name => " 86_delay", delay_value => 1)  port map(req => loadKernelChannel_CP_676_elements(18), ack => loadKernelChannel_CP_676_elements(86), clk => clk, reset =>reset);
    -- CP-element group 87:  join  transition  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	81 
    -- CP-element group 87: 	85 
    -- CP-element group 87: 	77 
    -- CP-element group 87: 	62 
    -- CP-element group 87: 	66 
    -- CP-element group 87: 	21 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	15 
    -- CP-element group 87:  members (1) 
      -- CP-element group 87: 	 branch_block_stmt_349/do_while_stmt_350/do_while_stmt_350_loop_body/$exit
      -- 
    loadKernelChannel_cp_element_group_87: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_87"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= loadKernelChannel_CP_676_elements(81) & loadKernelChannel_CP_676_elements(85) & loadKernelChannel_CP_676_elements(77) & loadKernelChannel_CP_676_elements(62) & loadKernelChannel_CP_676_elements(66) & loadKernelChannel_CP_676_elements(21);
      gj_loadKernelChannel_cp_element_group_87 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_676_elements(87), clk => clk, reset => reset); --
    end block;
    -- CP-element group 88:  transition  input  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	14 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (2) 
      -- CP-element group 88: 	 branch_block_stmt_349/do_while_stmt_350/loop_exit/ack
      -- CP-element group 88: 	 branch_block_stmt_349/do_while_stmt_350/loop_exit/$exit
      -- 
    ack_1083_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_350_branch_ack_0, ack => loadKernelChannel_CP_676_elements(88)); -- 
    -- CP-element group 89:  transition  input  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	14 
    -- CP-element group 89: successors 
    -- CP-element group 89:  members (2) 
      -- CP-element group 89: 	 branch_block_stmt_349/do_while_stmt_350/loop_taken/$exit
      -- CP-element group 89: 	 branch_block_stmt_349/do_while_stmt_350/loop_taken/ack
      -- 
    ack_1087_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_350_branch_ack_1, ack => loadKernelChannel_CP_676_elements(89)); -- 
    -- CP-element group 90:  transition  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	12 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	10 
    -- CP-element group 90:  members (1) 
      -- CP-element group 90: 	 branch_block_stmt_349/do_while_stmt_350/$exit
      -- 
    loadKernelChannel_CP_676_elements(90) <= loadKernelChannel_CP_676_elements(12);
    -- CP-element group 91:  transition  input  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	10 
    -- CP-element group 91: successors 
    -- CP-element group 91:  members (3) 
      -- CP-element group 91: 	 assign_stmt_433/type_cast_432_sample_completed_
      -- CP-element group 91: 	 assign_stmt_433/type_cast_432_Sample/ra
      -- CP-element group 91: 	 assign_stmt_433/type_cast_432_Sample/$exit
      -- 
    ra_1100_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_432_inst_ack_0, ack => loadKernelChannel_CP_676_elements(91)); -- 
    -- CP-element group 92:  transition  input  output  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	10 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	93 
    -- CP-element group 92:  members (6) 
      -- CP-element group 92: 	 assign_stmt_433/type_cast_432_Update/ca
      -- CP-element group 92: 	 assign_stmt_433/WPIPE_size_pipe_428_Sample/$entry
      -- CP-element group 92: 	 assign_stmt_433/WPIPE_size_pipe_428_Sample/req
      -- CP-element group 92: 	 assign_stmt_433/WPIPE_size_pipe_428_sample_start_
      -- CP-element group 92: 	 assign_stmt_433/type_cast_432_update_completed_
      -- CP-element group 92: 	 assign_stmt_433/type_cast_432_Update/$exit
      -- 
    ca_1105_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_432_inst_ack_1, ack => loadKernelChannel_CP_676_elements(92)); -- 
    req_1113_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1113_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(92), ack => WPIPE_size_pipe_428_inst_req_0); -- 
    -- CP-element group 93:  transition  input  output  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	92 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93:  members (6) 
      -- CP-element group 93: 	 assign_stmt_433/WPIPE_size_pipe_428_Sample/$exit
      -- CP-element group 93: 	 assign_stmt_433/WPIPE_size_pipe_428_update_start_
      -- CP-element group 93: 	 assign_stmt_433/WPIPE_size_pipe_428_Sample/ack
      -- CP-element group 93: 	 assign_stmt_433/WPIPE_size_pipe_428_Update/$entry
      -- CP-element group 93: 	 assign_stmt_433/WPIPE_size_pipe_428_sample_completed_
      -- CP-element group 93: 	 assign_stmt_433/WPIPE_size_pipe_428_Update/req
      -- 
    ack_1114_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_size_pipe_428_inst_ack_0, ack => loadKernelChannel_CP_676_elements(93)); -- 
    req_1118_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1118_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_676_elements(93), ack => WPIPE_size_pipe_428_inst_req_1); -- 
    -- CP-element group 94:  transition  input  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94:  members (5) 
      -- CP-element group 94: 	 assign_stmt_433/$exit
      -- CP-element group 94: 	 assign_stmt_433/WPIPE_size_pipe_428_update_completed_
      -- CP-element group 94: 	 assign_stmt_433/WPIPE_size_pipe_428_Update/$exit
      -- CP-element group 94: 	 assign_stmt_433/WPIPE_size_pipe_428_Update/ack
      -- CP-element group 94: 	 $exit
      -- 
    ack_1119_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_size_pipe_428_inst_ack_1, ack => loadKernelChannel_CP_676_elements(94)); -- 
    loadKernelChannel_do_while_stmt_350_terminator_1088: loop_terminator -- 
      generic map (name => " loadKernelChannel_do_while_stmt_350_terminator_1088", max_iterations_in_flight =>15) 
      port map(loop_body_exit => loadKernelChannel_CP_676_elements(15),loop_continue => loadKernelChannel_CP_676_elements(89),loop_terminate => loadKernelChannel_CP_676_elements(88),loop_back => loadKernelChannel_CP_676_elements(13),loop_exit => loadKernelChannel_CP_676_elements(12),clk => clk, reset => reset); -- 
    phi_stmt_352_phi_seq_872_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= loadKernelChannel_CP_676_elements(30);
      loadKernelChannel_CP_676_elements(35)<= src_sample_reqs(0);
      src_sample_acks(0)  <= loadKernelChannel_CP_676_elements(37);
      loadKernelChannel_CP_676_elements(36)<= src_update_reqs(0);
      src_update_acks(0)  <= loadKernelChannel_CP_676_elements(38);
      loadKernelChannel_CP_676_elements(31) <= phi_mux_reqs(0);
      triggers(1)  <= loadKernelChannel_CP_676_elements(32);
      loadKernelChannel_CP_676_elements(39)<= src_sample_reqs(1);
      src_sample_acks(1)  <= loadKernelChannel_CP_676_elements(41);
      loadKernelChannel_CP_676_elements(40)<= src_update_reqs(1);
      src_update_acks(1)  <= loadKernelChannel_CP_676_elements(42);
      loadKernelChannel_CP_676_elements(33) <= phi_mux_reqs(1);
      phi_stmt_352_phi_seq_872 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_352_phi_seq_872") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => loadKernelChannel_CP_676_elements(26), 
          phi_sample_ack => loadKernelChannel_CP_676_elements(27), 
          phi_update_req => loadKernelChannel_CP_676_elements(28), 
          phi_update_ack => loadKernelChannel_CP_676_elements(29), 
          phi_mux_ack => loadKernelChannel_CP_676_elements(34), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_356_phi_seq_926_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= loadKernelChannel_CP_676_elements(47);
      loadKernelChannel_CP_676_elements(52)<= src_sample_reqs(0);
      src_sample_acks(0)  <= loadKernelChannel_CP_676_elements(54);
      loadKernelChannel_CP_676_elements(53)<= src_update_reqs(0);
      src_update_acks(0)  <= loadKernelChannel_CP_676_elements(55);
      loadKernelChannel_CP_676_elements(48) <= phi_mux_reqs(0);
      triggers(1)  <= loadKernelChannel_CP_676_elements(49);
      loadKernelChannel_CP_676_elements(56)<= src_sample_reqs(1);
      src_sample_acks(1)  <= loadKernelChannel_CP_676_elements(58);
      loadKernelChannel_CP_676_elements(57)<= src_update_reqs(1);
      src_update_acks(1)  <= loadKernelChannel_CP_676_elements(59);
      loadKernelChannel_CP_676_elements(50) <= phi_mux_reqs(1);
      phi_stmt_356_phi_seq_926 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_356_phi_seq_926") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => loadKernelChannel_CP_676_elements(20), 
          phi_sample_ack => loadKernelChannel_CP_676_elements(45), 
          phi_update_req => loadKernelChannel_CP_676_elements(22), 
          phi_update_ack => loadKernelChannel_CP_676_elements(46), 
          phi_mux_ack => loadKernelChannel_CP_676_elements(51), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_814_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= loadKernelChannel_CP_676_elements(16);
        preds(1)  <= loadKernelChannel_CP_676_elements(17);
        entry_tmerge_814 : transition_merge -- 
          generic map(name => " entry_tmerge_814")
          port map (preds => preds, symbol_out => loadKernelChannel_CP_676_elements(18));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal AND_u64_u64_365_wire : std_logic_vector(63 downto 0);
    signal AND_u64_u64_387_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_378_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_396_resized : std_logic_vector(13 downto 0);
    signal LSHR_u64_u64_396_scaled : std_logic_vector(13 downto 0);
    signal LSHR_u64_u64_396_wire : std_logic_vector(63 downto 0);
    signal R_sh_start_332_resized : std_logic_vector(13 downto 0);
    signal R_sh_start_332_scaled : std_logic_vector(13 downto 0);
    signal SUB_u64_u64_366_wire : std_logic_vector(63 downto 0);
    signal SUB_u64_u64_424_wire : std_logic_vector(63 downto 0);
    signal SUB_u64_u64_431_wire : std_logic_vector(63 downto 0);
    signal ULT_u64_u1_425_wire : std_logic_vector(0 downto 0);
    signal array_obj_ref_333_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_333_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_333_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_333_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_333_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_333_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_397_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_397_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_397_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_397_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_397_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_397_root_address : std_logic_vector(13 downto 0);
    signal fetch_addr_335 : std_logic_vector(31 downto 0);
    signal fetch_addr_399 : std_logic_vector(31 downto 0);
    signal fetch_val_356 : std_logic_vector(63 downto 0);
    signal fetch_val_396_delayed_13_0_413 : std_logic_vector(63 downto 0);
    signal first_fill_344 : std_logic_vector(0 downto 0);
    signal fn_388_delayed_7_0_402 : std_logic_vector(0 downto 0);
    signal fn_390 : std_logic_vector(0 downto 0);
    signal fn_394_delayed_13_0_410 : std_logic_vector(0 downto 0);
    signal fv_407 : std_logic_vector(63 downto 0);
    signal konst_326_wire_constant : std_logic_vector(63 downto 0);
    signal konst_342_wire_constant : std_logic_vector(63 downto 0);
    signal konst_362_wire_constant : std_logic_vector(63 downto 0);
    signal konst_364_wire_constant : std_logic_vector(63 downto 0);
    signal konst_367_wire_constant : std_logic_vector(63 downto 0);
    signal konst_372_wire_constant : std_logic_vector(63 downto 0);
    signal konst_386_wire_constant : std_logic_vector(63 downto 0);
    signal konst_388_wire_constant : std_logic_vector(63 downto 0);
    signal konst_395_wire_constant : std_logic_vector(63 downto 0);
    signal konst_423_wire_constant : std_logic_vector(63 downto 0);
    signal my_fetch_339 : std_logic_vector(63 downto 0);
    signal my_fetch_339_359_buffered : std_logic_vector(63 downto 0);
    signal my_num1_369 : std_logic_vector(63 downto 0);
    signal mycount_352 : std_logic_vector(63 downto 0);
    signal nfetch_val_419 : std_logic_vector(63 downto 0);
    signal nfetch_val_419_358_buffered : std_logic_vector(63 downto 0);
    signal nmycount_374 : std_logic_vector(63 downto 0);
    signal nmycount_374_354_buffered : std_logic_vector(63 downto 0);
    signal ptr_deref_338_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_338_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_338_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_338_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_338_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_406_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_406_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_406_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_406_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_406_word_offset_0 : std_logic_vector(13 downto 0);
    signal sh_start_328 : std_logic_vector(63 downto 0);
    signal start_add_355_buffered : std_logic_vector(63 downto 0);
    signal start_next_348 : std_logic_vector(0 downto 0);
    signal type_cast_432_wire : std_logic_vector(31 downto 0);
    signal var_val_380 : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_333_constant_part_of_offset <= "00000000000000";
    array_obj_ref_333_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_333_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_333_resized_base_address <= "00000000000000";
    array_obj_ref_397_constant_part_of_offset <= "00000000000000";
    array_obj_ref_397_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_397_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_397_resized_base_address <= "00000000000000";
    konst_326_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    konst_342_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    konst_362_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_364_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_367_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000100";
    konst_372_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    konst_386_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_388_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    konst_395_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    konst_423_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    ptr_deref_338_word_offset_0 <= "00000000000000";
    ptr_deref_406_word_offset_0 <= "00000000000000";
    phi_stmt_352: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= nmycount_374_354_buffered & start_add_355_buffered;
      req <= phi_stmt_352_req_0 & phi_stmt_352_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_352",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_352_ack_0,
          idata => idata,
          odata => mycount_352,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_352
    phi_stmt_356: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= nfetch_val_419_358_buffered & my_fetch_339_359_buffered;
      req <= phi_stmt_356_req_0 & phi_stmt_356_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_356",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_356_ack_0,
          idata => idata,
          odata => fetch_val_356,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_356
    -- flow-through select operator MUX_418_inst
    nfetch_val_419 <= fv_407 when (fn_394_delayed_13_0_410(0) /=  '0') else fetch_val_396_delayed_13_0_413;
    W_fetch_val_396_delayed_13_0_411_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fetch_val_396_delayed_13_0_411_inst_req_0;
      W_fetch_val_396_delayed_13_0_411_inst_ack_0<= wack(0);
      rreq(0) <= W_fetch_val_396_delayed_13_0_411_inst_req_1;
      W_fetch_val_396_delayed_13_0_411_inst_ack_1<= rack(0);
      W_fetch_val_396_delayed_13_0_411_inst : InterlockBuffer generic map ( -- 
        name => "W_fetch_val_396_delayed_13_0_411_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fetch_val_356,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_val_396_delayed_13_0_413,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fn_388_delayed_7_0_400_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fn_388_delayed_7_0_400_inst_req_0;
      W_fn_388_delayed_7_0_400_inst_ack_0<= wack(0);
      rreq(0) <= W_fn_388_delayed_7_0_400_inst_req_1;
      W_fn_388_delayed_7_0_400_inst_ack_1<= rack(0);
      W_fn_388_delayed_7_0_400_inst : InterlockBuffer generic map ( -- 
        name => "W_fn_388_delayed_7_0_400_inst",
        buffer_size => 7,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fn_390,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fn_388_delayed_7_0_402,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fn_394_delayed_13_0_408_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fn_394_delayed_13_0_408_inst_req_0;
      W_fn_394_delayed_13_0_408_inst_ack_0<= wack(0);
      rreq(0) <= W_fn_394_delayed_13_0_408_inst_req_1;
      W_fn_394_delayed_13_0_408_inst_ack_1<= rack(0);
      W_fn_394_delayed_13_0_408_inst : InterlockBuffer generic map ( -- 
        name => "W_fn_394_delayed_13_0_408_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fn_390,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fn_394_delayed_13_0_410,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_334_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_334_final_reg_req_0;
      addr_of_334_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_334_final_reg_req_1;
      addr_of_334_final_reg_ack_1<= rack(0);
      addr_of_334_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_334_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_333_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr_335,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_398_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_398_final_reg_req_0;
      addr_of_398_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_398_final_reg_req_1;
      addr_of_398_final_reg_ack_1<= rack(0);
      addr_of_398_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_398_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_397_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr_399,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    my_fetch_339_359_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= my_fetch_339_359_buf_req_0;
      my_fetch_339_359_buf_ack_0<= wack(0);
      rreq(0) <= my_fetch_339_359_buf_req_1;
      my_fetch_339_359_buf_ack_1<= rack(0);
      my_fetch_339_359_buf : InterlockBuffer generic map ( -- 
        name => "my_fetch_339_359_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => my_fetch_339,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => my_fetch_339_359_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nfetch_val_419_358_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nfetch_val_419_358_buf_req_0;
      nfetch_val_419_358_buf_ack_0<= wack(0);
      rreq(0) <= nfetch_val_419_358_buf_req_1;
      nfetch_val_419_358_buf_ack_1<= rack(0);
      nfetch_val_419_358_buf : InterlockBuffer generic map ( -- 
        name => "nfetch_val_419_358_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nfetch_val_419,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nfetch_val_419_358_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nmycount_374_354_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nmycount_374_354_buf_req_0;
      nmycount_374_354_buf_ack_0<= wack(0);
      rreq(0) <= nmycount_374_354_buf_req_1;
      nmycount_374_354_buf_ack_1<= rack(0);
      nmycount_374_354_buf : InterlockBuffer generic map ( -- 
        name => "nmycount_374_354_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nmycount_374,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nmycount_374_354_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    start_add_355_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= start_add_355_buf_req_0;
      start_add_355_buf_ack_0<= wack(0);
      rreq(0) <= start_add_355_buf_req_1;
      start_add_355_buf_ack_1<= rack(0);
      start_add_355_buf : InterlockBuffer generic map ( -- 
        name => "start_add_355_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => start_add_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => start_add_355_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_379_inst
    process(LSHR_u64_u64_378_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := LSHR_u64_u64_378_wire(15 downto 0);
      var_val_380 <= tmp_var; -- 
    end process;
    type_cast_432_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_432_inst_req_0;
      type_cast_432_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_432_inst_req_1;
      type_cast_432_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  first_fill_344(0);
      type_cast_432_inst_gI: SplitGuardInterface generic map(name => "type_cast_432_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_432_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_432_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => SUB_u64_u64_431_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_432_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_333_index_1_rename
    process(R_sh_start_332_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_sh_start_332_resized;
      ov(13 downto 0) := iv;
      R_sh_start_332_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_333_index_1_resize
    process(sh_start_328) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := sh_start_328;
      ov := iv(13 downto 0);
      R_sh_start_332_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_333_root_address_inst
    process(array_obj_ref_333_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_333_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_333_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_397_index_1_rename
    process(LSHR_u64_u64_396_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LSHR_u64_u64_396_resized;
      ov(13 downto 0) := iv;
      LSHR_u64_u64_396_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_397_index_1_resize
    process(LSHR_u64_u64_396_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LSHR_u64_u64_396_wire;
      ov := iv(13 downto 0);
      LSHR_u64_u64_396_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_397_root_address_inst
    process(array_obj_ref_397_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_397_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_397_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_338_addr_0
    process(ptr_deref_338_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_338_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_338_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_338_base_resize
    process(fetch_addr_335) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr_335;
      ov := iv(13 downto 0);
      ptr_deref_338_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_338_gather_scatter
    process(ptr_deref_338_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_338_data_0;
      ov(63 downto 0) := iv;
      my_fetch_339 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_338_root_address_inst
    process(ptr_deref_338_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_338_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_338_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_406_addr_0
    process(ptr_deref_406_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_406_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_406_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_406_base_resize
    process(fetch_addr_399) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr_399;
      ov := iv(13 downto 0);
      ptr_deref_406_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_406_gather_scatter
    process(ptr_deref_406_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_406_data_0;
      ov(63 downto 0) := iv;
      fv_407 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_406_root_address_inst
    process(ptr_deref_406_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_406_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_406_root_address <= ov(13 downto 0);
      --
    end process;
    do_while_stmt_350_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= ULT_u64_u1_425_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_350_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_350_branch_req_0,
          ack0 => do_while_stmt_350_branch_ack_0,
          ack1 => do_while_stmt_350_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u64_u64_373_inst
    process(mycount_352) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mycount_352, konst_372_wire_constant, tmp_var);
      nmycount_374 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_365_inst
    process(mycount_352) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(mycount_352, konst_364_wire_constant, tmp_var);
      AND_u64_u64_365_wire <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_387_inst
    process(nmycount_374) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(nmycount_374, konst_386_wire_constant, tmp_var);
      AND_u64_u64_387_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_343_inst
    process(start_add_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(start_add_buffer, konst_342_wire_constant, tmp_var);
      first_fill_344 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_389_inst
    process(AND_u64_u64_387_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(AND_u64_u64_387_wire, konst_388_wire_constant, tmp_var);
      fn_390 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_327_inst
    process(start_add_buffer) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(start_add_buffer, konst_326_wire_constant, tmp_var);
      sh_start_328 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_378_inst
    process(fetch_val_356, my_num1_369) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(fetch_val_356, my_num1_369, tmp_var);
      LSHR_u64_u64_378_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_396_inst
    process(nmycount_374) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(nmycount_374, konst_395_wire_constant, tmp_var);
      LSHR_u64_u64_396_wire <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_368_inst
    process(SUB_u64_u64_366_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(SUB_u64_u64_366_wire, konst_367_wire_constant, tmp_var);
      my_num1_369 <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_366_inst
    process(konst_362_wire_constant, AND_u64_u64_365_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(konst_362_wire_constant, AND_u64_u64_365_wire, tmp_var);
      SUB_u64_u64_366_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_424_inst
    process(end_add_buffer) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(end_add_buffer, konst_423_wire_constant, tmp_var);
      SUB_u64_u64_424_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_431_inst
    process(end_add_buffer, start_add_buffer) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(end_add_buffer, start_add_buffer, tmp_var);
      SUB_u64_u64_431_wire <= tmp_var; --
    end process;
    -- binary operator ULT_u64_u1_425_inst
    process(mycount_352, SUB_u64_u64_424_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(mycount_352, SUB_u64_u64_424_wire, tmp_var);
      ULT_u64_u1_425_wire <= tmp_var; --
    end process;
    -- shared split operator group (13) : array_obj_ref_333_index_offset 
    ApIntAdd_group_13: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_sh_start_332_scaled;
      array_obj_ref_333_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_333_index_offset_req_0;
      array_obj_ref_333_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_333_index_offset_req_1;
      array_obj_ref_333_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_13_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_13_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_13",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 13
    -- shared split operator group (14) : array_obj_ref_397_index_offset 
    ApIntAdd_group_14: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= LSHR_u64_u64_396_scaled;
      array_obj_ref_397_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_397_index_offset_req_0;
      array_obj_ref_397_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_397_index_offset_req_1;
      array_obj_ref_397_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_14_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_14_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_14",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 14
    -- shared load operator group (0) : ptr_deref_338_load_0 ptr_deref_406_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(27 downto 0);
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 2);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 2);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => true, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 6, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_338_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_406_load_0_req_0;
      ptr_deref_338_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_406_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_338_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_406_load_0_req_1;
      ptr_deref_338_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_406_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= fn_388_delayed_7_0_402(0);
      guard_vector(1)  <=  '1';
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 2) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_338_word_address_0 & ptr_deref_406_word_address_0;
      ptr_deref_338_data_0 <= data_out(127 downto 64);
      ptr_deref_406_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(13 downto 0),
          mtag => memory_space_0_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared inport operator group (0) : RPIPE_input_done_pipe_347_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(0 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_input_done_pipe_347_inst_req_0;
      RPIPE_input_done_pipe_347_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_input_done_pipe_347_inst_req_1;
      RPIPE_input_done_pipe_347_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not first_fill_344(0);
      start_next_348 <= data_out(0 downto 0);
      input_done_pipe_read_0_gI: SplitGuardInterface generic map(name => "input_done_pipe_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      input_done_pipe_read_0: InputPortRevised -- 
        generic map ( name => "input_done_pipe_read_0", data_width => 1,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => input_done_pipe_pipe_read_req(0),
          oack => input_done_pipe_pipe_read_ack(0),
          odata => input_done_pipe_pipe_read_data(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_kernel_pipe1_381_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_kernel_pipe1_381_inst_req_0;
      WPIPE_kernel_pipe1_381_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_kernel_pipe1_381_inst_req_1;
      WPIPE_kernel_pipe1_381_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= var_val_380;
      kernel_pipe1_write_0_gI: SplitGuardInterface generic map(name => "kernel_pipe1_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      kernel_pipe1_write_0: OutputPortRevised -- 
        generic map ( name => "kernel_pipe1", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => kernel_pipe1_pipe_write_req(0),
          oack => kernel_pipe1_pipe_write_ack(0),
          odata => kernel_pipe1_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_size_pipe_428_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_size_pipe_428_inst_req_0;
      WPIPE_size_pipe_428_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_size_pipe_428_inst_req_1;
      WPIPE_size_pipe_428_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= first_fill_344(0);
      data_in <= type_cast_432_wire;
      size_pipe_write_1_gI: SplitGuardInterface generic map(name => "size_pipe_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      size_pipe_write_1: OutputPortRevised -- 
        generic map ( name => "size_pipe", data_width => 32, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => size_pipe_pipe_write_req(0),
          oack => size_pipe_pipe_write_ack(0),
          odata => size_pipe_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- 
  end Block; -- data_path
  -- 
end loadKernelChannel_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timer is -- 
  generic (tag_length : integer); 
  port ( -- 
    c : out  std_logic_vector(63 downto 0);
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timer;
architecture timer_arch of timer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal c_buffer :  std_logic_vector(63 downto 0);
  signal c_update_enable: Boolean;
  signal timer_CP_637_start: Boolean;
  signal timer_CP_637_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal LOAD_count_318_load_0_req_0 : boolean;
  signal LOAD_count_318_load_0_ack_0 : boolean;
  signal LOAD_count_318_load_0_req_1 : boolean;
  signal LOAD_count_318_load_0_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timer_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timer_CP_637_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timer_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= c_buffer;
  c <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_637_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timer_CP_637_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_637_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timer_CP_637: Block -- control-path 
    signal timer_CP_637_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    timer_CP_637_elements(0) <= timer_CP_637_start;
    timer_CP_637_symbol <= timer_CP_637_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_319/$entry
      -- CP-element group 0: 	 assign_stmt_319/LOAD_count_318_sample_start_
      -- CP-element group 0: 	 assign_stmt_319/LOAD_count_318_update_start_
      -- CP-element group 0: 	 assign_stmt_319/LOAD_count_318_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_319/LOAD_count_318_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_319/LOAD_count_318_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_319/LOAD_count_318_Sample/word_access_start/$entry
      -- CP-element group 0: 	 assign_stmt_319/LOAD_count_318_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_319/LOAD_count_318_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 assign_stmt_319/LOAD_count_318_Update/$entry
      -- CP-element group 0: 	 assign_stmt_319/LOAD_count_318_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_319/LOAD_count_318_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_319/LOAD_count_318_Update/word_access_complete/word_0/cr
      -- 
    cr_669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_637_elements(0), ack => LOAD_count_318_load_0_req_1); -- 
    rr_658_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_658_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_637_elements(0), ack => LOAD_count_318_load_0_req_0); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (5) 
      -- CP-element group 1: 	 assign_stmt_319/LOAD_count_318_sample_completed_
      -- CP-element group 1: 	 assign_stmt_319/LOAD_count_318_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_319/LOAD_count_318_Sample/word_access_start/$exit
      -- CP-element group 1: 	 assign_stmt_319/LOAD_count_318_Sample/word_access_start/word_0/$exit
      -- CP-element group 1: 	 assign_stmt_319/LOAD_count_318_Sample/word_access_start/word_0/ra
      -- 
    ra_659_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_count_318_load_0_ack_0, ack => timer_CP_637_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (11) 
      -- CP-element group 2: 	 $exit
      -- CP-element group 2: 	 assign_stmt_319/$exit
      -- CP-element group 2: 	 assign_stmt_319/LOAD_count_318_update_completed_
      -- CP-element group 2: 	 assign_stmt_319/LOAD_count_318_Update/$exit
      -- CP-element group 2: 	 assign_stmt_319/LOAD_count_318_Update/word_access_complete/$exit
      -- CP-element group 2: 	 assign_stmt_319/LOAD_count_318_Update/word_access_complete/word_0/$exit
      -- CP-element group 2: 	 assign_stmt_319/LOAD_count_318_Update/word_access_complete/word_0/ca
      -- CP-element group 2: 	 assign_stmt_319/LOAD_count_318_Update/LOAD_count_318_Merge/$entry
      -- CP-element group 2: 	 assign_stmt_319/LOAD_count_318_Update/LOAD_count_318_Merge/$exit
      -- CP-element group 2: 	 assign_stmt_319/LOAD_count_318_Update/LOAD_count_318_Merge/merge_req
      -- CP-element group 2: 	 assign_stmt_319/LOAD_count_318_Update/LOAD_count_318_Merge/merge_ack
      -- 
    ca_670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_count_318_load_0_ack_1, ack => timer_CP_637_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal LOAD_count_318_data_0 : std_logic_vector(63 downto 0);
    signal LOAD_count_318_word_address_0 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    LOAD_count_318_word_address_0 <= "0";
    -- equivalence LOAD_count_318_gather_scatter
    process(LOAD_count_318_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_count_318_data_0;
      ov(63 downto 0) := iv;
      c_buffer <= ov(63 downto 0);
      --
    end process;
    -- shared load operator group (0) : LOAD_count_318_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_count_318_load_0_req_0;
      LOAD_count_318_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_count_318_load_0_req_1;
      LOAD_count_318_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_count_318_word_address_0;
      LOAD_count_318_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(0 downto 0),
          mtag => memory_space_2_lr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(63 downto 0),
          mtag => memory_space_2_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- 
  end Block; -- data_path
  -- 
end timer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timerDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timerDaemon;
architecture timerDaemon_arch of timerDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal timerDaemon_CP_5052_start: Boolean;
  signal timerDaemon_CP_5052_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal do_while_stmt_2102_branch_req_0 : boolean;
  signal phi_stmt_2104_req_1 : boolean;
  signal phi_stmt_2104_req_0 : boolean;
  signal phi_stmt_2104_ack_0 : boolean;
  signal ADD_u64_u64_2110_inst_req_0 : boolean;
  signal ADD_u64_u64_2110_inst_ack_0 : boolean;
  signal ADD_u64_u64_2110_inst_req_1 : boolean;
  signal ADD_u64_u64_2110_inst_ack_1 : boolean;
  signal STORE_count_2112_store_0_req_0 : boolean;
  signal STORE_count_2112_store_0_ack_0 : boolean;
  signal STORE_count_2112_store_0_req_1 : boolean;
  signal STORE_count_2112_store_0_ack_1 : boolean;
  signal do_while_stmt_2102_branch_ack_0 : boolean;
  signal do_while_stmt_2102_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timerDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timerDaemon_CP_5052_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timerDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timerDaemon_CP_5052_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timerDaemon_CP_5052_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timerDaemon_CP_5052_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timerDaemon_CP_5052: Block -- control-path 
    signal timerDaemon_CP_5052_elements: BooleanArray(39 downto 0);
    -- 
  begin -- 
    timerDaemon_CP_5052_elements(0) <= timerDaemon_CP_5052_start;
    timerDaemon_CP_5052_symbol <= timerDaemon_CP_5052_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_2101/$entry
      -- CP-element group 0: 	 branch_block_stmt_2101/branch_block_stmt_2101__entry__
      -- CP-element group 0: 	 branch_block_stmt_2101/do_while_stmt_2102__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	39 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_2101/$exit
      -- CP-element group 1: 	 branch_block_stmt_2101/branch_block_stmt_2101__exit__
      -- CP-element group 1: 	 branch_block_stmt_2101/do_while_stmt_2102__exit__
      -- 
    timerDaemon_CP_5052_elements(1) <= timerDaemon_CP_5052_elements(39);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_2101/do_while_stmt_2102/$entry
      -- CP-element group 2: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102__entry__
      -- 
    timerDaemon_CP_5052_elements(2) <= timerDaemon_CP_5052_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	39 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102__exit__
      -- 
    -- Element group timerDaemon_CP_5052_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_2101/do_while_stmt_2102/loop_back
      -- 
    -- Element group timerDaemon_CP_5052_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	37 
    -- CP-element group 5: 	38 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_2101/do_while_stmt_2102/condition_done
      -- CP-element group 5: 	 branch_block_stmt_2101/do_while_stmt_2102/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_2101/do_while_stmt_2102/loop_taken/$entry
      -- 
    timerDaemon_CP_5052_elements(5) <= timerDaemon_CP_5052_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	36 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_2101/do_while_stmt_2102/loop_body_done
      -- 
    timerDaemon_CP_5052_elements(6) <= timerDaemon_CP_5052_elements(36);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	16 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/back_edge_to_loop_body
      -- 
    timerDaemon_CP_5052_elements(7) <= timerDaemon_CP_5052_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	18 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/first_time_through_loop_body
      -- 
    timerDaemon_CP_5052_elements(8) <= timerDaemon_CP_5052_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	12 
    -- CP-element group 9: 	13 
    -- CP-element group 9: 	31 
    -- CP-element group 9: 	35 
    -- CP-element group 9:  members (4) 
      -- CP-element group 9: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/STORE_count_2112_word_address_calculated
      -- CP-element group 9: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/STORE_count_2112_root_address_calculated
      -- 
    -- Element group timerDaemon_CP_5052_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	35 
    -- CP-element group 10: 	15 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/condition_evaluated
      -- 
    condition_evaluated_5076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_5076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_5052_elements(10), ack => do_while_stmt_2102_branch_req_0); -- 
    timerDaemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 3);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_5052_elements(35) & timerDaemon_CP_5052_elements(15);
      gj_timerDaemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_5052_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	12 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	15 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/phi_stmt_2104_sample_start__ps
      -- 
    timerDaemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_5052_elements(12) & timerDaemon_CP_5052_elements(15);
      gj_timerDaemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_5052_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	9 
    -- CP-element group 12: marked-predecessors 
    -- CP-element group 12: 	14 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	11 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/phi_stmt_2104_sample_start_
      -- 
    timerDaemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_5052_elements(9) & timerDaemon_CP_5052_elements(14);
      gj_timerDaemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_5052_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	9 
    -- CP-element group 13: marked-predecessors 
    -- CP-element group 13: 	33 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/phi_stmt_2104_update_start_
      -- CP-element group 13: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/phi_stmt_2104_update_start__ps
      -- 
    timerDaemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_5052_elements(9) & timerDaemon_CP_5052_elements(33);
      gj_timerDaemon_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_5052_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	36 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	12 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/aggregated_phi_sample_ack
      -- CP-element group 14: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/phi_stmt_2104_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/phi_stmt_2104_sample_completed__ps
      -- 
    -- Element group timerDaemon_CP_5052_elements(14) is bound as output of CP function.
    -- CP-element group 15:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	10 
    -- CP-element group 15: 	31 
    -- CP-element group 15: marked-successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/aggregated_phi_update_ack
      -- CP-element group 15: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/phi_stmt_2104_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/phi_stmt_2104_update_completed__ps
      -- 
    -- Element group timerDaemon_CP_5052_elements(15) is bound as output of CP function.
    -- CP-element group 16:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	7 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/phi_stmt_2104_loopback_trigger
      -- 
    timerDaemon_CP_5052_elements(16) <= timerDaemon_CP_5052_elements(7);
    -- CP-element group 17:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (2) 
      -- CP-element group 17: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/phi_stmt_2104_loopback_sample_req
      -- CP-element group 17: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/phi_stmt_2104_loopback_sample_req_ps
      -- 
    phi_stmt_2104_loopback_sample_req_5091_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2104_loopback_sample_req_5091_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_5052_elements(17), ack => phi_stmt_2104_req_1); -- 
    -- Element group timerDaemon_CP_5052_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	8 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/phi_stmt_2104_entry_trigger
      -- 
    timerDaemon_CP_5052_elements(18) <= timerDaemon_CP_5052_elements(8);
    -- CP-element group 19:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (2) 
      -- CP-element group 19: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/phi_stmt_2104_entry_sample_req
      -- CP-element group 19: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/phi_stmt_2104_entry_sample_req_ps
      -- 
    phi_stmt_2104_entry_sample_req_5094_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2104_entry_sample_req_5094_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_5052_elements(19), ack => phi_stmt_2104_req_0); -- 
    -- Element group timerDaemon_CP_5052_elements(19) is bound as output of CP function.
    -- CP-element group 20:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/phi_stmt_2104_phi_mux_ack
      -- CP-element group 20: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/phi_stmt_2104_phi_mux_ack_ps
      -- 
    phi_stmt_2104_phi_mux_ack_5097_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2104_ack_0, ack => timerDaemon_CP_5052_elements(20)); -- 
    -- CP-element group 21:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (4) 
      -- CP-element group 21: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/type_cast_2107_sample_start__ps
      -- CP-element group 21: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/type_cast_2107_sample_completed__ps
      -- CP-element group 21: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/type_cast_2107_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/type_cast_2107_sample_completed_
      -- 
    -- Element group timerDaemon_CP_5052_elements(21) is bound as output of CP function.
    -- CP-element group 22:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	24 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/type_cast_2107_update_start__ps
      -- CP-element group 22: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/type_cast_2107_update_start_
      -- 
    -- Element group timerDaemon_CP_5052_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	24 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/type_cast_2107_update_completed__ps
      -- 
    timerDaemon_CP_5052_elements(23) <= timerDaemon_CP_5052_elements(24);
    -- CP-element group 24:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	22 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	23 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/type_cast_2107_update_completed_
      -- 
    -- Element group timerDaemon_CP_5052_elements(24) is a control-delay.
    cp_element_24_delay: control_delay_element  generic map(name => " 24_delay", delay_value => 1)  port map(req => timerDaemon_CP_5052_elements(22), ack => timerDaemon_CP_5052_elements(24), clk => clk, reset =>reset);
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/ADD_u64_u64_2110_sample_start__ps
      -- 
    -- Element group timerDaemon_CP_5052_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	28 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/ADD_u64_u64_2110_update_start__ps
      -- 
    -- Element group timerDaemon_CP_5052_elements(26) is bound as output of CP function.
    -- CP-element group 27:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: marked-predecessors 
    -- CP-element group 27: 	29 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/ADD_u64_u64_2110_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/ADD_u64_u64_2110_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/ADD_u64_u64_2110_Sample/rr
      -- 
    rr_5118_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5118_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_5052_elements(27), ack => ADD_u64_u64_2110_inst_req_0); -- 
    timerDaemon_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_5052_elements(25) & timerDaemon_CP_5052_elements(29);
      gj_timerDaemon_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_5052_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: marked-predecessors 
    -- CP-element group 28: 	30 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/ADD_u64_u64_2110_update_start_
      -- CP-element group 28: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/ADD_u64_u64_2110_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/ADD_u64_u64_2110_Update/cr
      -- 
    cr_5123_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5123_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_5052_elements(28), ack => ADD_u64_u64_2110_inst_req_1); -- 
    timerDaemon_cp_element_group_28: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_28"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_5052_elements(26) & timerDaemon_CP_5052_elements(30);
      gj_timerDaemon_cp_element_group_28 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_5052_elements(28), clk => clk, reset => reset); --
    end block;
    -- CP-element group 29:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29: marked-successors 
    -- CP-element group 29: 	27 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/ADD_u64_u64_2110_sample_completed__ps
      -- CP-element group 29: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/ADD_u64_u64_2110_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/ADD_u64_u64_2110_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/ADD_u64_u64_2110_Sample/ra
      -- 
    ra_5119_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_2110_inst_ack_0, ack => timerDaemon_CP_5052_elements(29)); -- 
    -- CP-element group 30:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30: marked-successors 
    -- CP-element group 30: 	28 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/ADD_u64_u64_2110_update_completed__ps
      -- CP-element group 30: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/ADD_u64_u64_2110_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/ADD_u64_u64_2110_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/ADD_u64_u64_2110_Update/ca
      -- 
    ca_5124_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_2110_inst_ack_1, ack => timerDaemon_CP_5052_elements(30)); -- 
    -- CP-element group 31:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	9 
    -- CP-element group 31: 	15 
    -- CP-element group 31: marked-predecessors 
    -- CP-element group 31: 	33 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (9) 
      -- CP-element group 31: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/STORE_count_2112_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/STORE_count_2112_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/STORE_count_2112_Sample/STORE_count_2112_Split/$entry
      -- CP-element group 31: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/STORE_count_2112_Sample/STORE_count_2112_Split/$exit
      -- CP-element group 31: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/STORE_count_2112_Sample/STORE_count_2112_Split/split_req
      -- CP-element group 31: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/STORE_count_2112_Sample/STORE_count_2112_Split/split_ack
      -- CP-element group 31: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/STORE_count_2112_Sample/word_access_start/$entry
      -- CP-element group 31: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/STORE_count_2112_Sample/word_access_start/word_0/$entry
      -- CP-element group 31: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/STORE_count_2112_Sample/word_access_start/word_0/rr
      -- 
    rr_5146_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5146_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_5052_elements(31), ack => STORE_count_2112_store_0_req_0); -- 
    timerDaemon_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 3,1 => 3,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= timerDaemon_CP_5052_elements(9) & timerDaemon_CP_5052_elements(15) & timerDaemon_CP_5052_elements(33);
      gj_timerDaemon_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_5052_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	34 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	34 
    -- CP-element group 32:  members (5) 
      -- CP-element group 32: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/STORE_count_2112_update_start_
      -- CP-element group 32: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/STORE_count_2112_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/STORE_count_2112_Update/word_access_complete/$entry
      -- CP-element group 32: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/STORE_count_2112_Update/word_access_complete/word_0/$entry
      -- CP-element group 32: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/STORE_count_2112_Update/word_access_complete/word_0/cr
      -- 
    cr_5157_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5157_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_5052_elements(32), ack => STORE_count_2112_store_0_req_1); -- 
    timerDaemon_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= timerDaemon_CP_5052_elements(34);
      gj_timerDaemon_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_5052_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33: marked-successors 
    -- CP-element group 33: 	13 
    -- CP-element group 33: 	31 
    -- CP-element group 33:  members (5) 
      -- CP-element group 33: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/STORE_count_2112_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/STORE_count_2112_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/STORE_count_2112_Sample/word_access_start/$exit
      -- CP-element group 33: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/STORE_count_2112_Sample/word_access_start/word_0/$exit
      -- CP-element group 33: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/STORE_count_2112_Sample/word_access_start/word_0/ra
      -- 
    ra_5147_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_count_2112_store_0_ack_0, ack => timerDaemon_CP_5052_elements(33)); -- 
    -- CP-element group 34:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	32 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34: marked-successors 
    -- CP-element group 34: 	32 
    -- CP-element group 34:  members (5) 
      -- CP-element group 34: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/STORE_count_2112_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/STORE_count_2112_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/STORE_count_2112_Update/word_access_complete/$exit
      -- CP-element group 34: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/STORE_count_2112_Update/word_access_complete/word_0/$exit
      -- CP-element group 34: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/STORE_count_2112_Update/word_access_complete/word_0/ca
      -- 
    ca_5158_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_count_2112_store_0_ack_1, ack => timerDaemon_CP_5052_elements(34)); -- 
    -- CP-element group 35:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	9 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	10 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group timerDaemon_CP_5052_elements(35) is a control-delay.
    cp_element_35_delay: control_delay_element  generic map(name => " 35_delay", delay_value => 1)  port map(req => timerDaemon_CP_5052_elements(9), ack => timerDaemon_CP_5052_elements(35), clk => clk, reset =>reset);
    -- CP-element group 36:  join  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: 	14 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	6 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/$exit
      -- 
    timerDaemon_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 3);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_5052_elements(34) & timerDaemon_CP_5052_elements(14);
      gj_timerDaemon_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_5052_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  transition  input  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	5 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (2) 
      -- CP-element group 37: 	 branch_block_stmt_2101/do_while_stmt_2102/loop_exit/$exit
      -- CP-element group 37: 	 branch_block_stmt_2101/do_while_stmt_2102/loop_exit/ack
      -- 
    ack_5163_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_2102_branch_ack_0, ack => timerDaemon_CP_5052_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	5 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (2) 
      -- CP-element group 38: 	 branch_block_stmt_2101/do_while_stmt_2102/loop_taken/$exit
      -- CP-element group 38: 	 branch_block_stmt_2101/do_while_stmt_2102/loop_taken/ack
      -- 
    ack_5167_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_2102_branch_ack_1, ack => timerDaemon_CP_5052_elements(38)); -- 
    -- CP-element group 39:  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	3 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	1 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_2101/do_while_stmt_2102/$exit
      -- 
    timerDaemon_CP_5052_elements(39) <= timerDaemon_CP_5052_elements(3);
    timerDaemon_do_while_stmt_2102_terminator_5168: loop_terminator -- 
      generic map (name => " timerDaemon_do_while_stmt_2102_terminator_5168", max_iterations_in_flight =>3) 
      port map(loop_body_exit => timerDaemon_CP_5052_elements(6),loop_continue => timerDaemon_CP_5052_elements(38),loop_terminate => timerDaemon_CP_5052_elements(37),loop_back => timerDaemon_CP_5052_elements(4),loop_exit => timerDaemon_CP_5052_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_2104_phi_seq_5125_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= timerDaemon_CP_5052_elements(18);
      timerDaemon_CP_5052_elements(21)<= src_sample_reqs(0);
      src_sample_acks(0)  <= timerDaemon_CP_5052_elements(21);
      timerDaemon_CP_5052_elements(22)<= src_update_reqs(0);
      src_update_acks(0)  <= timerDaemon_CP_5052_elements(23);
      timerDaemon_CP_5052_elements(19) <= phi_mux_reqs(0);
      triggers(1)  <= timerDaemon_CP_5052_elements(16);
      timerDaemon_CP_5052_elements(25)<= src_sample_reqs(1);
      src_sample_acks(1)  <= timerDaemon_CP_5052_elements(29);
      timerDaemon_CP_5052_elements(26)<= src_update_reqs(1);
      src_update_acks(1)  <= timerDaemon_CP_5052_elements(30);
      timerDaemon_CP_5052_elements(17) <= phi_mux_reqs(1);
      phi_stmt_2104_phi_seq_5125 : phi_sequencer_v2-- 
        generic map (place_capacity => 3, ntriggers => 2, name => "phi_stmt_2104_phi_seq_5125") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => timerDaemon_CP_5052_elements(11), 
          phi_sample_ack => timerDaemon_CP_5052_elements(14), 
          phi_update_req => timerDaemon_CP_5052_elements(13), 
          phi_update_ack => timerDaemon_CP_5052_elements(15), 
          phi_mux_ack => timerDaemon_CP_5052_elements(20), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_5077_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= timerDaemon_CP_5052_elements(7);
        preds(1)  <= timerDaemon_CP_5052_elements(8);
        entry_tmerge_5077 : transition_merge -- 
          generic map(name => " entry_tmerge_5077")
          port map (preds => preds, symbol_out => timerDaemon_CP_5052_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u64_u64_2110_wire : std_logic_vector(63 downto 0);
    signal STORE_count_2112_data_0 : std_logic_vector(63 downto 0);
    signal STORE_count_2112_word_address_0 : std_logic_vector(0 downto 0);
    signal konst_2109_wire_constant : std_logic_vector(63 downto 0);
    signal konst_2116_wire_constant : std_logic_vector(0 downto 0);
    signal ncount_2104 : std_logic_vector(63 downto 0);
    signal type_cast_2107_wire_constant : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    STORE_count_2112_word_address_0 <= "0";
    konst_2109_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    konst_2116_wire_constant <= "1";
    type_cast_2107_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    phi_stmt_2104: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2107_wire_constant & ADD_u64_u64_2110_wire;
      req <= phi_stmt_2104_req_0 & phi_stmt_2104_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2104",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2104_ack_0,
          idata => idata,
          odata => ncount_2104,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2104
    -- equivalence STORE_count_2112_gather_scatter
    process(ncount_2104) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ncount_2104;
      ov(63 downto 0) := iv;
      STORE_count_2112_data_0 <= ov(63 downto 0);
      --
    end process;
    do_while_stmt_2102_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_2116_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_2102_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_2102_branch_req_0,
          ack0 => do_while_stmt_2102_branch_ack_0,
          ack1 => do_while_stmt_2102_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : ADD_u64_u64_2110_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ncount_2104;
      ADD_u64_u64_2110_wire <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u64_u64_2110_inst_req_0;
      ADD_u64_u64_2110_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u64_u64_2110_inst_req_1;
      ADD_u64_u64_2110_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000000001",
          constant_width => 64,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared store operator group (0) : STORE_count_2112_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 3);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= STORE_count_2112_store_0_req_0;
      STORE_count_2112_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= STORE_count_2112_store_0_req_1;
      STORE_count_2112_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_count_2112_word_address_0;
      data_in <= STORE_count_2112_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 1,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(0 downto 0),
          mdata => memory_space_2_sr_data(63 downto 0),
          mtag => memory_space_2_sr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end timerDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    elapsed_time_pipe_pipe_read_data: out std_logic_vector(63 downto 0);
    elapsed_time_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_read_ack : out std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_write_data: in std_logic_vector(7 downto 0);
    maxpool_input_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_read_data: out std_logic_vector(7 downto 0);
    maxpool_output_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(18 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(1 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(18 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(1 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_2_lr_tag : std_logic_vector(17 downto 0);
  signal memory_space_2_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_2_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(17 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(0 downto 0);
  -- declarations related to module access_T
  component access_T is -- 
    generic (tag_length : integer); 
    port ( -- 
      num_cont : in  std_logic_vector(15 downto 0);
      row1 : in  std_logic_vector(15 downto 0);
      col1 : in  std_logic_vector(15 downto 0);
      rk1 : in  std_logic_vector(15 downto 0);
      chl_in : in  std_logic_vector(15 downto 0);
      ct : in  std_logic_vector(15 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
      input_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module access_T
  signal access_T_num_cont :  std_logic_vector(15 downto 0);
  signal access_T_row1 :  std_logic_vector(15 downto 0);
  signal access_T_col1 :  std_logic_vector(15 downto 0);
  signal access_T_rk1 :  std_logic_vector(15 downto 0);
  signal access_T_chl_in :  std_logic_vector(15 downto 0);
  signal access_T_ct :  std_logic_vector(15 downto 0);
  signal access_T_in_args    : std_logic_vector(95 downto 0);
  signal access_T_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal access_T_tag_out   : std_logic_vector(1 downto 0);
  signal access_T_start_req : std_logic;
  signal access_T_start_ack : std_logic;
  signal access_T_fin_req   : std_logic;
  signal access_T_fin_ack : std_logic;
  -- caller side aggregated signals for module access_T
  signal access_T_call_reqs: std_logic_vector(0 downto 0);
  signal access_T_call_acks: std_logic_vector(0 downto 0);
  signal access_T_return_reqs: std_logic_vector(0 downto 0);
  signal access_T_return_acks: std_logic_vector(0 downto 0);
  signal access_T_call_data: std_logic_vector(95 downto 0);
  signal access_T_call_tag: std_logic_vector(0 downto 0);
  signal access_T_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module convolution3D
  component convolution3D is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(1 downto 0);
      maxpool_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      maxpool_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      maxpool_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      elapsed_time_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      elapsed_time_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      elapsed_time_pipe_pipe_write_data : out  std_logic_vector(63 downto 0);
      maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      num_out_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      num_out_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      num_out_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
      access_T_call_reqs : out  std_logic_vector(0 downto 0);
      access_T_call_acks : in   std_logic_vector(0 downto 0);
      access_T_call_data : out  std_logic_vector(95 downto 0);
      access_T_call_tag  :  out  std_logic_vector(0 downto 0);
      access_T_return_reqs : out  std_logic_vector(0 downto 0);
      access_T_return_acks : in   std_logic_vector(0 downto 0);
      access_T_return_tag :  in   std_logic_vector(0 downto 0);
      timer_call_reqs : out  std_logic_vector(0 downto 0);
      timer_call_acks : in   std_logic_vector(0 downto 0);
      timer_call_tag  :  out  std_logic_vector(1 downto 0);
      timer_return_reqs : out  std_logic_vector(0 downto 0);
      timer_return_acks : in   std_logic_vector(0 downto 0);
      timer_return_data : in   std_logic_vector(63 downto 0);
      timer_return_tag :  in   std_logic_vector(1 downto 0);
      loadKernelChannel_call_reqs : out  std_logic_vector(0 downto 0);
      loadKernelChannel_call_acks : in   std_logic_vector(0 downto 0);
      loadKernelChannel_call_data : out  std_logic_vector(127 downto 0);
      loadKernelChannel_call_tag  :  out  std_logic_vector(0 downto 0);
      loadKernelChannel_return_reqs : out  std_logic_vector(0 downto 0);
      loadKernelChannel_return_acks : in   std_logic_vector(0 downto 0);
      loadKernelChannel_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convolution3D
  signal convolution3D_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convolution3D_tag_out   : std_logic_vector(1 downto 0);
  signal convolution3D_start_req : std_logic;
  signal convolution3D_start_ack : std_logic;
  signal convolution3D_fin_req   : std_logic;
  signal convolution3D_fin_ack : std_logic;
  -- declarations related to module convolve
  component convolve is -- 
    generic (tag_length : integer); 
    port ( -- 
      input_pipe1_pipe_read_req : out  std_logic_vector(0 downto 0);
      input_pipe1_pipe_read_ack : in   std_logic_vector(0 downto 0);
      input_pipe1_pipe_read_data : in   std_logic_vector(15 downto 0);
      num_out_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      num_out_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      num_out_pipe_pipe_read_data : in   std_logic_vector(15 downto 0);
      size_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      size_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      size_pipe_pipe_read_data : in   std_logic_vector(31 downto 0);
      kernel_pipe1_pipe_read_req : out  std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_read_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_read_data : in   std_logic_vector(15 downto 0);
      input_done_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_done_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_done_pipe_pipe_write_data : out  std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      kernel_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convolve
  signal convolve_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convolve_tag_out   : std_logic_vector(1 downto 0);
  signal convolve_start_req : std_logic;
  signal convolve_start_ack : std_logic;
  signal convolve_fin_req   : std_logic;
  signal convolve_fin_ack : std_logic;
  -- declarations related to module loadKernelChannel
  component loadKernelChannel is -- 
    generic (tag_length : integer); 
    port ( -- 
      start_add : in  std_logic_vector(63 downto 0);
      end_add : in  std_logic_vector(63 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
      input_done_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_data : in   std_logic_vector(0 downto 0);
      size_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      size_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      size_pipe_pipe_write_data : out  std_logic_vector(31 downto 0);
      kernel_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module loadKernelChannel
  signal loadKernelChannel_start_add :  std_logic_vector(63 downto 0);
  signal loadKernelChannel_end_add :  std_logic_vector(63 downto 0);
  signal loadKernelChannel_in_args    : std_logic_vector(127 downto 0);
  signal loadKernelChannel_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal loadKernelChannel_tag_out   : std_logic_vector(1 downto 0);
  signal loadKernelChannel_start_req : std_logic;
  signal loadKernelChannel_start_ack : std_logic;
  signal loadKernelChannel_fin_req   : std_logic;
  signal loadKernelChannel_fin_ack : std_logic;
  -- caller side aggregated signals for module loadKernelChannel
  signal loadKernelChannel_call_reqs: std_logic_vector(0 downto 0);
  signal loadKernelChannel_call_acks: std_logic_vector(0 downto 0);
  signal loadKernelChannel_return_reqs: std_logic_vector(0 downto 0);
  signal loadKernelChannel_return_acks: std_logic_vector(0 downto 0);
  signal loadKernelChannel_call_data: std_logic_vector(127 downto 0);
  signal loadKernelChannel_call_tag: std_logic_vector(0 downto 0);
  signal loadKernelChannel_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module timer
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      c : out  std_logic_vector(63 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timer
  signal timer_c :  std_logic_vector(63 downto 0);
  signal timer_out_args   : std_logic_vector(63 downto 0);
  signal timer_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal timer_tag_out   : std_logic_vector(2 downto 0);
  signal timer_start_req : std_logic;
  signal timer_start_ack : std_logic;
  signal timer_fin_req   : std_logic;
  signal timer_fin_ack : std_logic;
  -- caller side aggregated signals for module timer
  signal timer_call_reqs: std_logic_vector(0 downto 0);
  signal timer_call_acks: std_logic_vector(0 downto 0);
  signal timer_return_reqs: std_logic_vector(0 downto 0);
  signal timer_return_acks: std_logic_vector(0 downto 0);
  signal timer_call_tag: std_logic_vector(1 downto 0);
  signal timer_return_data: std_logic_vector(63 downto 0);
  signal timer_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module timerDaemon
  component timerDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timerDaemon
  signal timerDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal timerDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal timerDaemon_start_req : std_logic;
  signal timerDaemon_start_ack : std_logic;
  signal timerDaemon_fin_req   : std_logic;
  signal timerDaemon_fin_ack : std_logic;
  -- aggregate signals for write to pipe elapsed_time_pipe
  signal elapsed_time_pipe_pipe_write_data: std_logic_vector(63 downto 0);
  signal elapsed_time_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal elapsed_time_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe input_done_pipe
  signal input_done_pipe_pipe_write_data: std_logic_vector(0 downto 0);
  signal input_done_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal input_done_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe input_done_pipe
  signal input_done_pipe_pipe_read_data: std_logic_vector(0 downto 0);
  signal input_done_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal input_done_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe input_pipe1
  signal input_pipe1_pipe_write_data: std_logic_vector(15 downto 0);
  signal input_pipe1_pipe_write_req: std_logic_vector(0 downto 0);
  signal input_pipe1_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe input_pipe1
  signal input_pipe1_pipe_read_data: std_logic_vector(15 downto 0);
  signal input_pipe1_pipe_read_req: std_logic_vector(0 downto 0);
  signal input_pipe1_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe kernel_pipe1
  signal kernel_pipe1_pipe_write_data: std_logic_vector(31 downto 0);
  signal kernel_pipe1_pipe_write_req: std_logic_vector(1 downto 0);
  signal kernel_pipe1_pipe_write_ack: std_logic_vector(1 downto 0);
  -- aggregate signals for read from pipe kernel_pipe1
  signal kernel_pipe1_pipe_read_data: std_logic_vector(15 downto 0);
  signal kernel_pipe1_pipe_read_req: std_logic_vector(0 downto 0);
  signal kernel_pipe1_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe maxpool_input_pipe
  signal maxpool_input_pipe_pipe_read_data: std_logic_vector(7 downto 0);
  signal maxpool_input_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal maxpool_input_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe maxpool_output_pipe
  signal maxpool_output_pipe_pipe_write_data: std_logic_vector(15 downto 0);
  signal maxpool_output_pipe_pipe_write_req: std_logic_vector(1 downto 0);
  signal maxpool_output_pipe_pipe_write_ack: std_logic_vector(1 downto 0);
  -- aggregate signals for write to pipe num_out_pipe
  signal num_out_pipe_pipe_write_data: std_logic_vector(15 downto 0);
  signal num_out_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal num_out_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe num_out_pipe
  signal num_out_pipe_pipe_read_data: std_logic_vector(15 downto 0);
  signal num_out_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal num_out_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe size_pipe
  signal size_pipe_pipe_write_data: std_logic_vector(31 downto 0);
  signal size_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal size_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe size_pipe
  signal size_pipe_pipe_read_data: std_logic_vector(31 downto 0);
  signal size_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal size_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module access_T
  access_T_num_cont <= access_T_in_args(95 downto 80);
  access_T_row1 <= access_T_in_args(79 downto 64);
  access_T_col1 <= access_T_in_args(63 downto 48);
  access_T_rk1 <= access_T_in_args(47 downto 32);
  access_T_chl_in <= access_T_in_args(31 downto 16);
  access_T_ct <= access_T_in_args(15 downto 0);
  -- call arbiter for module access_T
  access_T_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 96,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => access_T_call_reqs,
      call_acks => access_T_call_acks,
      return_reqs => access_T_return_reqs,
      return_acks => access_T_return_acks,
      call_data  => access_T_call_data,
      call_tag  => access_T_call_tag,
      return_tag  => access_T_return_tag,
      call_mtag => access_T_tag_in,
      return_mtag => access_T_tag_out,
      call_mreq => access_T_start_req,
      call_mack => access_T_start_ack,
      return_mreq => access_T_fin_req,
      return_mack => access_T_fin_ack,
      call_mdata => access_T_in_args,
      clk => clk, 
      reset => reset --
    ); --
  access_T_instance:access_T-- 
    generic map(tag_length => 2)
    port map(-- 
      num_cont => access_T_num_cont,
      row1 => access_T_row1,
      col1 => access_T_col1,
      rk1 => access_T_rk1,
      chl_in => access_T_chl_in,
      ct => access_T_ct,
      start_req => access_T_start_req,
      start_ack => access_T_start_ack,
      fin_req => access_T_fin_req,
      fin_ack => access_T_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(13 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(18 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(63 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(1 downto 0),
      input_pipe1_pipe_write_req => input_pipe1_pipe_write_req(0 downto 0),
      input_pipe1_pipe_write_ack => input_pipe1_pipe_write_ack(0 downto 0),
      input_pipe1_pipe_write_data => input_pipe1_pipe_write_data(15 downto 0),
      tag_in => access_T_tag_in,
      tag_out => access_T_tag_out-- 
    ); -- 
  -- module convolution3D
  convolution3D_instance:convolution3D-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convolution3D_start_req,
      start_ack => convolution3D_start_ack,
      fin_req => convolution3D_fin_req,
      fin_ack => convolution3D_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(13 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(63 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(18 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(1 downto 0),
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(13 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(63 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(18 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(1 downto 0),
      maxpool_input_pipe_pipe_read_req => maxpool_input_pipe_pipe_read_req(0 downto 0),
      maxpool_input_pipe_pipe_read_ack => maxpool_input_pipe_pipe_read_ack(0 downto 0),
      maxpool_input_pipe_pipe_read_data => maxpool_input_pipe_pipe_read_data(7 downto 0),
      elapsed_time_pipe_pipe_write_req => elapsed_time_pipe_pipe_write_req(0 downto 0),
      elapsed_time_pipe_pipe_write_ack => elapsed_time_pipe_pipe_write_ack(0 downto 0),
      elapsed_time_pipe_pipe_write_data => elapsed_time_pipe_pipe_write_data(63 downto 0),
      maxpool_output_pipe_pipe_write_req => maxpool_output_pipe_pipe_write_req(1 downto 1),
      maxpool_output_pipe_pipe_write_ack => maxpool_output_pipe_pipe_write_ack(1 downto 1),
      maxpool_output_pipe_pipe_write_data => maxpool_output_pipe_pipe_write_data(15 downto 8),
      num_out_pipe_pipe_write_req => num_out_pipe_pipe_write_req(0 downto 0),
      num_out_pipe_pipe_write_ack => num_out_pipe_pipe_write_ack(0 downto 0),
      num_out_pipe_pipe_write_data => num_out_pipe_pipe_write_data(15 downto 0),
      access_T_call_reqs => access_T_call_reqs(0 downto 0),
      access_T_call_acks => access_T_call_acks(0 downto 0),
      access_T_call_data => access_T_call_data(95 downto 0),
      access_T_call_tag => access_T_call_tag(0 downto 0),
      access_T_return_reqs => access_T_return_reqs(0 downto 0),
      access_T_return_acks => access_T_return_acks(0 downto 0),
      access_T_return_tag => access_T_return_tag(0 downto 0),
      timer_call_reqs => timer_call_reqs(0 downto 0),
      timer_call_acks => timer_call_acks(0 downto 0),
      timer_call_tag => timer_call_tag(1 downto 0),
      timer_return_reqs => timer_return_reqs(0 downto 0),
      timer_return_acks => timer_return_acks(0 downto 0),
      timer_return_data => timer_return_data(63 downto 0),
      timer_return_tag => timer_return_tag(1 downto 0),
      loadKernelChannel_call_reqs => loadKernelChannel_call_reqs(0 downto 0),
      loadKernelChannel_call_acks => loadKernelChannel_call_acks(0 downto 0),
      loadKernelChannel_call_data => loadKernelChannel_call_data(127 downto 0),
      loadKernelChannel_call_tag => loadKernelChannel_call_tag(0 downto 0),
      loadKernelChannel_return_reqs => loadKernelChannel_return_reqs(0 downto 0),
      loadKernelChannel_return_acks => loadKernelChannel_return_acks(0 downto 0),
      loadKernelChannel_return_tag => loadKernelChannel_return_tag(0 downto 0),
      tag_in => convolution3D_tag_in,
      tag_out => convolution3D_tag_out-- 
    ); -- 
  -- module will be run forever 
  convolution3D_tag_in <= (others => '0');
  convolution3D_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convolution3D_start_req, start_ack => convolution3D_start_ack,  fin_req => convolution3D_fin_req,  fin_ack => convolution3D_fin_ack);
  -- module convolve
  convolve_instance:convolve-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convolve_start_req,
      start_ack => convolve_start_ack,
      fin_req => convolve_fin_req,
      fin_ack => convolve_fin_ack,
      clk => clk,
      reset => reset,
      input_pipe1_pipe_read_req => input_pipe1_pipe_read_req(0 downto 0),
      input_pipe1_pipe_read_ack => input_pipe1_pipe_read_ack(0 downto 0),
      input_pipe1_pipe_read_data => input_pipe1_pipe_read_data(15 downto 0),
      num_out_pipe_pipe_read_req => num_out_pipe_pipe_read_req(0 downto 0),
      num_out_pipe_pipe_read_ack => num_out_pipe_pipe_read_ack(0 downto 0),
      num_out_pipe_pipe_read_data => num_out_pipe_pipe_read_data(15 downto 0),
      size_pipe_pipe_read_req => size_pipe_pipe_read_req(0 downto 0),
      size_pipe_pipe_read_ack => size_pipe_pipe_read_ack(0 downto 0),
      size_pipe_pipe_read_data => size_pipe_pipe_read_data(31 downto 0),
      kernel_pipe1_pipe_read_req => kernel_pipe1_pipe_read_req(0 downto 0),
      kernel_pipe1_pipe_read_ack => kernel_pipe1_pipe_read_ack(0 downto 0),
      kernel_pipe1_pipe_read_data => kernel_pipe1_pipe_read_data(15 downto 0),
      input_done_pipe_pipe_write_req => input_done_pipe_pipe_write_req(0 downto 0),
      input_done_pipe_pipe_write_ack => input_done_pipe_pipe_write_ack(0 downto 0),
      input_done_pipe_pipe_write_data => input_done_pipe_pipe_write_data(0 downto 0),
      maxpool_output_pipe_pipe_write_req => maxpool_output_pipe_pipe_write_req(0 downto 0),
      maxpool_output_pipe_pipe_write_ack => maxpool_output_pipe_pipe_write_ack(0 downto 0),
      maxpool_output_pipe_pipe_write_data => maxpool_output_pipe_pipe_write_data(7 downto 0),
      kernel_pipe1_pipe_write_req => kernel_pipe1_pipe_write_req(0 downto 0),
      kernel_pipe1_pipe_write_ack => kernel_pipe1_pipe_write_ack(0 downto 0),
      kernel_pipe1_pipe_write_data => kernel_pipe1_pipe_write_data(15 downto 0),
      tag_in => convolve_tag_in,
      tag_out => convolve_tag_out-- 
    ); -- 
  -- module will be run forever 
  convolve_tag_in <= (others => '0');
  convolve_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convolve_start_req, start_ack => convolve_start_ack,  fin_req => convolve_fin_req,  fin_ack => convolve_fin_ack);
  -- module loadKernelChannel
  loadKernelChannel_start_add <= loadKernelChannel_in_args(127 downto 64);
  loadKernelChannel_end_add <= loadKernelChannel_in_args(63 downto 0);
  -- call arbiter for module loadKernelChannel
  loadKernelChannel_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 128,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => loadKernelChannel_call_reqs,
      call_acks => loadKernelChannel_call_acks,
      return_reqs => loadKernelChannel_return_reqs,
      return_acks => loadKernelChannel_return_acks,
      call_data  => loadKernelChannel_call_data,
      call_tag  => loadKernelChannel_call_tag,
      return_tag  => loadKernelChannel_return_tag,
      call_mtag => loadKernelChannel_tag_in,
      return_mtag => loadKernelChannel_tag_out,
      call_mreq => loadKernelChannel_start_req,
      call_mack => loadKernelChannel_start_ack,
      return_mreq => loadKernelChannel_fin_req,
      return_mack => loadKernelChannel_fin_ack,
      call_mdata => loadKernelChannel_in_args,
      clk => clk, 
      reset => reset --
    ); --
  loadKernelChannel_instance:loadKernelChannel-- 
    generic map(tag_length => 2)
    port map(-- 
      start_add => loadKernelChannel_start_add,
      end_add => loadKernelChannel_end_add,
      start_req => loadKernelChannel_start_req,
      start_ack => loadKernelChannel_start_ack,
      fin_req => loadKernelChannel_fin_req,
      fin_ack => loadKernelChannel_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(13 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(18 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(1 downto 0),
      input_done_pipe_pipe_read_req => input_done_pipe_pipe_read_req(0 downto 0),
      input_done_pipe_pipe_read_ack => input_done_pipe_pipe_read_ack(0 downto 0),
      input_done_pipe_pipe_read_data => input_done_pipe_pipe_read_data(0 downto 0),
      size_pipe_pipe_write_req => size_pipe_pipe_write_req(0 downto 0),
      size_pipe_pipe_write_ack => size_pipe_pipe_write_ack(0 downto 0),
      size_pipe_pipe_write_data => size_pipe_pipe_write_data(31 downto 0),
      kernel_pipe1_pipe_write_req => kernel_pipe1_pipe_write_req(1 downto 1),
      kernel_pipe1_pipe_write_ack => kernel_pipe1_pipe_write_ack(1 downto 1),
      kernel_pipe1_pipe_write_data => kernel_pipe1_pipe_write_data(31 downto 16),
      tag_in => loadKernelChannel_tag_in,
      tag_out => loadKernelChannel_tag_out-- 
    ); -- 
  -- module timer
  timer_out_args <= timer_c ;
  -- call arbiter for module timer
  timer_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargs", num_reqs => 1,
      return_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => timer_call_reqs,
      call_acks => timer_call_acks,
      return_reqs => timer_return_reqs,
      return_acks => timer_return_acks,
      call_tag  => timer_call_tag,
      return_tag  => timer_return_tag,
      call_mtag => timer_tag_in,
      return_mtag => timer_tag_out,
      return_data =>timer_return_data,
      call_mreq => timer_start_req,
      call_mack => timer_start_ack,
      return_mreq => timer_fin_req,
      return_mack => timer_fin_ack,
      return_mdata => timer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  timer_instance:timer-- 
    generic map(tag_length => 3)
    port map(-- 
      c => timer_c,
      start_req => timer_start_req,
      start_ack => timer_start_ack,
      fin_req => timer_fin_req,
      fin_ack => timer_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_2_lr_req => memory_space_2_lr_req(0 downto 0),
      memory_space_2_lr_ack => memory_space_2_lr_ack(0 downto 0),
      memory_space_2_lr_addr => memory_space_2_lr_addr(0 downto 0),
      memory_space_2_lr_tag => memory_space_2_lr_tag(17 downto 0),
      memory_space_2_lc_req => memory_space_2_lc_req(0 downto 0),
      memory_space_2_lc_ack => memory_space_2_lc_ack(0 downto 0),
      memory_space_2_lc_data => memory_space_2_lc_data(63 downto 0),
      memory_space_2_lc_tag => memory_space_2_lc_tag(0 downto 0),
      tag_in => timer_tag_in,
      tag_out => timer_tag_out-- 
    ); -- 
  -- module timerDaemon
  timerDaemon_instance:timerDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => timerDaemon_start_req,
      start_ack => timerDaemon_start_ack,
      fin_req => timerDaemon_fin_req,
      fin_ack => timerDaemon_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_2_sr_req => memory_space_2_sr_req(0 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(0 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(0 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(63 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(17 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(0 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(0 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(0 downto 0),
      tag_in => timerDaemon_tag_in,
      tag_out => timerDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  timerDaemon_tag_in <= (others => '0');
  timerDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => timerDaemon_start_req, start_ack => timerDaemon_start_ack,  fin_req => timerDaemon_fin_req,  fin_ack => timerDaemon_fin_ack);
  elapsed_time_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe elapsed_time_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => elapsed_time_pipe_pipe_read_req,
      read_ack => elapsed_time_pipe_pipe_read_ack,
      read_data => elapsed_time_pipe_pipe_read_data,
      write_req => elapsed_time_pipe_pipe_write_req,
      write_ack => elapsed_time_pipe_pipe_write_ack,
      write_data => elapsed_time_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  input_done_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe input_done_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 1,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => input_done_pipe_pipe_read_req,
      read_ack => input_done_pipe_pipe_read_ack,
      read_data => input_done_pipe_pipe_read_data,
      write_req => input_done_pipe_pipe_write_req,
      write_ack => input_done_pipe_pipe_write_ack,
      write_data => input_done_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  input_pipe1_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe input_pipe1",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 100 --
    )
    port map( -- 
      read_req => input_pipe1_pipe_read_req,
      read_ack => input_pipe1_pipe_read_ack,
      read_data => input_pipe1_pipe_read_data,
      write_req => input_pipe1_pipe_write_req,
      write_ack => input_pipe1_pipe_write_ack,
      write_data => input_pipe1_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  kernel_pipe1_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe kernel_pipe1",
      num_reads => 1,
      num_writes => 2,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 100 --
    )
    port map( -- 
      read_req => kernel_pipe1_pipe_read_req,
      read_ack => kernel_pipe1_pipe_read_ack,
      read_data => kernel_pipe1_pipe_read_data,
      write_req => kernel_pipe1_pipe_write_req,
      write_ack => kernel_pipe1_pipe_write_ack,
      write_data => kernel_pipe1_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  maxpool_input_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe maxpool_input_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => maxpool_input_pipe_pipe_read_req,
      read_ack => maxpool_input_pipe_pipe_read_ack,
      read_data => maxpool_input_pipe_pipe_read_data,
      write_req => maxpool_input_pipe_pipe_write_req,
      write_ack => maxpool_input_pipe_pipe_write_ack,
      write_data => maxpool_input_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  maxpool_output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe maxpool_output_pipe",
      num_reads => 1,
      num_writes => 2,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => maxpool_output_pipe_pipe_read_req,
      read_ack => maxpool_output_pipe_pipe_read_ack,
      read_data => maxpool_output_pipe_pipe_read_data,
      write_req => maxpool_output_pipe_pipe_write_req,
      write_ack => maxpool_output_pipe_pipe_write_ack,
      write_data => maxpool_output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  num_out_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe num_out_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => num_out_pipe_pipe_read_req,
      read_ack => num_out_pipe_pipe_read_ack,
      read_data => num_out_pipe_pipe_read_data,
      write_req => num_out_pipe_pipe_write_req,
      write_ack => num_out_pipe_pipe_write_ack,
      write_data => num_out_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  size_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe size_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => size_pipe_pipe_read_req,
      read_ack => size_pipe_pipe_read_ack,
      read_data => size_pipe_pipe_read_data,
      write_req => size_pipe_pipe_write_req,
      write_ack => size_pipe_pipe_write_ack,
      write_data => size_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  MemorySpace_memory_space_0: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 2,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_1: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 2,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_2: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_2",
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_2_lr_addr,
      lr_req_in => memory_space_2_lr_req,
      lr_ack_out => memory_space_2_lr_ack,
      lr_tag_in => memory_space_2_lr_tag,
      lc_req_in => memory_space_2_lc_req,
      lc_ack_out => memory_space_2_lc_ack,
      lc_data_out => memory_space_2_lc_data,
      lc_tag_out => memory_space_2_lc_tag,
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
