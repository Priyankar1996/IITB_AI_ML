-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity sendOutput is -- 
  generic (tag_length : integer); 
  port ( -- 
    size : in  std_logic_vector(31 downto 0);
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
    zeropad_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    zeropad_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    zeropad_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity sendOutput;
architecture sendOutput_arch of sendOutput is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 32)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal size_buffer :  std_logic_vector(31 downto 0);
  signal size_update_enable: Boolean;
  -- output port buffer signals
  signal sendOutput_CP_26_start: Boolean;
  signal sendOutput_CP_26_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal if_stmt_44_branch_req_0 : boolean;
  signal if_stmt_44_branch_ack_1 : boolean;
  signal if_stmt_44_branch_ack_0 : boolean;
  signal type_cast_53_inst_req_0 : boolean;
  signal type_cast_53_inst_ack_0 : boolean;
  signal type_cast_53_inst_req_1 : boolean;
  signal type_cast_53_inst_ack_1 : boolean;
  signal array_obj_ref_69_index_offset_req_0 : boolean;
  signal array_obj_ref_69_index_offset_ack_0 : boolean;
  signal array_obj_ref_69_index_offset_req_1 : boolean;
  signal array_obj_ref_69_index_offset_ack_1 : boolean;
  signal addr_of_70_final_reg_req_0 : boolean;
  signal addr_of_70_final_reg_ack_0 : boolean;
  signal addr_of_70_final_reg_req_1 : boolean;
  signal addr_of_70_final_reg_ack_1 : boolean;
  signal ptr_deref_74_load_0_req_0 : boolean;
  signal ptr_deref_74_load_0_ack_0 : boolean;
  signal ptr_deref_74_load_0_req_1 : boolean;
  signal ptr_deref_74_load_0_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_165_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_165_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_168_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_168_inst_ack_0 : boolean;
  signal type_cast_78_inst_req_0 : boolean;
  signal type_cast_78_inst_ack_0 : boolean;
  signal type_cast_78_inst_req_1 : boolean;
  signal type_cast_78_inst_ack_1 : boolean;
  signal type_cast_88_inst_req_0 : boolean;
  signal type_cast_88_inst_ack_0 : boolean;
  signal type_cast_88_inst_req_1 : boolean;
  signal type_cast_88_inst_ack_1 : boolean;
  signal type_cast_98_inst_req_0 : boolean;
  signal type_cast_98_inst_ack_0 : boolean;
  signal type_cast_98_inst_req_1 : boolean;
  signal type_cast_98_inst_ack_1 : boolean;
  signal type_cast_108_inst_req_0 : boolean;
  signal type_cast_108_inst_ack_0 : boolean;
  signal type_cast_108_inst_req_1 : boolean;
  signal type_cast_108_inst_ack_1 : boolean;
  signal type_cast_118_inst_req_0 : boolean;
  signal type_cast_118_inst_ack_0 : boolean;
  signal type_cast_118_inst_req_1 : boolean;
  signal type_cast_118_inst_ack_1 : boolean;
  signal type_cast_128_inst_req_0 : boolean;
  signal type_cast_128_inst_ack_0 : boolean;
  signal type_cast_128_inst_req_1 : boolean;
  signal type_cast_128_inst_ack_1 : boolean;
  signal type_cast_138_inst_req_0 : boolean;
  signal type_cast_138_inst_ack_0 : boolean;
  signal type_cast_138_inst_req_1 : boolean;
  signal type_cast_138_inst_ack_1 : boolean;
  signal type_cast_148_inst_req_0 : boolean;
  signal type_cast_148_inst_ack_0 : boolean;
  signal type_cast_148_inst_req_1 : boolean;
  signal type_cast_148_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_150_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_150_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_150_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_150_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_153_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_153_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_153_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_153_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_156_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_156_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_156_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_156_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_159_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_159_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_159_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_159_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_162_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_162_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_162_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_162_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_165_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_165_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_168_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_168_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_171_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_171_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_171_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_171_inst_ack_1 : boolean;
  signal if_stmt_185_branch_req_0 : boolean;
  signal if_stmt_185_branch_ack_1 : boolean;
  signal if_stmt_185_branch_ack_0 : boolean;
  signal phi_stmt_57_req_0 : boolean;
  signal type_cast_63_inst_req_0 : boolean;
  signal type_cast_63_inst_ack_0 : boolean;
  signal type_cast_63_inst_req_1 : boolean;
  signal type_cast_63_inst_ack_1 : boolean;
  signal phi_stmt_57_req_1 : boolean;
  signal phi_stmt_57_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "sendOutput_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 32) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(31 downto 0) <= size;
  size_buffer <= in_buffer_data_out(31 downto 0);
  in_buffer_data_in(tag_length + 31 downto 32) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 31 downto 32);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  sendOutput_CP_26_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "sendOutput_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendOutput_CP_26_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= sendOutput_CP_26_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendOutput_CP_26_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  sendOutput_CP_26: Block -- control-path 
    signal sendOutput_CP_26_elements: BooleanArray(59 downto 0);
    -- 
  begin -- 
    sendOutput_CP_26_elements(0) <= sendOutput_CP_26_start;
    sendOutput_CP_26_symbol <= sendOutput_CP_26_elements(59);
    -- CP-element group 0:  branch  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (15) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_24/$entry
      -- CP-element group 0: 	 branch_block_stmt_24/branch_block_stmt_24__entry__
      -- CP-element group 0: 	 branch_block_stmt_24/assign_stmt_34_to_assign_stmt_43__entry__
      -- CP-element group 0: 	 branch_block_stmt_24/assign_stmt_34_to_assign_stmt_43__exit__
      -- CP-element group 0: 	 branch_block_stmt_24/if_stmt_44__entry__
      -- CP-element group 0: 	 branch_block_stmt_24/assign_stmt_34_to_assign_stmt_43/$entry
      -- CP-element group 0: 	 branch_block_stmt_24/assign_stmt_34_to_assign_stmt_43/$exit
      -- CP-element group 0: 	 branch_block_stmt_24/if_stmt_44_dead_link/$entry
      -- CP-element group 0: 	 branch_block_stmt_24/if_stmt_44_eval_test/$entry
      -- CP-element group 0: 	 branch_block_stmt_24/if_stmt_44_eval_test/$exit
      -- CP-element group 0: 	 branch_block_stmt_24/if_stmt_44_eval_test/branch_req
      -- CP-element group 0: 	 branch_block_stmt_24/R_cmp68_45_place
      -- CP-element group 0: 	 branch_block_stmt_24/if_stmt_44_if_link/$entry
      -- CP-element group 0: 	 branch_block_stmt_24/if_stmt_44_else_link/$entry
      -- 
    branch_req_64_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_64_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(0), ack => if_stmt_44_branch_req_0); -- 
    -- CP-element group 1:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	3 
    -- CP-element group 1: 	4 
    -- CP-element group 1:  members (18) 
      -- CP-element group 1: 	 branch_block_stmt_24/entry_bbx_xnph
      -- CP-element group 1: 	 branch_block_stmt_24/merge_stmt_50__exit__
      -- CP-element group 1: 	 branch_block_stmt_24/assign_stmt_54__entry__
      -- CP-element group 1: 	 branch_block_stmt_24/if_stmt_44_if_link/$exit
      -- CP-element group 1: 	 branch_block_stmt_24/if_stmt_44_if_link/if_choice_transition
      -- CP-element group 1: 	 branch_block_stmt_24/assign_stmt_54/$entry
      -- CP-element group 1: 	 branch_block_stmt_24/assign_stmt_54/type_cast_53_sample_start_
      -- CP-element group 1: 	 branch_block_stmt_24/assign_stmt_54/type_cast_53_update_start_
      -- CP-element group 1: 	 branch_block_stmt_24/assign_stmt_54/type_cast_53_Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_24/assign_stmt_54/type_cast_53_Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_24/assign_stmt_54/type_cast_53_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_24/assign_stmt_54/type_cast_53_Update/cr
      -- CP-element group 1: 	 branch_block_stmt_24/entry_bbx_xnph_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_24/entry_bbx_xnph_PhiReq/$exit
      -- CP-element group 1: 	 branch_block_stmt_24/merge_stmt_50_PhiReqMerge
      -- CP-element group 1: 	 branch_block_stmt_24/merge_stmt_50_PhiAck/$entry
      -- CP-element group 1: 	 branch_block_stmt_24/merge_stmt_50_PhiAck/$exit
      -- CP-element group 1: 	 branch_block_stmt_24/merge_stmt_50_PhiAck/dummy
      -- 
    if_choice_transition_69_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_44_branch_ack_1, ack => sendOutput_CP_26_elements(1)); -- 
    rr_86_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_86_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(1), ack => type_cast_53_inst_req_0); -- 
    cr_91_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_91_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(1), ack => type_cast_53_inst_req_1); -- 
    -- CP-element group 2:  transition  place  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	59 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 branch_block_stmt_24/entry_forx_xend
      -- CP-element group 2: 	 branch_block_stmt_24/if_stmt_44_else_link/$exit
      -- CP-element group 2: 	 branch_block_stmt_24/if_stmt_44_else_link/else_choice_transition
      -- CP-element group 2: 	 branch_block_stmt_24/entry_forx_xend_PhiReq/$entry
      -- CP-element group 2: 	 branch_block_stmt_24/entry_forx_xend_PhiReq/$exit
      -- 
    else_choice_transition_73_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_44_branch_ack_0, ack => sendOutput_CP_26_elements(2)); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	1 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_24/assign_stmt_54/type_cast_53_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_24/assign_stmt_54/type_cast_53_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_24/assign_stmt_54/type_cast_53_Sample/ra
      -- 
    ra_87_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_53_inst_ack_0, ack => sendOutput_CP_26_elements(3)); -- 
    -- CP-element group 4:  transition  place  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	1 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	53 
    -- CP-element group 4:  members (9) 
      -- CP-element group 4: 	 branch_block_stmt_24/assign_stmt_54__exit__
      -- CP-element group 4: 	 branch_block_stmt_24/bbx_xnph_forx_xbody
      -- CP-element group 4: 	 branch_block_stmt_24/assign_stmt_54/$exit
      -- CP-element group 4: 	 branch_block_stmt_24/assign_stmt_54/type_cast_53_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_24/assign_stmt_54/type_cast_53_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_24/assign_stmt_54/type_cast_53_Update/ca
      -- CP-element group 4: 	 branch_block_stmt_24/bbx_xnph_forx_xbody_PhiReq/$entry
      -- CP-element group 4: 	 branch_block_stmt_24/bbx_xnph_forx_xbody_PhiReq/phi_stmt_57/$entry
      -- CP-element group 4: 	 branch_block_stmt_24/bbx_xnph_forx_xbody_PhiReq/phi_stmt_57/phi_stmt_57_sources/$entry
      -- 
    ca_92_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_53_inst_ack_1, ack => sendOutput_CP_26_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	58 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	50 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/array_obj_ref_69_final_index_sum_regn_sample_complete
      -- CP-element group 5: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/array_obj_ref_69_final_index_sum_regn_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/array_obj_ref_69_final_index_sum_regn_Sample/ack
      -- 
    ack_121_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_69_index_offset_ack_0, ack => sendOutput_CP_26_elements(5)); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	58 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (11) 
      -- CP-element group 6: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/addr_of_70_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/array_obj_ref_69_root_address_calculated
      -- CP-element group 6: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/array_obj_ref_69_offset_calculated
      -- CP-element group 6: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/array_obj_ref_69_final_index_sum_regn_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/array_obj_ref_69_final_index_sum_regn_Update/ack
      -- CP-element group 6: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/array_obj_ref_69_base_plus_offset/$entry
      -- CP-element group 6: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/array_obj_ref_69_base_plus_offset/$exit
      -- CP-element group 6: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/array_obj_ref_69_base_plus_offset/sum_rename_req
      -- CP-element group 6: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/array_obj_ref_69_base_plus_offset/sum_rename_ack
      -- CP-element group 6: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/addr_of_70_request/$entry
      -- CP-element group 6: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/addr_of_70_request/req
      -- 
    ack_126_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_69_index_offset_ack_1, ack => sendOutput_CP_26_elements(6)); -- 
    req_135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(6), ack => addr_of_70_final_reg_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/addr_of_70_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/addr_of_70_request/$exit
      -- CP-element group 7: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/addr_of_70_request/ack
      -- 
    ack_136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_70_final_reg_ack_0, ack => sendOutput_CP_26_elements(7)); -- 
    -- CP-element group 8:  join  fork  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	58 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (24) 
      -- CP-element group 8: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/addr_of_70_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/addr_of_70_complete/$exit
      -- CP-element group 8: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/addr_of_70_complete/ack
      -- CP-element group 8: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/ptr_deref_74_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/ptr_deref_74_base_address_calculated
      -- CP-element group 8: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/ptr_deref_74_word_address_calculated
      -- CP-element group 8: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/ptr_deref_74_root_address_calculated
      -- CP-element group 8: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/ptr_deref_74_base_address_resized
      -- CP-element group 8: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/ptr_deref_74_base_addr_resize/$entry
      -- CP-element group 8: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/ptr_deref_74_base_addr_resize/$exit
      -- CP-element group 8: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/ptr_deref_74_base_addr_resize/base_resize_req
      -- CP-element group 8: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/ptr_deref_74_base_addr_resize/base_resize_ack
      -- CP-element group 8: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/ptr_deref_74_base_plus_offset/$entry
      -- CP-element group 8: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/ptr_deref_74_base_plus_offset/$exit
      -- CP-element group 8: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/ptr_deref_74_base_plus_offset/sum_rename_req
      -- CP-element group 8: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/ptr_deref_74_base_plus_offset/sum_rename_ack
      -- CP-element group 8: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/ptr_deref_74_word_addrgen/$entry
      -- CP-element group 8: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/ptr_deref_74_word_addrgen/$exit
      -- CP-element group 8: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/ptr_deref_74_word_addrgen/root_register_req
      -- CP-element group 8: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/ptr_deref_74_word_addrgen/root_register_ack
      -- CP-element group 8: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/ptr_deref_74_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/ptr_deref_74_Sample/word_access_start/$entry
      -- CP-element group 8: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/ptr_deref_74_Sample/word_access_start/word_0/$entry
      -- CP-element group 8: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/ptr_deref_74_Sample/word_access_start/word_0/rr
      -- 
    ack_141_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_70_final_reg_ack_1, ack => sendOutput_CP_26_elements(8)); -- 
    rr_174_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_174_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(8), ack => ptr_deref_74_load_0_req_0); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (5) 
      -- CP-element group 9: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/ptr_deref_74_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/ptr_deref_74_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/ptr_deref_74_Sample/word_access_start/$exit
      -- CP-element group 9: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/ptr_deref_74_Sample/word_access_start/word_0/$exit
      -- CP-element group 9: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/ptr_deref_74_Sample/word_access_start/word_0/ra
      -- 
    ra_175_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_74_load_0_ack_0, ack => sendOutput_CP_26_elements(9)); -- 
    -- CP-element group 10:  fork  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	58 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10: 	13 
    -- CP-element group 10: 	23 
    -- CP-element group 10: 	21 
    -- CP-element group 10: 	19 
    -- CP-element group 10: 	17 
    -- CP-element group 10: 	25 
    -- CP-element group 10: 	15 
    -- CP-element group 10:  members (33) 
      -- CP-element group 10: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_78_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/ptr_deref_74_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/ptr_deref_74_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/ptr_deref_74_Update/word_access_complete/$exit
      -- CP-element group 10: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/ptr_deref_74_Update/word_access_complete/word_0/$exit
      -- CP-element group 10: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/ptr_deref_74_Update/word_access_complete/word_0/ca
      -- CP-element group 10: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/ptr_deref_74_Update/ptr_deref_74_Merge/$entry
      -- CP-element group 10: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/ptr_deref_74_Update/ptr_deref_74_Merge/$exit
      -- CP-element group 10: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/ptr_deref_74_Update/ptr_deref_74_Merge/merge_req
      -- CP-element group 10: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/ptr_deref_74_Update/ptr_deref_74_Merge/merge_ack
      -- CP-element group 10: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_78_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_78_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_88_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_88_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_88_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_98_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_98_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_98_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_108_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_108_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_108_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_118_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_118_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_118_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_128_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_128_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_128_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_138_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_138_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_138_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_148_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_148_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_148_Sample/rr
      -- 
    ca_186_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_74_load_0_ack_1, ack => sendOutput_CP_26_elements(10)); -- 
    rr_213_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_213_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(10), ack => type_cast_88_inst_req_0); -- 
    rr_227_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_227_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(10), ack => type_cast_98_inst_req_0); -- 
    rr_199_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_199_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(10), ack => type_cast_78_inst_req_0); -- 
    rr_241_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_241_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(10), ack => type_cast_108_inst_req_0); -- 
    rr_283_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_283_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(10), ack => type_cast_138_inst_req_0); -- 
    rr_269_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_269_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(10), ack => type_cast_128_inst_req_0); -- 
    rr_255_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_255_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(10), ack => type_cast_118_inst_req_0); -- 
    rr_297_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_297_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(10), ack => type_cast_148_inst_req_0); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_78_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_78_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_78_Sample/ra
      -- 
    ra_200_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_78_inst_ack_0, ack => sendOutput_CP_26_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	58 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	47 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_78_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_78_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_78_Update/ca
      -- 
    ca_205_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_78_inst_ack_1, ack => sendOutput_CP_26_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	10 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_88_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_88_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_88_Sample/ra
      -- 
    ra_214_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_88_inst_ack_0, ack => sendOutput_CP_26_elements(13)); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	58 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	44 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_88_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_88_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_88_Update/ca
      -- 
    ca_219_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_88_inst_ack_1, ack => sendOutput_CP_26_elements(14)); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	10 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_98_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_98_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_98_Sample/ra
      -- 
    ra_228_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_98_inst_ack_0, ack => sendOutput_CP_26_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	58 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	41 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_98_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_98_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_98_Update/ca
      -- 
    ca_233_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_98_inst_ack_1, ack => sendOutput_CP_26_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	10 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_108_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_108_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_108_Sample/ra
      -- 
    ra_242_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_108_inst_ack_0, ack => sendOutput_CP_26_elements(17)); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	58 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	38 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_108_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_108_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_108_Update/ca
      -- 
    ca_247_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_108_inst_ack_1, ack => sendOutput_CP_26_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	10 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_118_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_118_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_118_Sample/ra
      -- 
    ra_256_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_118_inst_ack_0, ack => sendOutput_CP_26_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	58 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	35 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_118_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_118_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_118_Update/ca
      -- 
    ca_261_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_118_inst_ack_1, ack => sendOutput_CP_26_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	10 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_128_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_128_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_128_Sample/ra
      -- 
    ra_270_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_128_inst_ack_0, ack => sendOutput_CP_26_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	58 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	32 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_128_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_128_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_128_Update/ca
      -- 
    ca_275_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_128_inst_ack_1, ack => sendOutput_CP_26_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	10 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_138_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_138_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_138_Sample/ra
      -- 
    ra_284_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_138_inst_ack_0, ack => sendOutput_CP_26_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	58 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	29 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_138_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_138_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_138_Update/ca
      -- 
    ca_289_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_138_inst_ack_1, ack => sendOutput_CP_26_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	10 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_148_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_148_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_148_Sample/ra
      -- 
    ra_298_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_148_inst_ack_0, ack => sendOutput_CP_26_elements(25)); -- 
    -- CP-element group 26:  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	58 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (6) 
      -- CP-element group 26: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_148_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_148_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_148_Update/ca
      -- CP-element group 26: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_150_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_150_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_150_Sample/req
      -- 
    ca_303_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_148_inst_ack_1, ack => sendOutput_CP_26_elements(26)); -- 
    req_311_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_311_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(26), ack => WPIPE_zeropad_output_pipe_150_inst_req_0); -- 
    -- CP-element group 27:  transition  input  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27:  members (6) 
      -- CP-element group 27: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_150_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_150_update_start_
      -- CP-element group 27: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_150_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_150_Sample/ack
      -- CP-element group 27: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_150_Update/$entry
      -- CP-element group 27: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_150_Update/req
      -- 
    ack_312_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_150_inst_ack_0, ack => sendOutput_CP_26_elements(27)); -- 
    req_316_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_316_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(27), ack => WPIPE_zeropad_output_pipe_150_inst_req_1); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_150_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_150_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_150_Update/ack
      -- 
    ack_317_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_150_inst_ack_1, ack => sendOutput_CP_26_elements(28)); -- 
    -- CP-element group 29:  join  transition  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: 	24 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_153_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_153_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_153_Sample/req
      -- 
    req_325_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_325_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(29), ack => WPIPE_zeropad_output_pipe_153_inst_req_0); -- 
    sendOutput_cp_element_group_29: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_29"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(28) & sendOutput_CP_26_elements(24);
      gj_sendOutput_cp_element_group_29 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(29), clk => clk, reset => reset); --
    end block;
    -- CP-element group 30:  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (6) 
      -- CP-element group 30: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_153_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_153_update_start_
      -- CP-element group 30: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_153_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_153_Sample/ack
      -- CP-element group 30: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_153_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_153_Update/req
      -- 
    ack_326_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_153_inst_ack_0, ack => sendOutput_CP_26_elements(30)); -- 
    req_330_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_330_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(30), ack => WPIPE_zeropad_output_pipe_153_inst_req_1); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_153_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_153_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_153_Update/ack
      -- 
    ack_331_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_153_inst_ack_1, ack => sendOutput_CP_26_elements(31)); -- 
    -- CP-element group 32:  join  transition  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	22 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_156_sample_start_
      -- CP-element group 32: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_156_Sample/$entry
      -- CP-element group 32: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_156_Sample/req
      -- 
    req_339_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_339_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(32), ack => WPIPE_zeropad_output_pipe_156_inst_req_0); -- 
    sendOutput_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(22) & sendOutput_CP_26_elements(31);
      gj_sendOutput_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (6) 
      -- CP-element group 33: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_156_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_156_update_start_
      -- CP-element group 33: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_156_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_156_Sample/ack
      -- CP-element group 33: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_156_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_156_Update/req
      -- 
    ack_340_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_156_inst_ack_0, ack => sendOutput_CP_26_elements(33)); -- 
    req_344_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_344_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(33), ack => WPIPE_zeropad_output_pipe_156_inst_req_1); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_156_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_156_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_156_Update/ack
      -- 
    ack_345_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_156_inst_ack_1, ack => sendOutput_CP_26_elements(34)); -- 
    -- CP-element group 35:  join  transition  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: 	20 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_159_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_159_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_159_Sample/req
      -- 
    req_353_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_353_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(35), ack => WPIPE_zeropad_output_pipe_159_inst_req_0); -- 
    sendOutput_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(34) & sendOutput_CP_26_elements(20);
      gj_sendOutput_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  transition  input  output  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	37 
    -- CP-element group 36:  members (6) 
      -- CP-element group 36: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_159_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_159_update_start_
      -- CP-element group 36: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_159_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_159_Sample/ack
      -- CP-element group 36: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_159_Update/$entry
      -- CP-element group 36: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_159_Update/req
      -- 
    ack_354_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_159_inst_ack_0, ack => sendOutput_CP_26_elements(36)); -- 
    req_358_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_358_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(36), ack => WPIPE_zeropad_output_pipe_159_inst_req_1); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	36 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_159_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_159_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_159_Update/ack
      -- 
    ack_359_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_159_inst_ack_1, ack => sendOutput_CP_26_elements(37)); -- 
    -- CP-element group 38:  join  transition  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: 	18 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_162_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_162_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_162_Sample/req
      -- 
    req_367_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_367_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(38), ack => WPIPE_zeropad_output_pipe_162_inst_req_0); -- 
    sendOutput_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(37) & sendOutput_CP_26_elements(18);
      gj_sendOutput_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  transition  input  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (6) 
      -- CP-element group 39: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_162_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_162_update_start_
      -- CP-element group 39: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_162_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_162_Sample/ack
      -- CP-element group 39: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_162_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_162_Update/req
      -- 
    ack_368_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_162_inst_ack_0, ack => sendOutput_CP_26_elements(39)); -- 
    req_372_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_372_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(39), ack => WPIPE_zeropad_output_pipe_162_inst_req_1); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_162_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_162_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_162_Update/ack
      -- 
    ack_373_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_162_inst_ack_1, ack => sendOutput_CP_26_elements(40)); -- 
    -- CP-element group 41:  join  transition  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	40 
    -- CP-element group 41: 	16 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_165_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_165_Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_165_Sample/req
      -- 
    req_381_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_381_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(41), ack => WPIPE_zeropad_output_pipe_165_inst_req_0); -- 
    sendOutput_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(40) & sendOutput_CP_26_elements(16);
      gj_sendOutput_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (6) 
      -- CP-element group 42: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_165_Update/req
      -- CP-element group 42: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_165_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_165_update_start_
      -- CP-element group 42: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_165_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_165_Sample/ack
      -- CP-element group 42: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_165_Update/$entry
      -- 
    ack_382_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_165_inst_ack_0, ack => sendOutput_CP_26_elements(42)); -- 
    req_386_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_386_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(42), ack => WPIPE_zeropad_output_pipe_165_inst_req_1); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_165_Update/ack
      -- CP-element group 43: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_165_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_165_Update/$exit
      -- 
    ack_387_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_165_inst_ack_1, ack => sendOutput_CP_26_elements(43)); -- 
    -- CP-element group 44:  join  transition  output  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: 	14 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_168_sample_start_
      -- CP-element group 44: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_168_Sample/$entry
      -- CP-element group 44: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_168_Sample/req
      -- 
    req_395_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_395_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(44), ack => WPIPE_zeropad_output_pipe_168_inst_req_0); -- 
    sendOutput_cp_element_group_44: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_44"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(43) & sendOutput_CP_26_elements(14);
      gj_sendOutput_cp_element_group_44 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(44), clk => clk, reset => reset); --
    end block;
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	44 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (6) 
      -- CP-element group 45: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_168_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_168_update_start_
      -- CP-element group 45: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_168_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_168_Sample/ack
      -- CP-element group 45: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_168_Update/$entry
      -- CP-element group 45: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_168_Update/req
      -- 
    ack_396_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_168_inst_ack_0, ack => sendOutput_CP_26_elements(45)); -- 
    req_400_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_400_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(45), ack => WPIPE_zeropad_output_pipe_168_inst_req_1); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_168_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_168_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_168_Update/ack
      -- 
    ack_401_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_168_inst_ack_1, ack => sendOutput_CP_26_elements(46)); -- 
    -- CP-element group 47:  join  transition  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: 	12 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_171_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_171_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_171_Sample/req
      -- 
    req_409_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_409_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(47), ack => WPIPE_zeropad_output_pipe_171_inst_req_0); -- 
    sendOutput_cp_element_group_47: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_47"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(46) & sendOutput_CP_26_elements(12);
      gj_sendOutput_cp_element_group_47 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(47), clk => clk, reset => reset); --
    end block;
    -- CP-element group 48:  transition  input  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (6) 
      -- CP-element group 48: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_171_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_171_update_start_
      -- CP-element group 48: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_171_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_171_Sample/ack
      -- CP-element group 48: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_171_Update/$entry
      -- CP-element group 48: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_171_Update/req
      -- 
    ack_410_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_171_inst_ack_0, ack => sendOutput_CP_26_elements(48)); -- 
    req_414_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_414_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(48), ack => WPIPE_zeropad_output_pipe_171_inst_req_1); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_171_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_171_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/WPIPE_zeropad_output_pipe_171_Update/ack
      -- 
    ack_415_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_171_inst_ack_1, ack => sendOutput_CP_26_elements(49)); -- 
    -- CP-element group 50:  branch  join  transition  place  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: 	5 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (10) 
      -- CP-element group 50: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184__exit__
      -- CP-element group 50: 	 branch_block_stmt_24/if_stmt_185__entry__
      -- CP-element group 50: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/$exit
      -- CP-element group 50: 	 branch_block_stmt_24/if_stmt_185_dead_link/$entry
      -- CP-element group 50: 	 branch_block_stmt_24/if_stmt_185_eval_test/$entry
      -- CP-element group 50: 	 branch_block_stmt_24/if_stmt_185_eval_test/$exit
      -- CP-element group 50: 	 branch_block_stmt_24/if_stmt_185_eval_test/branch_req
      -- CP-element group 50: 	 branch_block_stmt_24/R_exitcond2_186_place
      -- CP-element group 50: 	 branch_block_stmt_24/if_stmt_185_if_link/$entry
      -- CP-element group 50: 	 branch_block_stmt_24/if_stmt_185_else_link/$entry
      -- 
    branch_req_423_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_423_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(50), ack => if_stmt_185_branch_req_0); -- 
    sendOutput_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(49) & sendOutput_CP_26_elements(5);
      gj_sendOutput_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  merge  transition  place  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	59 
    -- CP-element group 51:  members (13) 
      -- CP-element group 51: 	 branch_block_stmt_24/merge_stmt_191__exit__
      -- CP-element group 51: 	 branch_block_stmt_24/forx_xendx_xloopexit_forx_xend
      -- CP-element group 51: 	 branch_block_stmt_24/if_stmt_185_if_link/$exit
      -- CP-element group 51: 	 branch_block_stmt_24/if_stmt_185_if_link/if_choice_transition
      -- CP-element group 51: 	 branch_block_stmt_24/forx_xbody_forx_xendx_xloopexit
      -- CP-element group 51: 	 branch_block_stmt_24/forx_xbody_forx_xendx_xloopexit_PhiReq/$entry
      -- CP-element group 51: 	 branch_block_stmt_24/forx_xbody_forx_xendx_xloopexit_PhiReq/$exit
      -- CP-element group 51: 	 branch_block_stmt_24/merge_stmt_191_PhiReqMerge
      -- CP-element group 51: 	 branch_block_stmt_24/merge_stmt_191_PhiAck/$entry
      -- CP-element group 51: 	 branch_block_stmt_24/merge_stmt_191_PhiAck/$exit
      -- CP-element group 51: 	 branch_block_stmt_24/merge_stmt_191_PhiAck/dummy
      -- CP-element group 51: 	 branch_block_stmt_24/forx_xendx_xloopexit_forx_xend_PhiReq/$entry
      -- CP-element group 51: 	 branch_block_stmt_24/forx_xendx_xloopexit_forx_xend_PhiReq/$exit
      -- 
    if_choice_transition_428_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_185_branch_ack_1, ack => sendOutput_CP_26_elements(51)); -- 
    -- CP-element group 52:  fork  transition  place  input  output  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52: 	55 
    -- CP-element group 52:  members (12) 
      -- CP-element group 52: 	 branch_block_stmt_24/if_stmt_185_else_link/$exit
      -- CP-element group 52: 	 branch_block_stmt_24/if_stmt_185_else_link/else_choice_transition
      -- CP-element group 52: 	 branch_block_stmt_24/forx_xbody_forx_xbody
      -- CP-element group 52: 	 branch_block_stmt_24/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 52: 	 branch_block_stmt_24/forx_xbody_forx_xbody_PhiReq/phi_stmt_57/$entry
      -- CP-element group 52: 	 branch_block_stmt_24/forx_xbody_forx_xbody_PhiReq/phi_stmt_57/phi_stmt_57_sources/$entry
      -- CP-element group 52: 	 branch_block_stmt_24/forx_xbody_forx_xbody_PhiReq/phi_stmt_57/phi_stmt_57_sources/type_cast_63/$entry
      -- CP-element group 52: 	 branch_block_stmt_24/forx_xbody_forx_xbody_PhiReq/phi_stmt_57/phi_stmt_57_sources/type_cast_63/SplitProtocol/$entry
      -- CP-element group 52: 	 branch_block_stmt_24/forx_xbody_forx_xbody_PhiReq/phi_stmt_57/phi_stmt_57_sources/type_cast_63/SplitProtocol/Sample/$entry
      -- CP-element group 52: 	 branch_block_stmt_24/forx_xbody_forx_xbody_PhiReq/phi_stmt_57/phi_stmt_57_sources/type_cast_63/SplitProtocol/Sample/rr
      -- CP-element group 52: 	 branch_block_stmt_24/forx_xbody_forx_xbody_PhiReq/phi_stmt_57/phi_stmt_57_sources/type_cast_63/SplitProtocol/Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_24/forx_xbody_forx_xbody_PhiReq/phi_stmt_57/phi_stmt_57_sources/type_cast_63/SplitProtocol/Update/cr
      -- 
    else_choice_transition_432_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_185_branch_ack_0, ack => sendOutput_CP_26_elements(52)); -- 
    rr_476_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_476_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(52), ack => type_cast_63_inst_req_0); -- 
    cr_481_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_481_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(52), ack => type_cast_63_inst_req_1); -- 
    -- CP-element group 53:  transition  output  delay-element  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	4 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	57 
    -- CP-element group 53:  members (5) 
      -- CP-element group 53: 	 branch_block_stmt_24/bbx_xnph_forx_xbody_PhiReq/$exit
      -- CP-element group 53: 	 branch_block_stmt_24/bbx_xnph_forx_xbody_PhiReq/phi_stmt_57/$exit
      -- CP-element group 53: 	 branch_block_stmt_24/bbx_xnph_forx_xbody_PhiReq/phi_stmt_57/phi_stmt_57_sources/$exit
      -- CP-element group 53: 	 branch_block_stmt_24/bbx_xnph_forx_xbody_PhiReq/phi_stmt_57/phi_stmt_57_sources/type_cast_61_konst_delay_trans
      -- CP-element group 53: 	 branch_block_stmt_24/bbx_xnph_forx_xbody_PhiReq/phi_stmt_57/phi_stmt_57_req
      -- 
    phi_stmt_57_req_457_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_57_req_457_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(53), ack => phi_stmt_57_req_0); -- 
    -- Element group sendOutput_CP_26_elements(53) is a control-delay.
    cp_element_53_delay: control_delay_element  generic map(name => " 53_delay", delay_value => 1)  port map(req => sendOutput_CP_26_elements(4), ack => sendOutput_CP_26_elements(53), clk => clk, reset =>reset);
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	56 
    -- CP-element group 54:  members (2) 
      -- CP-element group 54: 	 branch_block_stmt_24/forx_xbody_forx_xbody_PhiReq/phi_stmt_57/phi_stmt_57_sources/type_cast_63/SplitProtocol/Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_24/forx_xbody_forx_xbody_PhiReq/phi_stmt_57/phi_stmt_57_sources/type_cast_63/SplitProtocol/Sample/ra
      -- 
    ra_477_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_63_inst_ack_0, ack => sendOutput_CP_26_elements(54)); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	52 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (2) 
      -- CP-element group 55: 	 branch_block_stmt_24/forx_xbody_forx_xbody_PhiReq/phi_stmt_57/phi_stmt_57_sources/type_cast_63/SplitProtocol/Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_24/forx_xbody_forx_xbody_PhiReq/phi_stmt_57/phi_stmt_57_sources/type_cast_63/SplitProtocol/Update/ca
      -- 
    ca_482_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_63_inst_ack_1, ack => sendOutput_CP_26_elements(55)); -- 
    -- CP-element group 56:  join  transition  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	54 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (6) 
      -- CP-element group 56: 	 branch_block_stmt_24/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 56: 	 branch_block_stmt_24/forx_xbody_forx_xbody_PhiReq/phi_stmt_57/$exit
      -- CP-element group 56: 	 branch_block_stmt_24/forx_xbody_forx_xbody_PhiReq/phi_stmt_57/phi_stmt_57_sources/$exit
      -- CP-element group 56: 	 branch_block_stmt_24/forx_xbody_forx_xbody_PhiReq/phi_stmt_57/phi_stmt_57_sources/type_cast_63/$exit
      -- CP-element group 56: 	 branch_block_stmt_24/forx_xbody_forx_xbody_PhiReq/phi_stmt_57/phi_stmt_57_sources/type_cast_63/SplitProtocol/$exit
      -- CP-element group 56: 	 branch_block_stmt_24/forx_xbody_forx_xbody_PhiReq/phi_stmt_57/phi_stmt_57_req
      -- 
    phi_stmt_57_req_483_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_57_req_483_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(56), ack => phi_stmt_57_req_1); -- 
    sendOutput_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_26_elements(54) & sendOutput_CP_26_elements(55);
      gj_sendOutput_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_26_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  merge  transition  place  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	53 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (2) 
      -- CP-element group 57: 	 branch_block_stmt_24/merge_stmt_56_PhiReqMerge
      -- CP-element group 57: 	 branch_block_stmt_24/merge_stmt_56_PhiAck/$entry
      -- 
    sendOutput_CP_26_elements(57) <= OrReduce(sendOutput_CP_26_elements(53) & sendOutput_CP_26_elements(56));
    -- CP-element group 58:  fork  transition  place  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	12 
    -- CP-element group 58: 	14 
    -- CP-element group 58: 	16 
    -- CP-element group 58: 	6 
    -- CP-element group 58: 	8 
    -- CP-element group 58: 	5 
    -- CP-element group 58: 	10 
    -- CP-element group 58: 	22 
    -- CP-element group 58: 	20 
    -- CP-element group 58: 	18 
    -- CP-element group 58: 	24 
    -- CP-element group 58: 	26 
    -- CP-element group 58:  members (53) 
      -- CP-element group 58: 	 branch_block_stmt_24/merge_stmt_56__exit__
      -- CP-element group 58: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184__entry__
      -- CP-element group 58: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_78_update_start_
      -- CP-element group 58: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/$entry
      -- CP-element group 58: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/addr_of_70_update_start_
      -- CP-element group 58: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/array_obj_ref_69_index_resized_1
      -- CP-element group 58: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/array_obj_ref_69_index_scaled_1
      -- CP-element group 58: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/array_obj_ref_69_index_computed_1
      -- CP-element group 58: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/array_obj_ref_69_index_resize_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/array_obj_ref_69_index_resize_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/array_obj_ref_69_index_resize_1/index_resize_req
      -- CP-element group 58: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/array_obj_ref_69_index_resize_1/index_resize_ack
      -- CP-element group 58: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/array_obj_ref_69_index_scale_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/array_obj_ref_69_index_scale_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/array_obj_ref_69_index_scale_1/scale_rename_req
      -- CP-element group 58: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/array_obj_ref_69_index_scale_1/scale_rename_ack
      -- CP-element group 58: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/array_obj_ref_69_final_index_sum_regn_update_start
      -- CP-element group 58: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/array_obj_ref_69_final_index_sum_regn_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/array_obj_ref_69_final_index_sum_regn_Sample/req
      -- CP-element group 58: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/array_obj_ref_69_final_index_sum_regn_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/array_obj_ref_69_final_index_sum_regn_Update/req
      -- CP-element group 58: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/addr_of_70_complete/$entry
      -- CP-element group 58: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/addr_of_70_complete/req
      -- CP-element group 58: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/ptr_deref_74_update_start_
      -- CP-element group 58: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/ptr_deref_74_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/ptr_deref_74_Update/word_access_complete/$entry
      -- CP-element group 58: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/ptr_deref_74_Update/word_access_complete/word_0/$entry
      -- CP-element group 58: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/ptr_deref_74_Update/word_access_complete/word_0/cr
      -- CP-element group 58: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_78_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_78_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_88_update_start_
      -- CP-element group 58: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_88_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_88_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_98_update_start_
      -- CP-element group 58: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_98_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_98_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_108_update_start_
      -- CP-element group 58: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_108_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_108_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_118_update_start_
      -- CP-element group 58: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_118_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_118_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_128_update_start_
      -- CP-element group 58: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_128_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_128_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_138_update_start_
      -- CP-element group 58: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_138_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_138_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_148_update_start_
      -- CP-element group 58: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_148_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_24/assign_stmt_71_to_assign_stmt_184/type_cast_148_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_24/merge_stmt_56_PhiAck/$exit
      -- CP-element group 58: 	 branch_block_stmt_24/merge_stmt_56_PhiAck/phi_stmt_57_ack
      -- 
    phi_stmt_57_ack_488_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_57_ack_0, ack => sendOutput_CP_26_elements(58)); -- 
    req_120_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_120_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(58), ack => array_obj_ref_69_index_offset_req_0); -- 
    req_125_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_125_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(58), ack => array_obj_ref_69_index_offset_req_1); -- 
    req_140_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_140_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(58), ack => addr_of_70_final_reg_req_1); -- 
    cr_185_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_185_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(58), ack => ptr_deref_74_load_0_req_1); -- 
    cr_204_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_204_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(58), ack => type_cast_78_inst_req_1); -- 
    cr_218_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_218_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(58), ack => type_cast_88_inst_req_1); -- 
    cr_232_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_232_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(58), ack => type_cast_98_inst_req_1); -- 
    cr_246_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_246_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(58), ack => type_cast_108_inst_req_1); -- 
    cr_260_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_260_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(58), ack => type_cast_118_inst_req_1); -- 
    cr_274_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_274_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(58), ack => type_cast_128_inst_req_1); -- 
    cr_288_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_288_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(58), ack => type_cast_138_inst_req_1); -- 
    cr_302_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_302_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_26_elements(58), ack => type_cast_148_inst_req_1); -- 
    -- CP-element group 59:  merge  transition  place  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	51 
    -- CP-element group 59: 	2 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (16) 
      -- CP-element group 59: 	 $exit
      -- CP-element group 59: 	 branch_block_stmt_24/$exit
      -- CP-element group 59: 	 branch_block_stmt_24/branch_block_stmt_24__exit__
      -- CP-element group 59: 	 branch_block_stmt_24/merge_stmt_193__exit__
      -- CP-element group 59: 	 branch_block_stmt_24/return__
      -- CP-element group 59: 	 branch_block_stmt_24/merge_stmt_195__exit__
      -- CP-element group 59: 	 branch_block_stmt_24/merge_stmt_193_PhiReqMerge
      -- CP-element group 59: 	 branch_block_stmt_24/merge_stmt_193_PhiAck/$entry
      -- CP-element group 59: 	 branch_block_stmt_24/merge_stmt_193_PhiAck/$exit
      -- CP-element group 59: 	 branch_block_stmt_24/merge_stmt_193_PhiAck/dummy
      -- CP-element group 59: 	 branch_block_stmt_24/return___PhiReq/$entry
      -- CP-element group 59: 	 branch_block_stmt_24/return___PhiReq/$exit
      -- CP-element group 59: 	 branch_block_stmt_24/merge_stmt_195_PhiReqMerge
      -- CP-element group 59: 	 branch_block_stmt_24/merge_stmt_195_PhiAck/$entry
      -- CP-element group 59: 	 branch_block_stmt_24/merge_stmt_195_PhiAck/$exit
      -- CP-element group 59: 	 branch_block_stmt_24/merge_stmt_195_PhiAck/dummy
      -- 
    sendOutput_CP_26_elements(59) <= OrReduce(sendOutput_CP_26_elements(51) & sendOutput_CP_26_elements(2));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i32_i32_32_wire : std_logic_vector(31 downto 0);
    signal R_indvar_68_resized : std_logic_vector(13 downto 0);
    signal R_indvar_68_scaled : std_logic_vector(13 downto 0);
    signal array_obj_ref_69_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_69_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_69_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_69_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_69_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_69_root_address : std_logic_vector(13 downto 0);
    signal arrayidx_71 : std_logic_vector(31 downto 0);
    signal cmp68_43 : std_logic_vector(0 downto 0);
    signal conv12_89 : std_logic_vector(7 downto 0);
    signal conv18_99 : std_logic_vector(7 downto 0);
    signal conv24_109 : std_logic_vector(7 downto 0);
    signal conv30_119 : std_logic_vector(7 downto 0);
    signal conv36_129 : std_logic_vector(7 downto 0);
    signal conv42_139 : std_logic_vector(7 downto 0);
    signal conv48_149 : std_logic_vector(7 downto 0);
    signal conv_79 : std_logic_vector(7 downto 0);
    signal exitcond2_184 : std_logic_vector(0 downto 0);
    signal indvar_57 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_179 : std_logic_vector(63 downto 0);
    signal ptr_deref_74_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_74_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_74_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_74_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_74_word_offset_0 : std_logic_vector(13 downto 0);
    signal shr15_95 : std_logic_vector(63 downto 0);
    signal shr21_105 : std_logic_vector(63 downto 0);
    signal shr27_115 : std_logic_vector(63 downto 0);
    signal shr33_125 : std_logic_vector(63 downto 0);
    signal shr39_135 : std_logic_vector(63 downto 0);
    signal shr45_145 : std_logic_vector(63 downto 0);
    signal shr67_34 : std_logic_vector(31 downto 0);
    signal shr9_85 : std_logic_vector(63 downto 0);
    signal tmp1_54 : std_logic_vector(63 downto 0);
    signal tmp4_75 : std_logic_vector(63 downto 0);
    signal type_cast_103_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_113_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_123_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_133_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_143_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_177_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_28_wire : std_logic_vector(31 downto 0);
    signal type_cast_31_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_37_wire : std_logic_vector(31 downto 0);
    signal type_cast_40_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_61_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_63_wire : std_logic_vector(63 downto 0);
    signal type_cast_83_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_93_wire_constant : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    array_obj_ref_69_constant_part_of_offset <= "00000000000000";
    array_obj_ref_69_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_69_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_69_resized_base_address <= "00000000000000";
    ptr_deref_74_word_offset_0 <= "00000000000000";
    type_cast_103_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_113_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_123_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_133_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_143_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_177_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_31_wire_constant <= "00000000000000000000000000000010";
    type_cast_40_wire_constant <= "00000000000000000000000000000000";
    type_cast_61_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_83_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_93_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    phi_stmt_57: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_61_wire_constant & type_cast_63_wire;
      req <= phi_stmt_57_req_0 & phi_stmt_57_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_57",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_57_ack_0,
          idata => idata,
          odata => indvar_57,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_57
    addr_of_70_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_70_final_reg_req_0;
      addr_of_70_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_70_final_reg_req_1;
      addr_of_70_final_reg_ack_1<= rack(0);
      addr_of_70_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_70_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_69_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_71,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_108_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_108_inst_req_0;
      type_cast_108_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_108_inst_req_1;
      type_cast_108_inst_ack_1<= rack(0);
      type_cast_108_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_108_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr21_105,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv24_109,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_118_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_118_inst_req_0;
      type_cast_118_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_118_inst_req_1;
      type_cast_118_inst_ack_1<= rack(0);
      type_cast_118_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_118_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr27_115,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv30_119,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_128_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_128_inst_req_0;
      type_cast_128_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_128_inst_req_1;
      type_cast_128_inst_ack_1<= rack(0);
      type_cast_128_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_128_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr33_125,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv36_129,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_138_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_138_inst_req_0;
      type_cast_138_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_138_inst_req_1;
      type_cast_138_inst_ack_1<= rack(0);
      type_cast_138_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_138_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr39_135,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv42_139,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_148_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_148_inst_req_0;
      type_cast_148_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_148_inst_req_1;
      type_cast_148_inst_ack_1<= rack(0);
      type_cast_148_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_148_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr45_145,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv48_149,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_28_inst
    process(size_buffer) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := size_buffer(31 downto 0);
      type_cast_28_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_33_inst
    process(ASHR_i32_i32_32_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_32_wire(31 downto 0);
      shr67_34 <= tmp_var; -- 
    end process;
    -- interlock type_cast_37_inst
    process(shr67_34) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := shr67_34(31 downto 0);
      type_cast_37_wire <= tmp_var; -- 
    end process;
    type_cast_53_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_53_inst_req_0;
      type_cast_53_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_53_inst_req_1;
      type_cast_53_inst_ack_1<= rack(0);
      type_cast_53_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_53_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr67_34,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp1_54,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_63_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_63_inst_req_0;
      type_cast_63_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_63_inst_req_1;
      type_cast_63_inst_ack_1<= rack(0);
      type_cast_63_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_63_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_179,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_63_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_78_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_78_inst_req_0;
      type_cast_78_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_78_inst_req_1;
      type_cast_78_inst_ack_1<= rack(0);
      type_cast_78_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_78_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp4_75,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_79,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_88_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_88_inst_req_0;
      type_cast_88_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_88_inst_req_1;
      type_cast_88_inst_ack_1<= rack(0);
      type_cast_88_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_88_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr9_85,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv12_89,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_98_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_98_inst_req_0;
      type_cast_98_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_98_inst_req_1;
      type_cast_98_inst_ack_1<= rack(0);
      type_cast_98_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_98_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr15_95,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv18_99,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_69_index_1_rename
    process(R_indvar_68_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_68_resized;
      ov(13 downto 0) := iv;
      R_indvar_68_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_69_index_1_resize
    process(indvar_57) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_57;
      ov := iv(13 downto 0);
      R_indvar_68_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_69_root_address_inst
    process(array_obj_ref_69_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_69_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_69_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_74_addr_0
    process(ptr_deref_74_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_74_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_74_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_74_base_resize
    process(arrayidx_71) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_71;
      ov := iv(13 downto 0);
      ptr_deref_74_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_74_gather_scatter
    process(ptr_deref_74_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_74_data_0;
      ov(63 downto 0) := iv;
      tmp4_75 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_74_root_address_inst
    process(ptr_deref_74_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_74_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_74_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_185_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond2_184;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_185_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_185_branch_req_0,
          ack0 => if_stmt_185_branch_ack_0,
          ack1 => if_stmt_185_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_44_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp68_43;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_44_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_44_branch_req_0,
          ack0 => if_stmt_44_branch_ack_0,
          ack1 => if_stmt_44_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u64_u64_178_inst
    process(indvar_57) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_57, type_cast_177_wire_constant, tmp_var);
      indvarx_xnext_179 <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_32_inst
    process(type_cast_28_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_28_wire, type_cast_31_wire_constant, tmp_var);
      ASHR_i32_i32_32_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_183_inst
    process(indvarx_xnext_179, tmp1_54) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_179, tmp1_54, tmp_var);
      exitcond2_184 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_104_inst
    process(tmp4_75) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_75, type_cast_103_wire_constant, tmp_var);
      shr21_105 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_114_inst
    process(tmp4_75) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_75, type_cast_113_wire_constant, tmp_var);
      shr27_115 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_124_inst
    process(tmp4_75) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_75, type_cast_123_wire_constant, tmp_var);
      shr33_125 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_134_inst
    process(tmp4_75) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_75, type_cast_133_wire_constant, tmp_var);
      shr39_135 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_144_inst
    process(tmp4_75) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_75, type_cast_143_wire_constant, tmp_var);
      shr45_145 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_84_inst
    process(tmp4_75) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_75, type_cast_83_wire_constant, tmp_var);
      shr9_85 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_94_inst
    process(tmp4_75) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_75, type_cast_93_wire_constant, tmp_var);
      shr15_95 <= tmp_var; --
    end process;
    -- binary operator SGT_i32_u1_41_inst
    process(type_cast_37_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(type_cast_37_wire, type_cast_40_wire_constant, tmp_var);
      cmp68_43 <= tmp_var; --
    end process;
    -- shared split operator group (11) : array_obj_ref_69_index_offset 
    ApIntAdd_group_11: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_68_scaled;
      array_obj_ref_69_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_69_index_offset_req_0;
      array_obj_ref_69_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_69_index_offset_req_1;
      array_obj_ref_69_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_11_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_11_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_11",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 11
    -- shared load operator group (0) : ptr_deref_74_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_74_load_0_req_0;
      ptr_deref_74_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_74_load_0_req_1;
      ptr_deref_74_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_74_word_address_0;
      ptr_deref_74_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(13 downto 0),
          mtag => memory_space_0_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared outport operator group (0) : WPIPE_zeropad_output_pipe_150_inst WPIPE_zeropad_output_pipe_153_inst WPIPE_zeropad_output_pipe_156_inst WPIPE_zeropad_output_pipe_159_inst WPIPE_zeropad_output_pipe_162_inst WPIPE_zeropad_output_pipe_165_inst WPIPE_zeropad_output_pipe_168_inst WPIPE_zeropad_output_pipe_171_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 7 downto 0);
      signal update_req, update_ack : BooleanArray( 7 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 7 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 7 downto 0);
      signal guard_vector : std_logic_vector( 7 downto 0);
      constant inBUFs : IntegerArray(7 downto 0) := (7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(7 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false);
      constant guardBuffering: IntegerArray(7 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2);
      -- 
    begin -- 
      sample_req_unguarded(7) <= WPIPE_zeropad_output_pipe_150_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_zeropad_output_pipe_153_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_zeropad_output_pipe_156_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_zeropad_output_pipe_159_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_zeropad_output_pipe_162_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_zeropad_output_pipe_165_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_zeropad_output_pipe_168_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_zeropad_output_pipe_171_inst_req_0;
      WPIPE_zeropad_output_pipe_150_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_zeropad_output_pipe_153_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_zeropad_output_pipe_156_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_zeropad_output_pipe_159_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_zeropad_output_pipe_162_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_zeropad_output_pipe_165_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_zeropad_output_pipe_168_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_zeropad_output_pipe_171_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(7) <= WPIPE_zeropad_output_pipe_150_inst_req_1;
      update_req_unguarded(6) <= WPIPE_zeropad_output_pipe_153_inst_req_1;
      update_req_unguarded(5) <= WPIPE_zeropad_output_pipe_156_inst_req_1;
      update_req_unguarded(4) <= WPIPE_zeropad_output_pipe_159_inst_req_1;
      update_req_unguarded(3) <= WPIPE_zeropad_output_pipe_162_inst_req_1;
      update_req_unguarded(2) <= WPIPE_zeropad_output_pipe_165_inst_req_1;
      update_req_unguarded(1) <= WPIPE_zeropad_output_pipe_168_inst_req_1;
      update_req_unguarded(0) <= WPIPE_zeropad_output_pipe_171_inst_req_1;
      WPIPE_zeropad_output_pipe_150_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_zeropad_output_pipe_153_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_zeropad_output_pipe_156_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_zeropad_output_pipe_159_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_zeropad_output_pipe_162_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_zeropad_output_pipe_165_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_zeropad_output_pipe_168_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_zeropad_output_pipe_171_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      data_in <= conv48_149 & conv42_139 & conv36_129 & conv30_119 & conv24_109 & conv18_99 & conv12_89 & conv_79;
      zeropad_output_pipe_write_0_gI: SplitGuardInterface generic map(name => "zeropad_output_pipe_write_0_gI", nreqs => 8, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      zeropad_output_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "zeropad_output_pipe", data_width => 8, num_reqs => 8, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => zeropad_output_pipe_pipe_write_req(0),
          oack => zeropad_output_pipe_pipe_write_ack(0),
          odata => zeropad_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end sendOutput_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timer is -- 
  generic (tag_length : integer); 
  port ( -- 
    c : out  std_logic_vector(63 downto 0);
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(0 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timer;
architecture timer_arch of timer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal c_buffer :  std_logic_vector(63 downto 0);
  signal c_update_enable: Boolean;
  signal timer_CP_520_start: Boolean;
  signal timer_CP_520_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal LOAD_count_201_load_0_req_0 : boolean;
  signal LOAD_count_201_load_0_ack_0 : boolean;
  signal LOAD_count_201_load_0_req_1 : boolean;
  signal LOAD_count_201_load_0_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timer_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timer_CP_520_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timer_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= c_buffer;
  c <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_520_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timer_CP_520_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_520_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timer_CP_520: Block -- control-path 
    signal timer_CP_520_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    timer_CP_520_elements(0) <= timer_CP_520_start;
    timer_CP_520_symbol <= timer_CP_520_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_202/$entry
      -- CP-element group 0: 	 assign_stmt_202/LOAD_count_201_sample_start_
      -- CP-element group 0: 	 assign_stmt_202/LOAD_count_201_update_start_
      -- CP-element group 0: 	 assign_stmt_202/LOAD_count_201_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_202/LOAD_count_201_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_202/LOAD_count_201_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_202/LOAD_count_201_Sample/word_access_start/$entry
      -- CP-element group 0: 	 assign_stmt_202/LOAD_count_201_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_202/LOAD_count_201_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 assign_stmt_202/LOAD_count_201_Update/$entry
      -- CP-element group 0: 	 assign_stmt_202/LOAD_count_201_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_202/LOAD_count_201_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_202/LOAD_count_201_Update/word_access_complete/word_0/cr
      -- 
    cr_552_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_552_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_520_elements(0), ack => LOAD_count_201_load_0_req_1); -- 
    rr_541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_520_elements(0), ack => LOAD_count_201_load_0_req_0); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (5) 
      -- CP-element group 1: 	 assign_stmt_202/LOAD_count_201_sample_completed_
      -- CP-element group 1: 	 assign_stmt_202/LOAD_count_201_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_202/LOAD_count_201_Sample/word_access_start/$exit
      -- CP-element group 1: 	 assign_stmt_202/LOAD_count_201_Sample/word_access_start/word_0/$exit
      -- CP-element group 1: 	 assign_stmt_202/LOAD_count_201_Sample/word_access_start/word_0/ra
      -- 
    ra_542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_count_201_load_0_ack_0, ack => timer_CP_520_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (11) 
      -- CP-element group 2: 	 $exit
      -- CP-element group 2: 	 assign_stmt_202/$exit
      -- CP-element group 2: 	 assign_stmt_202/LOAD_count_201_update_completed_
      -- CP-element group 2: 	 assign_stmt_202/LOAD_count_201_Update/$exit
      -- CP-element group 2: 	 assign_stmt_202/LOAD_count_201_Update/word_access_complete/$exit
      -- CP-element group 2: 	 assign_stmt_202/LOAD_count_201_Update/word_access_complete/word_0/$exit
      -- CP-element group 2: 	 assign_stmt_202/LOAD_count_201_Update/word_access_complete/word_0/ca
      -- CP-element group 2: 	 assign_stmt_202/LOAD_count_201_Update/LOAD_count_201_Merge/$entry
      -- CP-element group 2: 	 assign_stmt_202/LOAD_count_201_Update/LOAD_count_201_Merge/$exit
      -- CP-element group 2: 	 assign_stmt_202/LOAD_count_201_Update/LOAD_count_201_Merge/merge_req
      -- CP-element group 2: 	 assign_stmt_202/LOAD_count_201_Update/LOAD_count_201_Merge/merge_ack
      -- 
    ca_553_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_count_201_load_0_ack_1, ack => timer_CP_520_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal LOAD_count_201_data_0 : std_logic_vector(63 downto 0);
    signal LOAD_count_201_word_address_0 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    LOAD_count_201_word_address_0 <= "0";
    -- equivalence LOAD_count_201_gather_scatter
    process(LOAD_count_201_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_count_201_data_0;
      ov(63 downto 0) := iv;
      c_buffer <= ov(63 downto 0);
      --
    end process;
    -- shared load operator group (0) : LOAD_count_201_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_count_201_load_0_req_0;
      LOAD_count_201_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_count_201_load_0_req_1;
      LOAD_count_201_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_count_201_word_address_0;
      LOAD_count_201_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 0,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(0 downto 0),
          mtag => memory_space_2_lr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(63 downto 0),
          mtag => memory_space_2_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- 
  end Block; -- data_path
  -- 
end timer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity zeropad3D is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
    Block0_complete_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block0_complete_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block0_complete_pipe_read_data : in   std_logic_vector(7 downto 0);
    zeropad_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    zeropad_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    zeropad_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    zeropad_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    zeropad_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    zeropad_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    Block0_starting_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block0_starting_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block0_starting_pipe_write_data : out  std_logic_vector(7 downto 0);
    sendOutput_call_reqs : out  std_logic_vector(0 downto 0);
    sendOutput_call_acks : in   std_logic_vector(0 downto 0);
    sendOutput_call_data : out  std_logic_vector(31 downto 0);
    sendOutput_call_tag  :  out  std_logic_vector(0 downto 0);
    sendOutput_return_reqs : out  std_logic_vector(0 downto 0);
    sendOutput_return_acks : in   std_logic_vector(0 downto 0);
    sendOutput_return_tag :  in   std_logic_vector(0 downto 0);
    timer_call_reqs : out  std_logic_vector(0 downto 0);
    timer_call_acks : in   std_logic_vector(0 downto 0);
    timer_call_tag  :  out  std_logic_vector(1 downto 0);
    timer_return_reqs : out  std_logic_vector(0 downto 0);
    timer_return_acks : in   std_logic_vector(0 downto 0);
    timer_return_data : in   std_logic_vector(63 downto 0);
    timer_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity zeropad3D;
architecture zeropad3D_arch of zeropad3D is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal zeropad3D_CP_676_start: Boolean;
  signal zeropad3D_CP_676_symbol: Boolean;
  -- volatile/operator module components. 
  component sendOutput is -- 
    generic (tag_length : integer); 
    port ( -- 
      size : in  std_logic_vector(31 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
      zeropad_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      zeropad_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      zeropad_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      c : out  std_logic_vector(63 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal RPIPE_zeropad_input_pipe_238_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_226_inst_ack_1 : boolean;
  signal type_cast_305_inst_req_1 : boolean;
  signal type_cast_709_inst_ack_0 : boolean;
  signal type_cast_305_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_313_inst_req_0 : boolean;
  signal type_cast_689_inst_ack_0 : boolean;
  signal type_cast_292_inst_req_0 : boolean;
  signal type_cast_242_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_747_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_263_inst_req_0 : boolean;
  signal if_stmt_613_branch_ack_0 : boolean;
  signal type_cast_679_inst_req_1 : boolean;
  signal type_cast_729_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_226_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_226_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_747_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_235_inst_req_1 : boolean;
  signal type_cast_267_inst_ack_1 : boolean;
  signal WPIPE_Block0_starting_642_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_741_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_232_inst_ack_0 : boolean;
  signal type_cast_679_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_229_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_741_inst_req_1 : boolean;
  signal WPIPE_Block0_starting_642_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_235_inst_ack_0 : boolean;
  signal type_cast_267_inst_req_1 : boolean;
  signal WPIPE_Block0_starting_630_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_235_inst_req_0 : boolean;
  signal call_stmt_624_call_req_1 : boolean;
  signal type_cast_267_inst_ack_0 : boolean;
  signal WPIPE_Block0_starting_645_inst_req_1 : boolean;
  signal type_cast_267_inst_req_0 : boolean;
  signal type_cast_709_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_747_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_747_inst_ack_1 : boolean;
  signal call_stmt_624_call_req_0 : boolean;
  signal WPIPE_Block0_starting_642_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_226_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_753_inst_req_1 : boolean;
  signal WPIPE_Block0_starting_645_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_229_inst_ack_1 : boolean;
  signal WPIPE_Block0_starting_645_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_229_inst_req_1 : boolean;
  signal WPIPE_Block0_starting_642_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_232_inst_ack_1 : boolean;
  signal WPIPE_Block0_starting_630_inst_ack_0 : boolean;
  signal type_cast_679_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_232_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_741_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_313_inst_ack_1 : boolean;
  signal call_stmt_777_call_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_316_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_316_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_759_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_316_inst_req_1 : boolean;
  signal type_cast_709_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_316_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_238_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_229_inst_req_0 : boolean;
  signal call_stmt_624_call_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_238_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_232_inst_req_0 : boolean;
  signal type_cast_679_inst_ack_0 : boolean;
  signal call_stmt_624_call_ack_1 : boolean;
  signal type_cast_729_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_753_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_276_inst_ack_1 : boolean;
  signal WPIPE_Block0_starting_639_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_288_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_288_inst_ack_0 : boolean;
  signal WPIPE_Block0_starting_639_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_756_inst_ack_1 : boolean;
  signal type_cast_280_inst_ack_1 : boolean;
  signal type_cast_280_inst_req_1 : boolean;
  signal call_stmt_777_call_req_1 : boolean;
  signal type_cast_242_inst_ack_0 : boolean;
  signal type_cast_242_inst_req_0 : boolean;
  signal WPIPE_Block0_starting_645_inst_req_0 : boolean;
  signal type_cast_669_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_753_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_238_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_762_inst_ack_0 : boolean;
  signal type_cast_729_inst_req_0 : boolean;
  signal type_cast_255_inst_ack_1 : boolean;
  signal type_cast_255_inst_req_1 : boolean;
  signal type_cast_255_inst_ack_0 : boolean;
  signal type_cast_255_inst_req_0 : boolean;
  signal WPIPE_Block0_starting_639_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_276_inst_req_1 : boolean;
  signal type_cast_669_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_276_inst_req_0 : boolean;
  signal type_cast_709_inst_req_1 : boolean;
  signal type_cast_292_inst_ack_0 : boolean;
  signal type_cast_292_inst_req_1 : boolean;
  signal type_cast_292_inst_ack_1 : boolean;
  signal type_cast_669_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_753_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_263_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_288_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_288_inst_ack_1 : boolean;
  signal type_cast_729_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_251_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_251_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_741_inst_req_0 : boolean;
  signal WPIPE_Block0_starting_630_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_251_inst_ack_0 : boolean;
  signal type_cast_242_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_251_inst_req_0 : boolean;
  signal type_cast_628_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_301_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_756_inst_req_1 : boolean;
  signal call_stmt_777_call_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_313_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_313_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_301_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_301_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_301_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_263_inst_ack_1 : boolean;
  signal type_cast_280_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_263_inst_req_1 : boolean;
  signal type_cast_280_inst_req_0 : boolean;
  signal type_cast_689_inst_req_0 : boolean;
  signal type_cast_305_inst_ack_0 : boolean;
  signal WPIPE_Block0_starting_639_inst_ack_1 : boolean;
  signal type_cast_305_inst_req_0 : boolean;
  signal if_stmt_613_branch_ack_1 : boolean;
  signal type_cast_669_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_276_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_235_inst_ack_1 : boolean;
  signal WPIPE_Block0_starting_630_inst_ack_1 : boolean;
  signal type_cast_320_inst_req_0 : boolean;
  signal type_cast_320_inst_ack_0 : boolean;
  signal type_cast_320_inst_req_1 : boolean;
  signal type_cast_320_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_756_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_329_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_329_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_759_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_329_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_329_inst_ack_1 : boolean;
  signal call_stmt_777_call_req_0 : boolean;
  signal type_cast_333_inst_req_0 : boolean;
  signal type_cast_333_inst_ack_0 : boolean;
  signal type_cast_333_inst_req_1 : boolean;
  signal type_cast_333_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_756_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_341_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_341_inst_ack_0 : boolean;
  signal WPIPE_Block0_starting_636_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_341_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_341_inst_ack_1 : boolean;
  signal type_cast_660_inst_ack_1 : boolean;
  signal type_cast_345_inst_req_0 : boolean;
  signal type_cast_345_inst_ack_0 : boolean;
  signal type_cast_345_inst_req_1 : boolean;
  signal type_cast_345_inst_ack_1 : boolean;
  signal type_cast_739_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_354_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_354_inst_ack_0 : boolean;
  signal WPIPE_Block0_starting_636_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_759_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_354_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_354_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_750_inst_ack_1 : boolean;
  signal type_cast_660_inst_req_1 : boolean;
  signal WPIPE_zeropad_output_pipe_750_inst_req_1 : boolean;
  signal type_cast_358_inst_req_0 : boolean;
  signal type_cast_358_inst_ack_0 : boolean;
  signal type_cast_358_inst_req_1 : boolean;
  signal type_cast_358_inst_ack_1 : boolean;
  signal type_cast_739_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_366_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_366_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_759_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_366_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_366_inst_ack_1 : boolean;
  signal type_cast_660_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_744_inst_ack_1 : boolean;
  signal type_cast_370_inst_req_0 : boolean;
  signal type_cast_370_inst_ack_0 : boolean;
  signal type_cast_370_inst_req_1 : boolean;
  signal type_cast_370_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_379_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_379_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_379_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_379_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_762_inst_ack_1 : boolean;
  signal WPIPE_zeropad_output_pipe_750_inst_ack_0 : boolean;
  signal type_cast_719_inst_ack_1 : boolean;
  signal type_cast_660_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_744_inst_req_1 : boolean;
  signal type_cast_383_inst_req_0 : boolean;
  signal type_cast_383_inst_ack_0 : boolean;
  signal type_cast_383_inst_req_1 : boolean;
  signal type_cast_383_inst_ack_1 : boolean;
  signal WPIPE_Block0_starting_636_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_762_inst_req_0 : boolean;
  signal type_cast_628_inst_req_1 : boolean;
  signal if_stmt_422_branch_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_750_inst_req_0 : boolean;
  signal type_cast_689_inst_ack_1 : boolean;
  signal if_stmt_422_branch_ack_1 : boolean;
  signal type_cast_628_inst_ack_0 : boolean;
  signal if_stmt_422_branch_ack_0 : boolean;
  signal type_cast_689_inst_req_1 : boolean;
  signal type_cast_739_inst_ack_0 : boolean;
  signal type_cast_739_inst_req_0 : boolean;
  signal type_cast_719_inst_req_1 : boolean;
  signal type_cast_628_inst_req_0 : boolean;
  signal WPIPE_zeropad_output_pipe_762_inst_req_1 : boolean;
  signal call_stmt_656_call_ack_1 : boolean;
  signal array_obj_ref_462_index_offset_req_0 : boolean;
  signal array_obj_ref_462_index_offset_ack_0 : boolean;
  signal WPIPE_Block0_starting_636_inst_req_0 : boolean;
  signal array_obj_ref_462_index_offset_req_1 : boolean;
  signal array_obj_ref_462_index_offset_ack_1 : boolean;
  signal call_stmt_656_call_req_1 : boolean;
  signal type_cast_699_inst_ack_1 : boolean;
  signal addr_of_463_final_reg_req_0 : boolean;
  signal type_cast_699_inst_req_1 : boolean;
  signal addr_of_463_final_reg_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_744_inst_ack_0 : boolean;
  signal addr_of_463_final_reg_req_1 : boolean;
  signal addr_of_463_final_reg_ack_1 : boolean;
  signal type_cast_719_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_466_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_466_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_466_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_466_inst_ack_1 : boolean;
  signal call_stmt_656_call_ack_0 : boolean;
  signal call_stmt_656_call_req_0 : boolean;
  signal type_cast_470_inst_req_0 : boolean;
  signal type_cast_470_inst_ack_0 : boolean;
  signal WPIPE_zeropad_output_pipe_744_inst_req_0 : boolean;
  signal type_cast_470_inst_req_1 : boolean;
  signal type_cast_699_inst_ack_0 : boolean;
  signal type_cast_470_inst_ack_1 : boolean;
  signal if_stmt_613_branch_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_479_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_479_inst_ack_0 : boolean;
  signal WPIPE_Block0_starting_633_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_479_inst_req_1 : boolean;
  signal type_cast_699_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_479_inst_ack_1 : boolean;
  signal type_cast_483_inst_req_0 : boolean;
  signal type_cast_483_inst_ack_0 : boolean;
  signal type_cast_483_inst_req_1 : boolean;
  signal type_cast_483_inst_ack_1 : boolean;
  signal WPIPE_Block0_starting_633_inst_req_1 : boolean;
  signal type_cast_719_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_497_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_497_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_497_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_497_inst_ack_1 : boolean;
  signal RPIPE_Block0_complete_652_inst_ack_1 : boolean;
  signal RPIPE_Block0_complete_652_inst_req_1 : boolean;
  signal RPIPE_Block0_complete_652_inst_ack_0 : boolean;
  signal RPIPE_Block0_complete_652_inst_req_0 : boolean;
  signal type_cast_501_inst_req_0 : boolean;
  signal type_cast_501_inst_ack_0 : boolean;
  signal type_cast_501_inst_req_1 : boolean;
  signal type_cast_501_inst_ack_1 : boolean;
  signal WPIPE_Block0_starting_633_inst_ack_0 : boolean;
  signal WPIPE_Block0_starting_633_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_515_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_515_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_515_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_515_inst_ack_1 : boolean;
  signal type_cast_519_inst_req_0 : boolean;
  signal type_cast_519_inst_ack_0 : boolean;
  signal type_cast_519_inst_req_1 : boolean;
  signal type_cast_519_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_533_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_533_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_533_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_533_inst_ack_1 : boolean;
  signal WPIPE_Block0_starting_648_inst_ack_1 : boolean;
  signal WPIPE_Block0_starting_648_inst_req_1 : boolean;
  signal WPIPE_Block0_starting_648_inst_ack_0 : boolean;
  signal WPIPE_Block0_starting_648_inst_req_0 : boolean;
  signal type_cast_537_inst_req_0 : boolean;
  signal type_cast_537_inst_ack_0 : boolean;
  signal type_cast_537_inst_req_1 : boolean;
  signal type_cast_537_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_551_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_551_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_551_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_551_inst_ack_1 : boolean;
  signal type_cast_555_inst_req_0 : boolean;
  signal type_cast_555_inst_ack_0 : boolean;
  signal type_cast_555_inst_req_1 : boolean;
  signal type_cast_555_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_569_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_569_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_569_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_569_inst_ack_1 : boolean;
  signal type_cast_573_inst_req_0 : boolean;
  signal type_cast_573_inst_ack_0 : boolean;
  signal type_cast_573_inst_req_1 : boolean;
  signal type_cast_573_inst_ack_1 : boolean;
  signal RPIPE_zeropad_input_pipe_587_inst_req_0 : boolean;
  signal RPIPE_zeropad_input_pipe_587_inst_ack_0 : boolean;
  signal RPIPE_zeropad_input_pipe_587_inst_req_1 : boolean;
  signal RPIPE_zeropad_input_pipe_587_inst_ack_1 : boolean;
  signal type_cast_591_inst_req_0 : boolean;
  signal type_cast_591_inst_ack_0 : boolean;
  signal type_cast_591_inst_req_1 : boolean;
  signal type_cast_591_inst_ack_1 : boolean;
  signal ptr_deref_599_store_0_req_0 : boolean;
  signal ptr_deref_599_store_0_ack_0 : boolean;
  signal ptr_deref_599_store_0_req_1 : boolean;
  signal ptr_deref_599_store_0_ack_1 : boolean;
  signal phi_stmt_450_req_0 : boolean;
  signal type_cast_456_inst_req_0 : boolean;
  signal type_cast_456_inst_ack_0 : boolean;
  signal type_cast_456_inst_req_1 : boolean;
  signal type_cast_456_inst_ack_1 : boolean;
  signal phi_stmt_450_req_1 : boolean;
  signal phi_stmt_450_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "zeropad3D_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  zeropad3D_CP_676_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "zeropad3D_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= zeropad3D_CP_676_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= zeropad3D_CP_676_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= zeropad3D_CP_676_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  zeropad3D_CP_676: Block -- control-path 
    signal zeropad3D_CP_676_elements: BooleanArray(176 downto 0);
    -- 
  begin -- 
    zeropad3D_CP_676_elements(0) <= zeropad3D_CP_676_start;
    zeropad3D_CP_676_symbol <= zeropad3D_CP_676_elements(169);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	20 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	24 
    -- CP-element group 0: 	28 
    -- CP-element group 0: 	32 
    -- CP-element group 0: 	38 
    -- CP-element group 0: 	42 
    -- CP-element group 0: 	46 
    -- CP-element group 0: 	50 
    -- CP-element group 0: 	54 
    -- CP-element group 0: 	58 
    -- CP-element group 0: 	12 
    -- CP-element group 0: 	16 
    -- CP-element group 0:  members (44) 
      -- CP-element group 0: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_305_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_242_update_start_
      -- CP-element group 0: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_242_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_226_sample_start_
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_267_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_267_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_226_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421__entry__
      -- CP-element group 0: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_226_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_224/branch_block_stmt_224__entry__
      -- CP-element group 0: 	 branch_block_stmt_224/$entry
      -- CP-element group 0: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_292_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/$entry
      -- CP-element group 0: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_292_update_start_
      -- CP-element group 0: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_280_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_242_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_255_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_255_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_280_update_start_
      -- CP-element group 0: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_292_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_267_update_start_
      -- CP-element group 0: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_280_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_305_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_255_update_start_
      -- CP-element group 0: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_305_update_start_
      -- CP-element group 0: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_320_update_start_
      -- CP-element group 0: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_320_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_320_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_333_update_start_
      -- CP-element group 0: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_333_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_333_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_345_update_start_
      -- CP-element group 0: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_345_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_345_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_358_update_start_
      -- CP-element group 0: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_358_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_358_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_370_update_start_
      -- CP-element group 0: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_370_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_370_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_383_update_start_
      -- CP-element group 0: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_383_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_383_Update/cr
      -- 
    cr_935_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_935_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(0), ack => type_cast_305_inst_req_1); -- 
    cr_795_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_795_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(0), ack => type_cast_242_inst_req_1); -- 
    cr_851_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_851_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(0), ack => type_cast_267_inst_req_1); -- 
    rr_720_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_720_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(0), ack => RPIPE_zeropad_input_pipe_226_inst_req_0); -- 
    cr_879_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_879_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(0), ack => type_cast_280_inst_req_1); -- 
    cr_823_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_823_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(0), ack => type_cast_255_inst_req_1); -- 
    cr_907_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_907_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(0), ack => type_cast_292_inst_req_1); -- 
    cr_977_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_977_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(0), ack => type_cast_320_inst_req_1); -- 
    cr_1005_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1005_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(0), ack => type_cast_333_inst_req_1); -- 
    cr_1033_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1033_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(0), ack => type_cast_345_inst_req_1); -- 
    cr_1061_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1061_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(0), ack => type_cast_358_inst_req_1); -- 
    cr_1089_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1089_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(0), ack => type_cast_370_inst_req_1); -- 
    cr_1117_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1117_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(0), ack => type_cast_383_inst_req_1); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_226_Update/cr
      -- CP-element group 1: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_226_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_226_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_226_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_226_update_start_
      -- CP-element group 1: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_226_sample_completed_
      -- 
    ra_721_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_226_inst_ack_0, ack => zeropad3D_CP_676_elements(1)); -- 
    cr_725_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_725_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(1), ack => RPIPE_zeropad_input_pipe_226_inst_req_1); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_226_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_226_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_229_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_226_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_229_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_229_Sample/$entry
      -- 
    ca_726_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_226_inst_ack_1, ack => zeropad3D_CP_676_elements(2)); -- 
    rr_734_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_734_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(2), ack => RPIPE_zeropad_input_pipe_229_inst_req_0); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_229_update_start_
      -- CP-element group 3: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_229_Sample/ra
      -- CP-element group 3: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_229_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_229_Update/cr
      -- CP-element group 3: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_229_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_229_Sample/$exit
      -- 
    ra_735_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_229_inst_ack_0, ack => zeropad3D_CP_676_elements(3)); -- 
    cr_739_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_739_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(3), ack => RPIPE_zeropad_input_pipe_229_inst_req_1); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_232_sample_start_
      -- CP-element group 4: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_229_Update/ca
      -- CP-element group 4: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_229_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_232_Sample/rr
      -- CP-element group 4: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_232_Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_229_update_completed_
      -- 
    ca_740_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_229_inst_ack_1, ack => zeropad3D_CP_676_elements(4)); -- 
    rr_748_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_748_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(4), ack => RPIPE_zeropad_input_pipe_232_inst_req_0); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_232_update_start_
      -- CP-element group 5: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_232_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_232_Sample/ra
      -- CP-element group 5: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_232_Update/cr
      -- CP-element group 5: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_232_Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_232_Sample/$exit
      -- 
    ra_749_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_232_inst_ack_0, ack => zeropad3D_CP_676_elements(5)); -- 
    cr_753_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_753_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(5), ack => RPIPE_zeropad_input_pipe_232_inst_req_1); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_232_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_235_Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_235_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_232_Update/ca
      -- CP-element group 6: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_232_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_235_sample_start_
      -- 
    ca_754_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_232_inst_ack_1, ack => zeropad3D_CP_676_elements(6)); -- 
    rr_762_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_762_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(6), ack => RPIPE_zeropad_input_pipe_235_inst_req_0); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_235_Update/$entry
      -- CP-element group 7: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_235_Update/cr
      -- CP-element group 7: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_235_Sample/ra
      -- CP-element group 7: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_235_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_235_update_start_
      -- CP-element group 7: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_235_sample_completed_
      -- 
    ra_763_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_235_inst_ack_0, ack => zeropad3D_CP_676_elements(7)); -- 
    cr_767_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_767_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(7), ack => RPIPE_zeropad_input_pipe_235_inst_req_1); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_238_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_235_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_238_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_238_Sample/rr
      -- CP-element group 8: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_235_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_235_Update/ca
      -- 
    ca_768_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_235_inst_ack_1, ack => zeropad3D_CP_676_elements(8)); -- 
    rr_776_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_776_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(8), ack => RPIPE_zeropad_input_pipe_238_inst_req_0); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_238_Sample/ra
      -- CP-element group 9: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_238_update_start_
      -- CP-element group 9: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_238_Update/cr
      -- CP-element group 9: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_238_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_238_Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_238_Sample/$exit
      -- 
    ra_777_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_238_inst_ack_0, ack => zeropad3D_CP_676_elements(9)); -- 
    cr_781_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_781_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(9), ack => RPIPE_zeropad_input_pipe_238_inst_req_1); -- 
    -- CP-element group 10:  fork  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10: 	13 
    -- CP-element group 10:  members (9) 
      -- CP-element group 10: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_238_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_238_Update/ca
      -- CP-element group 10: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_238_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_242_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_242_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_251_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_251_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_251_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_242_sample_start_
      -- 
    ca_782_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_238_inst_ack_1, ack => zeropad3D_CP_676_elements(10)); -- 
    rr_790_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_790_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(10), ack => type_cast_242_inst_req_0); -- 
    rr_804_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_804_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(10), ack => RPIPE_zeropad_input_pipe_251_inst_req_0); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_242_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_242_Sample/ra
      -- CP-element group 11: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_242_Sample/$exit
      -- 
    ra_791_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_242_inst_ack_0, ack => zeropad3D_CP_676_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	0 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	59 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_242_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_242_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_242_Update/ca
      -- 
    ca_796_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_242_inst_ack_1, ack => zeropad3D_CP_676_elements(12)); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	10 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_251_update_start_
      -- CP-element group 13: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_251_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_251_Update/cr
      -- CP-element group 13: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_251_Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_251_Sample/ra
      -- CP-element group 13: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_251_Sample/$exit
      -- 
    ra_805_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_251_inst_ack_0, ack => zeropad3D_CP_676_elements(13)); -- 
    cr_809_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_809_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(13), ack => RPIPE_zeropad_input_pipe_251_inst_req_1); -- 
    -- CP-element group 14:  fork  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	17 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (9) 
      -- CP-element group 14: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_263_Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_263_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_255_Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_255_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_251_Update/ca
      -- CP-element group 14: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_251_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_263_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_255_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_251_update_completed_
      -- 
    ca_810_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_251_inst_ack_1, ack => zeropad3D_CP_676_elements(14)); -- 
    rr_818_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_818_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(14), ack => type_cast_255_inst_req_0); -- 
    rr_832_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_832_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(14), ack => RPIPE_zeropad_input_pipe_263_inst_req_0); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_255_Sample/ra
      -- CP-element group 15: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_255_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_255_sample_completed_
      -- 
    ra_819_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_255_inst_ack_0, ack => zeropad3D_CP_676_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	0 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	59 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_255_Update/ca
      -- CP-element group 16: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_255_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_255_update_completed_
      -- 
    ca_824_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_255_inst_ack_1, ack => zeropad3D_CP_676_elements(16)); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	14 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_263_update_start_
      -- CP-element group 17: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_263_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_263_Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_263_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_263_Update/cr
      -- CP-element group 17: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_263_Update/$entry
      -- 
    ra_833_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_263_inst_ack_0, ack => zeropad3D_CP_676_elements(17)); -- 
    cr_837_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_837_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(17), ack => RPIPE_zeropad_input_pipe_263_inst_req_1); -- 
    -- CP-element group 18:  fork  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18: 	21 
    -- CP-element group 18:  members (9) 
      -- CP-element group 18: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_263_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_267_Sample/rr
      -- CP-element group 18: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_267_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_276_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_267_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_276_Sample/rr
      -- CP-element group 18: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_276_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_263_Update/ca
      -- CP-element group 18: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_263_Update/$exit
      -- 
    ca_838_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_263_inst_ack_1, ack => zeropad3D_CP_676_elements(18)); -- 
    rr_846_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_846_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(18), ack => type_cast_267_inst_req_0); -- 
    rr_860_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_860_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(18), ack => RPIPE_zeropad_input_pipe_276_inst_req_0); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_267_Sample/ra
      -- CP-element group 19: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_267_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_267_sample_completed_
      -- 
    ra_847_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_267_inst_ack_0, ack => zeropad3D_CP_676_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	0 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	59 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_267_Update/ca
      -- CP-element group 20: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_267_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_267_update_completed_
      -- 
    ca_852_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_267_inst_ack_1, ack => zeropad3D_CP_676_elements(20)); -- 
    -- CP-element group 21:  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	18 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (6) 
      -- CP-element group 21: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_276_Update/$entry
      -- CP-element group 21: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_276_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_276_Update/cr
      -- CP-element group 21: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_276_update_start_
      -- CP-element group 21: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_276_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_276_Sample/ra
      -- 
    ra_861_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_276_inst_ack_0, ack => zeropad3D_CP_676_elements(21)); -- 
    cr_865_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_865_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(21), ack => RPIPE_zeropad_input_pipe_276_inst_req_1); -- 
    -- CP-element group 22:  fork  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22: 	25 
    -- CP-element group 22:  members (9) 
      -- CP-element group 22: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_280_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_276_Update/ca
      -- CP-element group 22: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_288_Sample/rr
      -- CP-element group 22: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_288_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_276_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_288_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_276_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_280_Sample/rr
      -- CP-element group 22: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_280_Sample/$entry
      -- 
    ca_866_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_276_inst_ack_1, ack => zeropad3D_CP_676_elements(22)); -- 
    rr_874_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_874_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(22), ack => type_cast_280_inst_req_0); -- 
    rr_888_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_888_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(22), ack => RPIPE_zeropad_input_pipe_288_inst_req_0); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_280_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_280_Sample/ra
      -- CP-element group 23: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_280_Sample/$exit
      -- 
    ra_875_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_280_inst_ack_0, ack => zeropad3D_CP_676_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	0 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	59 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_280_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_280_Update/ca
      -- CP-element group 24: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_280_Update/$exit
      -- 
    ca_880_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_280_inst_ack_1, ack => zeropad3D_CP_676_elements(24)); -- 
    -- CP-element group 25:  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	22 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25:  members (6) 
      -- CP-element group 25: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_288_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_288_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_288_Sample/ra
      -- CP-element group 25: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_288_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_288_Update/cr
      -- CP-element group 25: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_288_update_start_
      -- 
    ra_889_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_288_inst_ack_0, ack => zeropad3D_CP_676_elements(25)); -- 
    cr_893_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_893_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(25), ack => RPIPE_zeropad_input_pipe_288_inst_req_1); -- 
    -- CP-element group 26:  fork  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: 	29 
    -- CP-element group 26:  members (9) 
      -- CP-element group 26: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_292_Sample/rr
      -- CP-element group 26: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_288_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_301_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_292_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_288_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_292_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_288_Update/ca
      -- CP-element group 26: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_301_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_301_Sample/rr
      -- 
    ca_894_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_288_inst_ack_1, ack => zeropad3D_CP_676_elements(26)); -- 
    rr_902_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_902_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(26), ack => type_cast_292_inst_req_0); -- 
    rr_916_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_916_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(26), ack => RPIPE_zeropad_input_pipe_301_inst_req_0); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_292_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_292_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_292_Sample/ra
      -- 
    ra_903_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_292_inst_ack_0, ack => zeropad3D_CP_676_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	0 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	59 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_292_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_292_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_292_Update/ca
      -- 
    ca_908_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_292_inst_ack_1, ack => zeropad3D_CP_676_elements(28)); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	26 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_301_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_301_update_start_
      -- CP-element group 29: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_301_Sample/ra
      -- CP-element group 29: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_301_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_301_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_301_Update/cr
      -- 
    ra_917_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_301_inst_ack_0, ack => zeropad3D_CP_676_elements(29)); -- 
    cr_921_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_921_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(29), ack => RPIPE_zeropad_input_pipe_301_inst_req_1); -- 
    -- CP-element group 30:  fork  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30: 	33 
    -- CP-element group 30:  members (9) 
      -- CP-element group 30: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_313_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_313_Sample/rr
      -- CP-element group 30: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_301_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_301_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_301_Update/ca
      -- CP-element group 30: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_313_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_305_Sample/rr
      -- CP-element group 30: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_305_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_305_sample_start_
      -- 
    ca_922_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_301_inst_ack_1, ack => zeropad3D_CP_676_elements(30)); -- 
    rr_930_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_930_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(30), ack => type_cast_305_inst_req_0); -- 
    rr_944_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_944_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(30), ack => RPIPE_zeropad_input_pipe_313_inst_req_0); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_305_Sample/ra
      -- CP-element group 31: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_305_Sample/$exit
      -- CP-element group 31: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_305_sample_completed_
      -- 
    ra_931_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_305_inst_ack_0, ack => zeropad3D_CP_676_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	0 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	59 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_305_Update/ca
      -- CP-element group 32: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_305_Update/$exit
      -- CP-element group 32: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_305_update_completed_
      -- 
    ca_936_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_305_inst_ack_1, ack => zeropad3D_CP_676_elements(32)); -- 
    -- CP-element group 33:  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	30 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (6) 
      -- CP-element group 33: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_313_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_313_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_313_update_start_
      -- CP-element group 33: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_313_Sample/ra
      -- CP-element group 33: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_313_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_313_Update/cr
      -- 
    ra_945_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_313_inst_ack_0, ack => zeropad3D_CP_676_elements(33)); -- 
    cr_949_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_949_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(33), ack => RPIPE_zeropad_input_pipe_313_inst_req_1); -- 
    -- CP-element group 34:  transition  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34:  members (6) 
      -- CP-element group 34: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_313_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_313_Update/ca
      -- CP-element group 34: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_316_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_316_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_316_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_313_Update/$exit
      -- 
    ca_950_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_313_inst_ack_1, ack => zeropad3D_CP_676_elements(34)); -- 
    rr_958_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_958_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(34), ack => RPIPE_zeropad_input_pipe_316_inst_req_0); -- 
    -- CP-element group 35:  transition  input  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (6) 
      -- CP-element group 35: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_316_update_start_
      -- CP-element group 35: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_316_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_316_Sample/ra
      -- CP-element group 35: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_316_Update/$entry
      -- CP-element group 35: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_316_Update/cr
      -- CP-element group 35: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_316_sample_completed_
      -- 
    ra_959_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_316_inst_ack_0, ack => zeropad3D_CP_676_elements(35)); -- 
    cr_963_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_963_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(35), ack => RPIPE_zeropad_input_pipe_316_inst_req_1); -- 
    -- CP-element group 36:  fork  transition  input  output  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	37 
    -- CP-element group 36: 	39 
    -- CP-element group 36:  members (9) 
      -- CP-element group 36: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_316_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_316_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_316_Update/ca
      -- CP-element group 36: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_320_sample_start_
      -- CP-element group 36: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_320_Sample/$entry
      -- CP-element group 36: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_320_Sample/rr
      -- CP-element group 36: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_329_sample_start_
      -- CP-element group 36: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_329_Sample/$entry
      -- CP-element group 36: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_329_Sample/rr
      -- 
    ca_964_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_316_inst_ack_1, ack => zeropad3D_CP_676_elements(36)); -- 
    rr_972_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_972_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(36), ack => type_cast_320_inst_req_0); -- 
    rr_986_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_986_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(36), ack => RPIPE_zeropad_input_pipe_329_inst_req_0); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	36 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_320_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_320_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_320_Sample/ra
      -- 
    ra_973_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_320_inst_ack_0, ack => zeropad3D_CP_676_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	0 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	59 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_320_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_320_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_320_Update/ca
      -- 
    ca_978_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_320_inst_ack_1, ack => zeropad3D_CP_676_elements(38)); -- 
    -- CP-element group 39:  transition  input  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	36 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (6) 
      -- CP-element group 39: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_329_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_329_update_start_
      -- CP-element group 39: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_329_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_329_Sample/ra
      -- CP-element group 39: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_329_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_329_Update/cr
      -- 
    ra_987_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_329_inst_ack_0, ack => zeropad3D_CP_676_elements(39)); -- 
    cr_991_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_991_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(39), ack => RPIPE_zeropad_input_pipe_329_inst_req_1); -- 
    -- CP-element group 40:  fork  transition  input  output  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40: 	43 
    -- CP-element group 40:  members (9) 
      -- CP-element group 40: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_329_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_329_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_329_Update/ca
      -- CP-element group 40: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_333_sample_start_
      -- CP-element group 40: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_333_Sample/$entry
      -- CP-element group 40: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_333_Sample/rr
      -- CP-element group 40: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_341_sample_start_
      -- CP-element group 40: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_341_Sample/$entry
      -- CP-element group 40: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_341_Sample/rr
      -- 
    ca_992_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_329_inst_ack_1, ack => zeropad3D_CP_676_elements(40)); -- 
    rr_1000_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1000_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(40), ack => type_cast_333_inst_req_0); -- 
    rr_1014_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1014_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(40), ack => RPIPE_zeropad_input_pipe_341_inst_req_0); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_333_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_333_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_333_Sample/ra
      -- 
    ra_1001_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_333_inst_ack_0, ack => zeropad3D_CP_676_elements(41)); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	0 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	59 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_333_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_333_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_333_Update/ca
      -- 
    ca_1006_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_333_inst_ack_1, ack => zeropad3D_CP_676_elements(42)); -- 
    -- CP-element group 43:  transition  input  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	40 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (6) 
      -- CP-element group 43: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_341_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_341_update_start_
      -- CP-element group 43: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_341_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_341_Sample/ra
      -- CP-element group 43: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_341_Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_341_Update/cr
      -- 
    ra_1015_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_341_inst_ack_0, ack => zeropad3D_CP_676_elements(43)); -- 
    cr_1019_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1019_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(43), ack => RPIPE_zeropad_input_pipe_341_inst_req_1); -- 
    -- CP-element group 44:  fork  transition  input  output  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44: 	47 
    -- CP-element group 44:  members (9) 
      -- CP-element group 44: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_341_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_341_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_341_Update/ca
      -- CP-element group 44: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_345_sample_start_
      -- CP-element group 44: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_345_Sample/$entry
      -- CP-element group 44: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_345_Sample/rr
      -- CP-element group 44: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_354_sample_start_
      -- CP-element group 44: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_354_Sample/$entry
      -- CP-element group 44: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_354_Sample/rr
      -- 
    ca_1020_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_341_inst_ack_1, ack => zeropad3D_CP_676_elements(44)); -- 
    rr_1028_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1028_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(44), ack => type_cast_345_inst_req_0); -- 
    rr_1042_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1042_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(44), ack => RPIPE_zeropad_input_pipe_354_inst_req_0); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	44 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_345_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_345_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_345_Sample/ra
      -- 
    ra_1029_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_345_inst_ack_0, ack => zeropad3D_CP_676_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	0 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	59 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_345_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_345_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_345_Update/ca
      -- 
    ca_1034_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_345_inst_ack_1, ack => zeropad3D_CP_676_elements(46)); -- 
    -- CP-element group 47:  transition  input  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	44 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (6) 
      -- CP-element group 47: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_354_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_354_update_start_
      -- CP-element group 47: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_354_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_354_Sample/ra
      -- CP-element group 47: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_354_Update/$entry
      -- CP-element group 47: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_354_Update/cr
      -- 
    ra_1043_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_354_inst_ack_0, ack => zeropad3D_CP_676_elements(47)); -- 
    cr_1047_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1047_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(47), ack => RPIPE_zeropad_input_pipe_354_inst_req_1); -- 
    -- CP-element group 48:  fork  transition  input  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48: 	51 
    -- CP-element group 48:  members (9) 
      -- CP-element group 48: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_354_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_354_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_354_Update/ca
      -- CP-element group 48: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_358_sample_start_
      -- CP-element group 48: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_358_Sample/$entry
      -- CP-element group 48: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_358_Sample/rr
      -- CP-element group 48: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_366_sample_start_
      -- CP-element group 48: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_366_Sample/$entry
      -- CP-element group 48: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_366_Sample/rr
      -- 
    ca_1048_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_354_inst_ack_1, ack => zeropad3D_CP_676_elements(48)); -- 
    rr_1056_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1056_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(48), ack => type_cast_358_inst_req_0); -- 
    rr_1070_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1070_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(48), ack => RPIPE_zeropad_input_pipe_366_inst_req_0); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_358_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_358_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_358_Sample/ra
      -- 
    ra_1057_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_358_inst_ack_0, ack => zeropad3D_CP_676_elements(49)); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	0 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	59 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_358_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_358_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_358_Update/ca
      -- 
    ca_1062_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_358_inst_ack_1, ack => zeropad3D_CP_676_elements(50)); -- 
    -- CP-element group 51:  transition  input  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	48 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (6) 
      -- CP-element group 51: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_366_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_366_update_start_
      -- CP-element group 51: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_366_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_366_Sample/ra
      -- CP-element group 51: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_366_Update/$entry
      -- CP-element group 51: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_366_Update/cr
      -- 
    ra_1071_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_366_inst_ack_0, ack => zeropad3D_CP_676_elements(51)); -- 
    cr_1075_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1075_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(51), ack => RPIPE_zeropad_input_pipe_366_inst_req_1); -- 
    -- CP-element group 52:  fork  transition  input  output  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	53 
    -- CP-element group 52: 	55 
    -- CP-element group 52:  members (9) 
      -- CP-element group 52: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_366_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_366_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_366_Update/ca
      -- CP-element group 52: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_370_sample_start_
      -- CP-element group 52: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_370_Sample/$entry
      -- CP-element group 52: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_370_Sample/rr
      -- CP-element group 52: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_379_sample_start_
      -- CP-element group 52: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_379_Sample/$entry
      -- CP-element group 52: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_379_Sample/rr
      -- 
    ca_1076_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_366_inst_ack_1, ack => zeropad3D_CP_676_elements(52)); -- 
    rr_1084_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1084_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(52), ack => type_cast_370_inst_req_0); -- 
    rr_1098_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1098_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(52), ack => RPIPE_zeropad_input_pipe_379_inst_req_0); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	52 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_370_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_370_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_370_Sample/ra
      -- 
    ra_1085_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_370_inst_ack_0, ack => zeropad3D_CP_676_elements(53)); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	0 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	59 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_370_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_370_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_370_Update/ca
      -- 
    ca_1090_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_370_inst_ack_1, ack => zeropad3D_CP_676_elements(54)); -- 
    -- CP-element group 55:  transition  input  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	52 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (6) 
      -- CP-element group 55: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_379_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_379_update_start_
      -- CP-element group 55: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_379_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_379_Sample/ra
      -- CP-element group 55: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_379_Update/$entry
      -- CP-element group 55: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_379_Update/cr
      -- 
    ra_1099_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_379_inst_ack_0, ack => zeropad3D_CP_676_elements(55)); -- 
    cr_1103_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1103_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(55), ack => RPIPE_zeropad_input_pipe_379_inst_req_1); -- 
    -- CP-element group 56:  transition  input  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (6) 
      -- CP-element group 56: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_379_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_379_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/RPIPE_zeropad_input_pipe_379_Update/ca
      -- CP-element group 56: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_383_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_383_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_383_Sample/rr
      -- 
    ca_1104_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_379_inst_ack_1, ack => zeropad3D_CP_676_elements(56)); -- 
    rr_1112_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1112_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(56), ack => type_cast_383_inst_req_0); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_383_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_383_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_383_Sample/ra
      -- 
    ra_1113_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_383_inst_ack_0, ack => zeropad3D_CP_676_elements(57)); -- 
    -- CP-element group 58:  transition  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	0 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_383_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_383_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/type_cast_383_Update/ca
      -- 
    ca_1118_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_383_inst_ack_1, ack => zeropad3D_CP_676_elements(58)); -- 
    -- CP-element group 59:  branch  join  transition  place  output  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	20 
    -- CP-element group 59: 	24 
    -- CP-element group 59: 	28 
    -- CP-element group 59: 	32 
    -- CP-element group 59: 	38 
    -- CP-element group 59: 	42 
    -- CP-element group 59: 	46 
    -- CP-element group 59: 	50 
    -- CP-element group 59: 	54 
    -- CP-element group 59: 	58 
    -- CP-element group 59: 	12 
    -- CP-element group 59: 	16 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59: 	61 
    -- CP-element group 59:  members (10) 
      -- CP-element group 59: 	 branch_block_stmt_224/if_stmt_422__entry__
      -- CP-element group 59: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421__exit__
      -- CP-element group 59: 	 branch_block_stmt_224/assign_stmt_227_to_assign_stmt_421/$exit
      -- CP-element group 59: 	 branch_block_stmt_224/if_stmt_422_dead_link/$entry
      -- CP-element group 59: 	 branch_block_stmt_224/if_stmt_422_eval_test/$entry
      -- CP-element group 59: 	 branch_block_stmt_224/if_stmt_422_eval_test/$exit
      -- CP-element group 59: 	 branch_block_stmt_224/if_stmt_422_eval_test/branch_req
      -- CP-element group 59: 	 branch_block_stmt_224/R_cmp229_423_place
      -- CP-element group 59: 	 branch_block_stmt_224/if_stmt_422_if_link/$entry
      -- CP-element group 59: 	 branch_block_stmt_224/if_stmt_422_else_link/$entry
      -- 
    branch_req_1126_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1126_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(59), ack => if_stmt_422_branch_req_0); -- 
    zeropad3D_cp_element_group_59: block -- 
      constant place_capacities: IntegerArray(0 to 11) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1);
      constant place_markings: IntegerArray(0 to 11)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0);
      constant place_delays: IntegerArray(0 to 11) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0);
      constant joinName: string(1 to 29) := "zeropad3D_cp_element_group_59"; 
      signal preds: BooleanArray(1 to 12); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(20) & zeropad3D_CP_676_elements(24) & zeropad3D_CP_676_elements(28) & zeropad3D_CP_676_elements(32) & zeropad3D_CP_676_elements(38) & zeropad3D_CP_676_elements(42) & zeropad3D_CP_676_elements(46) & zeropad3D_CP_676_elements(50) & zeropad3D_CP_676_elements(54) & zeropad3D_CP_676_elements(58) & zeropad3D_CP_676_elements(12) & zeropad3D_CP_676_elements(16);
      gj_zeropad3D_cp_element_group_59 : generic_join generic map(name => joinName, number_of_predecessors => 12, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(59), clk => clk, reset => reset); --
    end block;
    -- CP-element group 60:  merge  transition  place  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	170 
    -- CP-element group 60:  members (18) 
      -- CP-element group 60: 	 branch_block_stmt_224/bbx_xnph_forx_xbody
      -- CP-element group 60: 	 branch_block_stmt_224/assign_stmt_434_to_assign_stmt_447__exit__
      -- CP-element group 60: 	 branch_block_stmt_224/assign_stmt_434_to_assign_stmt_447__entry__
      -- CP-element group 60: 	 branch_block_stmt_224/merge_stmt_428__exit__
      -- CP-element group 60: 	 branch_block_stmt_224/if_stmt_422_if_link/$exit
      -- CP-element group 60: 	 branch_block_stmt_224/if_stmt_422_if_link/if_choice_transition
      -- CP-element group 60: 	 branch_block_stmt_224/entry_bbx_xnph
      -- CP-element group 60: 	 branch_block_stmt_224/assign_stmt_434_to_assign_stmt_447/$entry
      -- CP-element group 60: 	 branch_block_stmt_224/assign_stmt_434_to_assign_stmt_447/$exit
      -- CP-element group 60: 	 branch_block_stmt_224/entry_bbx_xnph_PhiReq/$entry
      -- CP-element group 60: 	 branch_block_stmt_224/entry_bbx_xnph_PhiReq/$exit
      -- CP-element group 60: 	 branch_block_stmt_224/merge_stmt_428_PhiReqMerge
      -- CP-element group 60: 	 branch_block_stmt_224/merge_stmt_428_PhiAck/$entry
      -- CP-element group 60: 	 branch_block_stmt_224/merge_stmt_428_PhiAck/$exit
      -- CP-element group 60: 	 branch_block_stmt_224/merge_stmt_428_PhiAck/dummy
      -- CP-element group 60: 	 branch_block_stmt_224/bbx_xnph_forx_xbody_PhiReq/$entry
      -- CP-element group 60: 	 branch_block_stmt_224/bbx_xnph_forx_xbody_PhiReq/phi_stmt_450/$entry
      -- CP-element group 60: 	 branch_block_stmt_224/bbx_xnph_forx_xbody_PhiReq/phi_stmt_450/phi_stmt_450_sources/$entry
      -- 
    if_choice_transition_1131_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_422_branch_ack_1, ack => zeropad3D_CP_676_elements(60)); -- 
    -- CP-element group 61:  transition  place  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	59 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	176 
    -- CP-element group 61:  members (5) 
      -- CP-element group 61: 	 branch_block_stmt_224/if_stmt_422_else_link/$exit
      -- CP-element group 61: 	 branch_block_stmt_224/if_stmt_422_else_link/else_choice_transition
      -- CP-element group 61: 	 branch_block_stmt_224/entry_forx_xend
      -- CP-element group 61: 	 branch_block_stmt_224/entry_forx_xend_PhiReq/$entry
      -- CP-element group 61: 	 branch_block_stmt_224/entry_forx_xend_PhiReq/$exit
      -- 
    else_choice_transition_1135_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_422_branch_ack_0, ack => zeropad3D_CP_676_elements(61)); -- 
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	175 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	101 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/array_obj_ref_462_final_index_sum_regn_sample_complete
      -- CP-element group 62: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/array_obj_ref_462_final_index_sum_regn_Sample/$exit
      -- CP-element group 62: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/array_obj_ref_462_final_index_sum_regn_Sample/ack
      -- 
    ack_1169_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_462_index_offset_ack_0, ack => zeropad3D_CP_676_elements(62)); -- 
    -- CP-element group 63:  transition  input  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	175 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (11) 
      -- CP-element group 63: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/addr_of_463_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/array_obj_ref_462_root_address_calculated
      -- CP-element group 63: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/array_obj_ref_462_offset_calculated
      -- CP-element group 63: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/array_obj_ref_462_final_index_sum_regn_Update/$exit
      -- CP-element group 63: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/array_obj_ref_462_final_index_sum_regn_Update/ack
      -- CP-element group 63: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/array_obj_ref_462_base_plus_offset/$entry
      -- CP-element group 63: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/array_obj_ref_462_base_plus_offset/$exit
      -- CP-element group 63: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/array_obj_ref_462_base_plus_offset/sum_rename_req
      -- CP-element group 63: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/array_obj_ref_462_base_plus_offset/sum_rename_ack
      -- CP-element group 63: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/addr_of_463_request/$entry
      -- CP-element group 63: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/addr_of_463_request/req
      -- 
    ack_1174_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_462_index_offset_ack_1, ack => zeropad3D_CP_676_elements(63)); -- 
    req_1183_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1183_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(63), ack => addr_of_463_final_reg_req_0); -- 
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/addr_of_463_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/addr_of_463_request/$exit
      -- CP-element group 64: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/addr_of_463_request/ack
      -- 
    ack_1184_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_463_final_reg_ack_0, ack => zeropad3D_CP_676_elements(64)); -- 
    -- CP-element group 65:  fork  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	175 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	98 
    -- CP-element group 65:  members (19) 
      -- CP-element group 65: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/addr_of_463_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/addr_of_463_complete/$exit
      -- CP-element group 65: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/addr_of_463_complete/ack
      -- CP-element group 65: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/ptr_deref_599_base_address_calculated
      -- CP-element group 65: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/ptr_deref_599_word_address_calculated
      -- CP-element group 65: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/ptr_deref_599_root_address_calculated
      -- CP-element group 65: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/ptr_deref_599_base_address_resized
      -- CP-element group 65: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/ptr_deref_599_base_addr_resize/$entry
      -- CP-element group 65: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/ptr_deref_599_base_addr_resize/$exit
      -- CP-element group 65: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/ptr_deref_599_base_addr_resize/base_resize_req
      -- CP-element group 65: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/ptr_deref_599_base_addr_resize/base_resize_ack
      -- CP-element group 65: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/ptr_deref_599_base_plus_offset/$entry
      -- CP-element group 65: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/ptr_deref_599_base_plus_offset/$exit
      -- CP-element group 65: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/ptr_deref_599_base_plus_offset/sum_rename_req
      -- CP-element group 65: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/ptr_deref_599_base_plus_offset/sum_rename_ack
      -- CP-element group 65: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/ptr_deref_599_word_addrgen/$entry
      -- CP-element group 65: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/ptr_deref_599_word_addrgen/$exit
      -- CP-element group 65: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/ptr_deref_599_word_addrgen/root_register_req
      -- CP-element group 65: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/ptr_deref_599_word_addrgen/root_register_ack
      -- 
    ack_1189_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_463_final_reg_ack_1, ack => zeropad3D_CP_676_elements(65)); -- 
    -- CP-element group 66:  transition  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	175 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (6) 
      -- CP-element group 66: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_466_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_466_update_start_
      -- CP-element group 66: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_466_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_466_Sample/ra
      -- CP-element group 66: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_466_Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_466_Update/cr
      -- 
    ra_1198_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_466_inst_ack_0, ack => zeropad3D_CP_676_elements(66)); -- 
    cr_1202_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1202_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(66), ack => RPIPE_zeropad_input_pipe_466_inst_req_1); -- 
    -- CP-element group 67:  fork  transition  input  output  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67: 	70 
    -- CP-element group 67:  members (9) 
      -- CP-element group 67: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_466_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_466_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_466_Update/ca
      -- CP-element group 67: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_470_sample_start_
      -- CP-element group 67: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_470_Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_470_Sample/rr
      -- CP-element group 67: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_479_sample_start_
      -- CP-element group 67: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_479_Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_479_Sample/rr
      -- 
    ca_1203_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_466_inst_ack_1, ack => zeropad3D_CP_676_elements(67)); -- 
    rr_1211_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1211_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(67), ack => type_cast_470_inst_req_0); -- 
    rr_1225_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1225_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(67), ack => RPIPE_zeropad_input_pipe_479_inst_req_0); -- 
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_470_sample_completed_
      -- CP-element group 68: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_470_Sample/$exit
      -- CP-element group 68: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_470_Sample/ra
      -- 
    ra_1212_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_470_inst_ack_0, ack => zeropad3D_CP_676_elements(68)); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	175 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	98 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_470_update_completed_
      -- CP-element group 69: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_470_Update/$exit
      -- CP-element group 69: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_470_Update/ca
      -- 
    ca_1217_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_470_inst_ack_1, ack => zeropad3D_CP_676_elements(69)); -- 
    -- CP-element group 70:  transition  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	67 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70:  members (6) 
      -- CP-element group 70: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_479_sample_completed_
      -- CP-element group 70: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_479_update_start_
      -- CP-element group 70: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_479_Sample/$exit
      -- CP-element group 70: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_479_Sample/ra
      -- CP-element group 70: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_479_Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_479_Update/cr
      -- 
    ra_1226_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_479_inst_ack_0, ack => zeropad3D_CP_676_elements(70)); -- 
    cr_1230_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1230_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(70), ack => RPIPE_zeropad_input_pipe_479_inst_req_1); -- 
    -- CP-element group 71:  fork  transition  input  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	72 
    -- CP-element group 71: 	74 
    -- CP-element group 71:  members (9) 
      -- CP-element group 71: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_479_update_completed_
      -- CP-element group 71: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_479_Update/$exit
      -- CP-element group 71: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_479_Update/ca
      -- CP-element group 71: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_483_sample_start_
      -- CP-element group 71: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_483_Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_483_Sample/rr
      -- CP-element group 71: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_497_sample_start_
      -- CP-element group 71: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_497_Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_497_Sample/rr
      -- 
    ca_1231_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_479_inst_ack_1, ack => zeropad3D_CP_676_elements(71)); -- 
    rr_1239_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1239_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(71), ack => type_cast_483_inst_req_0); -- 
    rr_1253_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1253_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(71), ack => RPIPE_zeropad_input_pipe_497_inst_req_0); -- 
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	71 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_483_sample_completed_
      -- CP-element group 72: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_483_Sample/$exit
      -- CP-element group 72: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_483_Sample/ra
      -- 
    ra_1240_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_483_inst_ack_0, ack => zeropad3D_CP_676_elements(72)); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	175 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	98 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_483_update_completed_
      -- CP-element group 73: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_483_Update/$exit
      -- CP-element group 73: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_483_Update/ca
      -- 
    ca_1245_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_483_inst_ack_1, ack => zeropad3D_CP_676_elements(73)); -- 
    -- CP-element group 74:  transition  input  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	71 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74:  members (6) 
      -- CP-element group 74: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_497_sample_completed_
      -- CP-element group 74: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_497_update_start_
      -- CP-element group 74: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_497_Sample/$exit
      -- CP-element group 74: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_497_Sample/ra
      -- CP-element group 74: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_497_Update/$entry
      -- CP-element group 74: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_497_Update/cr
      -- 
    ra_1254_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_497_inst_ack_0, ack => zeropad3D_CP_676_elements(74)); -- 
    cr_1258_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1258_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(74), ack => RPIPE_zeropad_input_pipe_497_inst_req_1); -- 
    -- CP-element group 75:  fork  transition  input  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	76 
    -- CP-element group 75: 	78 
    -- CP-element group 75:  members (9) 
      -- CP-element group 75: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_497_update_completed_
      -- CP-element group 75: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_497_Update/$exit
      -- CP-element group 75: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_497_Update/ca
      -- CP-element group 75: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_501_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_501_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_501_Sample/rr
      -- CP-element group 75: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_515_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_515_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_515_Sample/rr
      -- 
    ca_1259_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_497_inst_ack_1, ack => zeropad3D_CP_676_elements(75)); -- 
    rr_1267_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1267_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(75), ack => type_cast_501_inst_req_0); -- 
    rr_1281_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1281_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(75), ack => RPIPE_zeropad_input_pipe_515_inst_req_0); -- 
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	75 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_501_sample_completed_
      -- CP-element group 76: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_501_Sample/$exit
      -- CP-element group 76: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_501_Sample/ra
      -- 
    ra_1268_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_501_inst_ack_0, ack => zeropad3D_CP_676_elements(76)); -- 
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	175 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	98 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_501_update_completed_
      -- CP-element group 77: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_501_Update/$exit
      -- CP-element group 77: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_501_Update/ca
      -- 
    ca_1273_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_501_inst_ack_1, ack => zeropad3D_CP_676_elements(77)); -- 
    -- CP-element group 78:  transition  input  output  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	75 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78:  members (6) 
      -- CP-element group 78: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_515_sample_completed_
      -- CP-element group 78: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_515_update_start_
      -- CP-element group 78: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_515_Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_515_Sample/ra
      -- CP-element group 78: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_515_Update/$entry
      -- CP-element group 78: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_515_Update/cr
      -- 
    ra_1282_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_515_inst_ack_0, ack => zeropad3D_CP_676_elements(78)); -- 
    cr_1286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(78), ack => RPIPE_zeropad_input_pipe_515_inst_req_1); -- 
    -- CP-element group 79:  fork  transition  input  output  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79: 	82 
    -- CP-element group 79:  members (9) 
      -- CP-element group 79: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_515_update_completed_
      -- CP-element group 79: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_515_Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_515_Update/ca
      -- CP-element group 79: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_519_sample_start_
      -- CP-element group 79: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_519_Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_519_Sample/rr
      -- CP-element group 79: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_533_sample_start_
      -- CP-element group 79: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_533_Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_533_Sample/rr
      -- 
    ca_1287_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_515_inst_ack_1, ack => zeropad3D_CP_676_elements(79)); -- 
    rr_1295_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1295_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(79), ack => type_cast_519_inst_req_0); -- 
    rr_1309_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1309_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(79), ack => RPIPE_zeropad_input_pipe_533_inst_req_0); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_519_sample_completed_
      -- CP-element group 80: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_519_Sample/$exit
      -- CP-element group 80: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_519_Sample/ra
      -- 
    ra_1296_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_519_inst_ack_0, ack => zeropad3D_CP_676_elements(80)); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	175 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	98 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_519_update_completed_
      -- CP-element group 81: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_519_Update/$exit
      -- CP-element group 81: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_519_Update/ca
      -- 
    ca_1301_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_519_inst_ack_1, ack => zeropad3D_CP_676_elements(81)); -- 
    -- CP-element group 82:  transition  input  output  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	79 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (6) 
      -- CP-element group 82: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_533_sample_completed_
      -- CP-element group 82: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_533_update_start_
      -- CP-element group 82: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_533_Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_533_Sample/ra
      -- CP-element group 82: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_533_Update/$entry
      -- CP-element group 82: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_533_Update/cr
      -- 
    ra_1310_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_533_inst_ack_0, ack => zeropad3D_CP_676_elements(82)); -- 
    cr_1314_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1314_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(82), ack => RPIPE_zeropad_input_pipe_533_inst_req_1); -- 
    -- CP-element group 83:  fork  transition  input  output  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83: 	86 
    -- CP-element group 83:  members (9) 
      -- CP-element group 83: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_533_update_completed_
      -- CP-element group 83: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_533_Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_533_Update/ca
      -- CP-element group 83: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_537_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_537_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_537_Sample/rr
      -- CP-element group 83: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_551_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_551_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_551_Sample/rr
      -- 
    ca_1315_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_533_inst_ack_1, ack => zeropad3D_CP_676_elements(83)); -- 
    rr_1323_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1323_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(83), ack => type_cast_537_inst_req_0); -- 
    rr_1337_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1337_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(83), ack => RPIPE_zeropad_input_pipe_551_inst_req_0); -- 
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_537_sample_completed_
      -- CP-element group 84: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_537_Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_537_Sample/ra
      -- 
    ra_1324_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_537_inst_ack_0, ack => zeropad3D_CP_676_elements(84)); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	175 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	98 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_537_update_completed_
      -- CP-element group 85: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_537_Update/$exit
      -- CP-element group 85: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_537_Update/ca
      -- 
    ca_1329_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_537_inst_ack_1, ack => zeropad3D_CP_676_elements(85)); -- 
    -- CP-element group 86:  transition  input  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	83 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (6) 
      -- CP-element group 86: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_551_sample_completed_
      -- CP-element group 86: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_551_update_start_
      -- CP-element group 86: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_551_Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_551_Sample/ra
      -- CP-element group 86: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_551_Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_551_Update/cr
      -- 
    ra_1338_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_551_inst_ack_0, ack => zeropad3D_CP_676_elements(86)); -- 
    cr_1342_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1342_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(86), ack => RPIPE_zeropad_input_pipe_551_inst_req_1); -- 
    -- CP-element group 87:  fork  transition  input  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87: 	90 
    -- CP-element group 87:  members (9) 
      -- CP-element group 87: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_551_update_completed_
      -- CP-element group 87: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_551_Update/$exit
      -- CP-element group 87: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_551_Update/ca
      -- CP-element group 87: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_555_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_555_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_555_Sample/rr
      -- CP-element group 87: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_569_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_569_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_569_Sample/rr
      -- 
    ca_1343_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_551_inst_ack_1, ack => zeropad3D_CP_676_elements(87)); -- 
    rr_1351_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1351_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(87), ack => type_cast_555_inst_req_0); -- 
    rr_1365_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1365_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(87), ack => RPIPE_zeropad_input_pipe_569_inst_req_0); -- 
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_555_sample_completed_
      -- CP-element group 88: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_555_Sample/$exit
      -- CP-element group 88: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_555_Sample/ra
      -- 
    ra_1352_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_555_inst_ack_0, ack => zeropad3D_CP_676_elements(88)); -- 
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	175 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	98 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_555_update_completed_
      -- CP-element group 89: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_555_Update/$exit
      -- CP-element group 89: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_555_Update/ca
      -- 
    ca_1357_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_555_inst_ack_1, ack => zeropad3D_CP_676_elements(89)); -- 
    -- CP-element group 90:  transition  input  output  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	87 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (6) 
      -- CP-element group 90: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_569_sample_completed_
      -- CP-element group 90: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_569_update_start_
      -- CP-element group 90: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_569_Sample/$exit
      -- CP-element group 90: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_569_Sample/ra
      -- CP-element group 90: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_569_Update/$entry
      -- CP-element group 90: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_569_Update/cr
      -- 
    ra_1366_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_569_inst_ack_0, ack => zeropad3D_CP_676_elements(90)); -- 
    cr_1370_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1370_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(90), ack => RPIPE_zeropad_input_pipe_569_inst_req_1); -- 
    -- CP-element group 91:  fork  transition  input  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91: 	94 
    -- CP-element group 91:  members (9) 
      -- CP-element group 91: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_569_update_completed_
      -- CP-element group 91: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_569_Update/$exit
      -- CP-element group 91: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_569_Update/ca
      -- CP-element group 91: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_573_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_573_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_573_Sample/rr
      -- CP-element group 91: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_587_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_587_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_587_Sample/rr
      -- 
    ca_1371_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_569_inst_ack_1, ack => zeropad3D_CP_676_elements(91)); -- 
    rr_1379_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1379_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(91), ack => type_cast_573_inst_req_0); -- 
    rr_1393_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1393_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(91), ack => RPIPE_zeropad_input_pipe_587_inst_req_0); -- 
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92:  members (3) 
      -- CP-element group 92: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_573_sample_completed_
      -- CP-element group 92: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_573_Sample/$exit
      -- CP-element group 92: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_573_Sample/ra
      -- 
    ra_1380_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_573_inst_ack_0, ack => zeropad3D_CP_676_elements(92)); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	175 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	98 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_573_update_completed_
      -- CP-element group 93: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_573_Update/$exit
      -- CP-element group 93: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_573_Update/ca
      -- 
    ca_1385_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_573_inst_ack_1, ack => zeropad3D_CP_676_elements(93)); -- 
    -- CP-element group 94:  transition  input  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	91 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94:  members (6) 
      -- CP-element group 94: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_587_sample_completed_
      -- CP-element group 94: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_587_update_start_
      -- CP-element group 94: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_587_Sample/$exit
      -- CP-element group 94: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_587_Sample/ra
      -- CP-element group 94: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_587_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_587_Update/cr
      -- 
    ra_1394_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_587_inst_ack_0, ack => zeropad3D_CP_676_elements(94)); -- 
    cr_1398_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1398_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(94), ack => RPIPE_zeropad_input_pipe_587_inst_req_1); -- 
    -- CP-element group 95:  transition  input  output  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95:  members (6) 
      -- CP-element group 95: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_587_update_completed_
      -- CP-element group 95: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_587_Update/$exit
      -- CP-element group 95: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_587_Update/ca
      -- CP-element group 95: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_591_sample_start_
      -- CP-element group 95: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_591_Sample/$entry
      -- CP-element group 95: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_591_Sample/rr
      -- 
    ca_1399_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_zeropad_input_pipe_587_inst_ack_1, ack => zeropad3D_CP_676_elements(95)); -- 
    rr_1407_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1407_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(95), ack => type_cast_591_inst_req_0); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_591_sample_completed_
      -- CP-element group 96: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_591_Sample/$exit
      -- CP-element group 96: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_591_Sample/ra
      -- 
    ra_1408_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_591_inst_ack_0, ack => zeropad3D_CP_676_elements(96)); -- 
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	175 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_591_update_completed_
      -- CP-element group 97: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_591_Update/$exit
      -- CP-element group 97: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_591_Update/ca
      -- 
    ca_1413_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_591_inst_ack_1, ack => zeropad3D_CP_676_elements(97)); -- 
    -- CP-element group 98:  join  transition  output  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	65 
    -- CP-element group 98: 	69 
    -- CP-element group 98: 	73 
    -- CP-element group 98: 	77 
    -- CP-element group 98: 	81 
    -- CP-element group 98: 	85 
    -- CP-element group 98: 	89 
    -- CP-element group 98: 	93 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (9) 
      -- CP-element group 98: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/ptr_deref_599_sample_start_
      -- CP-element group 98: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/ptr_deref_599_Sample/$entry
      -- CP-element group 98: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/ptr_deref_599_Sample/ptr_deref_599_Split/$entry
      -- CP-element group 98: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/ptr_deref_599_Sample/ptr_deref_599_Split/$exit
      -- CP-element group 98: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/ptr_deref_599_Sample/ptr_deref_599_Split/split_req
      -- CP-element group 98: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/ptr_deref_599_Sample/ptr_deref_599_Split/split_ack
      -- CP-element group 98: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/ptr_deref_599_Sample/word_access_start/$entry
      -- CP-element group 98: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/ptr_deref_599_Sample/word_access_start/word_0/$entry
      -- CP-element group 98: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/ptr_deref_599_Sample/word_access_start/word_0/rr
      -- 
    rr_1451_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1451_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(98), ack => ptr_deref_599_store_0_req_0); -- 
    zeropad3D_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 29) := "zeropad3D_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(65) & zeropad3D_CP_676_elements(69) & zeropad3D_CP_676_elements(73) & zeropad3D_CP_676_elements(77) & zeropad3D_CP_676_elements(81) & zeropad3D_CP_676_elements(85) & zeropad3D_CP_676_elements(89) & zeropad3D_CP_676_elements(93) & zeropad3D_CP_676_elements(97);
      gj_zeropad3D_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99:  members (5) 
      -- CP-element group 99: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/ptr_deref_599_sample_completed_
      -- CP-element group 99: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/ptr_deref_599_Sample/$exit
      -- CP-element group 99: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/ptr_deref_599_Sample/word_access_start/$exit
      -- CP-element group 99: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/ptr_deref_599_Sample/word_access_start/word_0/$exit
      -- CP-element group 99: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/ptr_deref_599_Sample/word_access_start/word_0/ra
      -- 
    ra_1452_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_599_store_0_ack_0, ack => zeropad3D_CP_676_elements(99)); -- 
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	175 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	101 
    -- CP-element group 100:  members (5) 
      -- CP-element group 100: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/ptr_deref_599_update_completed_
      -- CP-element group 100: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/ptr_deref_599_Update/$exit
      -- CP-element group 100: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/ptr_deref_599_Update/word_access_complete/$exit
      -- CP-element group 100: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/ptr_deref_599_Update/word_access_complete/word_0/$exit
      -- CP-element group 100: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/ptr_deref_599_Update/word_access_complete/word_0/ca
      -- 
    ca_1463_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_599_store_0_ack_1, ack => zeropad3D_CP_676_elements(100)); -- 
    -- CP-element group 101:  branch  join  transition  place  output  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	62 
    -- CP-element group 101: 	100 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	102 
    -- CP-element group 101: 	103 
    -- CP-element group 101:  members (10) 
      -- CP-element group 101: 	 branch_block_stmt_224/if_stmt_613__entry__
      -- CP-element group 101: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612__exit__
      -- CP-element group 101: 	 branch_block_stmt_224/if_stmt_613_else_link/$entry
      -- CP-element group 101: 	 branch_block_stmt_224/R_exitcond3_614_place
      -- CP-element group 101: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/$exit
      -- CP-element group 101: 	 branch_block_stmt_224/if_stmt_613_if_link/$entry
      -- CP-element group 101: 	 branch_block_stmt_224/if_stmt_613_eval_test/branch_req
      -- CP-element group 101: 	 branch_block_stmt_224/if_stmt_613_eval_test/$exit
      -- CP-element group 101: 	 branch_block_stmt_224/if_stmt_613_dead_link/$entry
      -- CP-element group 101: 	 branch_block_stmt_224/if_stmt_613_eval_test/$entry
      -- 
    branch_req_1471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(101), ack => if_stmt_613_branch_req_0); -- 
    zeropad3D_cp_element_group_101: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_101"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(62) & zeropad3D_CP_676_elements(100);
      gj_zeropad3D_cp_element_group_101 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(101), clk => clk, reset => reset); --
    end block;
    -- CP-element group 102:  merge  transition  place  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	101 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	176 
    -- CP-element group 102:  members (13) 
      -- CP-element group 102: 	 branch_block_stmt_224/forx_xendx_xloopexit_forx_xend
      -- CP-element group 102: 	 branch_block_stmt_224/merge_stmt_619__exit__
      -- CP-element group 102: 	 branch_block_stmt_224/forx_xbody_forx_xendx_xloopexit
      -- CP-element group 102: 	 branch_block_stmt_224/if_stmt_613_if_link/if_choice_transition
      -- CP-element group 102: 	 branch_block_stmt_224/if_stmt_613_if_link/$exit
      -- CP-element group 102: 	 branch_block_stmt_224/forx_xbody_forx_xendx_xloopexit_PhiReq/$entry
      -- CP-element group 102: 	 branch_block_stmt_224/forx_xbody_forx_xendx_xloopexit_PhiReq/$exit
      -- CP-element group 102: 	 branch_block_stmt_224/merge_stmt_619_PhiReqMerge
      -- CP-element group 102: 	 branch_block_stmt_224/merge_stmt_619_PhiAck/$entry
      -- CP-element group 102: 	 branch_block_stmt_224/merge_stmt_619_PhiAck/$exit
      -- CP-element group 102: 	 branch_block_stmt_224/merge_stmt_619_PhiAck/dummy
      -- CP-element group 102: 	 branch_block_stmt_224/forx_xendx_xloopexit_forx_xend_PhiReq/$entry
      -- CP-element group 102: 	 branch_block_stmt_224/forx_xendx_xloopexit_forx_xend_PhiReq/$exit
      -- 
    if_choice_transition_1476_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_613_branch_ack_1, ack => zeropad3D_CP_676_elements(102)); -- 
    -- CP-element group 103:  fork  transition  place  input  output  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	101 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	171 
    -- CP-element group 103: 	172 
    -- CP-element group 103:  members (12) 
      -- CP-element group 103: 	 branch_block_stmt_224/if_stmt_613_else_link/$exit
      -- CP-element group 103: 	 branch_block_stmt_224/if_stmt_613_else_link/else_choice_transition
      -- CP-element group 103: 	 branch_block_stmt_224/forx_xbody_forx_xbody
      -- CP-element group 103: 	 branch_block_stmt_224/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 103: 	 branch_block_stmt_224/forx_xbody_forx_xbody_PhiReq/phi_stmt_450/$entry
      -- CP-element group 103: 	 branch_block_stmt_224/forx_xbody_forx_xbody_PhiReq/phi_stmt_450/phi_stmt_450_sources/$entry
      -- CP-element group 103: 	 branch_block_stmt_224/forx_xbody_forx_xbody_PhiReq/phi_stmt_450/phi_stmt_450_sources/type_cast_456/$entry
      -- CP-element group 103: 	 branch_block_stmt_224/forx_xbody_forx_xbody_PhiReq/phi_stmt_450/phi_stmt_450_sources/type_cast_456/SplitProtocol/$entry
      -- CP-element group 103: 	 branch_block_stmt_224/forx_xbody_forx_xbody_PhiReq/phi_stmt_450/phi_stmt_450_sources/type_cast_456/SplitProtocol/Sample/$entry
      -- CP-element group 103: 	 branch_block_stmt_224/forx_xbody_forx_xbody_PhiReq/phi_stmt_450/phi_stmt_450_sources/type_cast_456/SplitProtocol/Sample/rr
      -- CP-element group 103: 	 branch_block_stmt_224/forx_xbody_forx_xbody_PhiReq/phi_stmt_450/phi_stmt_450_sources/type_cast_456/SplitProtocol/Update/$entry
      -- CP-element group 103: 	 branch_block_stmt_224/forx_xbody_forx_xbody_PhiReq/phi_stmt_450/phi_stmt_450_sources/type_cast_456/SplitProtocol/Update/cr
      -- 
    else_choice_transition_1480_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_613_branch_ack_0, ack => zeropad3D_CP_676_elements(103)); -- 
    rr_1939_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1939_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(103), ack => type_cast_456_inst_req_0); -- 
    cr_1944_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1944_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(103), ack => type_cast_456_inst_req_1); -- 
    -- CP-element group 104:  transition  input  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	176 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (3) 
      -- CP-element group 104: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/call_stmt_624_sample_completed_
      -- CP-element group 104: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/call_stmt_624_Sample/cra
      -- CP-element group 104: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/call_stmt_624_Sample/$exit
      -- 
    cra_1494_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_624_call_ack_0, ack => zeropad3D_CP_676_elements(104)); -- 
    -- CP-element group 105:  transition  input  output  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	176 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	106 
    -- CP-element group 105:  members (6) 
      -- CP-element group 105: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/type_cast_628_sample_start_
      -- CP-element group 105: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/call_stmt_624_Update/$exit
      -- CP-element group 105: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/call_stmt_624_update_completed_
      -- CP-element group 105: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/call_stmt_624_Update/cca
      -- CP-element group 105: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/type_cast_628_Sample/rr
      -- CP-element group 105: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/type_cast_628_Sample/$entry
      -- 
    cca_1499_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_624_call_ack_1, ack => zeropad3D_CP_676_elements(105)); -- 
    rr_1507_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1507_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(105), ack => type_cast_628_inst_req_0); -- 
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	105 
    -- CP-element group 106: successors 
    -- CP-element group 106:  members (3) 
      -- CP-element group 106: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/type_cast_628_sample_completed_
      -- CP-element group 106: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/type_cast_628_Sample/ra
      -- CP-element group 106: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/type_cast_628_Sample/$exit
      -- 
    ra_1508_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_628_inst_ack_0, ack => zeropad3D_CP_676_elements(106)); -- 
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	176 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	124 
    -- CP-element group 107:  members (3) 
      -- CP-element group 107: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/type_cast_628_Update/ca
      -- CP-element group 107: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/type_cast_628_Update/$exit
      -- CP-element group 107: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/type_cast_628_update_completed_
      -- 
    ca_1513_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_628_inst_ack_1, ack => zeropad3D_CP_676_elements(107)); -- 
    -- CP-element group 108:  transition  input  output  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	176 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	109 
    -- CP-element group 108:  members (6) 
      -- CP-element group 108: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_630_Update/$entry
      -- CP-element group 108: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_630_Sample/ack
      -- CP-element group 108: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_630_Sample/$exit
      -- CP-element group 108: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_630_Update/req
      -- CP-element group 108: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_630_sample_completed_
      -- CP-element group 108: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_630_update_start_
      -- 
    ack_1522_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_starting_630_inst_ack_0, ack => zeropad3D_CP_676_elements(108)); -- 
    req_1526_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1526_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(108), ack => WPIPE_Block0_starting_630_inst_req_1); -- 
    -- CP-element group 109:  transition  input  output  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	108 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	110 
    -- CP-element group 109:  members (6) 
      -- CP-element group 109: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_630_Update/$exit
      -- CP-element group 109: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_633_sample_start_
      -- CP-element group 109: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_630_update_completed_
      -- CP-element group 109: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_630_Update/ack
      -- CP-element group 109: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_633_Sample/req
      -- CP-element group 109: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_633_Sample/$entry
      -- 
    ack_1527_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_starting_630_inst_ack_1, ack => zeropad3D_CP_676_elements(109)); -- 
    req_1535_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1535_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(109), ack => WPIPE_Block0_starting_633_inst_req_0); -- 
    -- CP-element group 110:  transition  input  output  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	109 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (6) 
      -- CP-element group 110: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_633_sample_completed_
      -- CP-element group 110: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_633_Update/req
      -- CP-element group 110: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_633_Update/$entry
      -- CP-element group 110: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_633_Sample/ack
      -- CP-element group 110: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_633_Sample/$exit
      -- CP-element group 110: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_633_update_start_
      -- 
    ack_1536_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_starting_633_inst_ack_0, ack => zeropad3D_CP_676_elements(110)); -- 
    req_1540_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1540_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(110), ack => WPIPE_Block0_starting_633_inst_req_1); -- 
    -- CP-element group 111:  transition  input  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111:  members (6) 
      -- CP-element group 111: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_636_Sample/req
      -- CP-element group 111: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_636_Sample/$entry
      -- CP-element group 111: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_636_sample_start_
      -- CP-element group 111: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_633_Update/ack
      -- CP-element group 111: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_633_Update/$exit
      -- CP-element group 111: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_633_update_completed_
      -- 
    ack_1541_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_starting_633_inst_ack_1, ack => zeropad3D_CP_676_elements(111)); -- 
    req_1549_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1549_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(111), ack => WPIPE_Block0_starting_636_inst_req_0); -- 
    -- CP-element group 112:  transition  input  output  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	113 
    -- CP-element group 112:  members (6) 
      -- CP-element group 112: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_636_Update/req
      -- CP-element group 112: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_636_Update/$entry
      -- CP-element group 112: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_636_Sample/ack
      -- CP-element group 112: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_636_Sample/$exit
      -- CP-element group 112: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_636_update_start_
      -- CP-element group 112: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_636_sample_completed_
      -- 
    ack_1550_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_starting_636_inst_ack_0, ack => zeropad3D_CP_676_elements(112)); -- 
    req_1554_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1554_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(112), ack => WPIPE_Block0_starting_636_inst_req_1); -- 
    -- CP-element group 113:  transition  input  output  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	112 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	114 
    -- CP-element group 113:  members (6) 
      -- CP-element group 113: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_639_Sample/$entry
      -- CP-element group 113: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_639_Sample/req
      -- CP-element group 113: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_639_sample_start_
      -- CP-element group 113: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_636_Update/ack
      -- CP-element group 113: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_636_Update/$exit
      -- CP-element group 113: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_636_update_completed_
      -- 
    ack_1555_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_starting_636_inst_ack_1, ack => zeropad3D_CP_676_elements(113)); -- 
    req_1563_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1563_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(113), ack => WPIPE_Block0_starting_639_inst_req_0); -- 
    -- CP-element group 114:  transition  input  output  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	113 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (6) 
      -- CP-element group 114: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_639_sample_completed_
      -- CP-element group 114: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_639_Sample/ack
      -- CP-element group 114: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_639_Sample/$exit
      -- CP-element group 114: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_639_Update/$entry
      -- CP-element group 114: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_639_Update/req
      -- CP-element group 114: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_639_update_start_
      -- 
    ack_1564_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_starting_639_inst_ack_0, ack => zeropad3D_CP_676_elements(114)); -- 
    req_1568_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1568_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(114), ack => WPIPE_Block0_starting_639_inst_req_1); -- 
    -- CP-element group 115:  transition  input  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	116 
    -- CP-element group 115:  members (6) 
      -- CP-element group 115: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_642_Sample/req
      -- CP-element group 115: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_639_Update/$exit
      -- CP-element group 115: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_642_Sample/$entry
      -- CP-element group 115: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_642_sample_start_
      -- CP-element group 115: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_639_update_completed_
      -- CP-element group 115: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_639_Update/ack
      -- 
    ack_1569_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_starting_639_inst_ack_1, ack => zeropad3D_CP_676_elements(115)); -- 
    req_1577_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1577_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(115), ack => WPIPE_Block0_starting_642_inst_req_0); -- 
    -- CP-element group 116:  transition  input  output  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	115 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	117 
    -- CP-element group 116:  members (6) 
      -- CP-element group 116: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_642_update_start_
      -- CP-element group 116: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_642_Update/req
      -- CP-element group 116: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_642_Sample/$exit
      -- CP-element group 116: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_642_Sample/ack
      -- CP-element group 116: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_642_Update/$entry
      -- CP-element group 116: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_642_sample_completed_
      -- 
    ack_1578_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_starting_642_inst_ack_0, ack => zeropad3D_CP_676_elements(116)); -- 
    req_1582_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1582_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(116), ack => WPIPE_Block0_starting_642_inst_req_1); -- 
    -- CP-element group 117:  transition  input  output  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	116 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	118 
    -- CP-element group 117:  members (6) 
      -- CP-element group 117: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_642_update_completed_
      -- CP-element group 117: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_642_Update/ack
      -- CP-element group 117: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_645_sample_start_
      -- CP-element group 117: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_645_Sample/req
      -- CP-element group 117: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_645_Sample/$entry
      -- CP-element group 117: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_642_Update/$exit
      -- 
    ack_1583_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_starting_642_inst_ack_1, ack => zeropad3D_CP_676_elements(117)); -- 
    req_1591_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1591_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(117), ack => WPIPE_Block0_starting_645_inst_req_0); -- 
    -- CP-element group 118:  transition  input  output  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	117 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	119 
    -- CP-element group 118:  members (6) 
      -- CP-element group 118: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_645_Sample/$exit
      -- CP-element group 118: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_645_update_start_
      -- CP-element group 118: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_645_Update/req
      -- CP-element group 118: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_645_Sample/ack
      -- CP-element group 118: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_645_sample_completed_
      -- CP-element group 118: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_645_Update/$entry
      -- 
    ack_1592_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_starting_645_inst_ack_0, ack => zeropad3D_CP_676_elements(118)); -- 
    req_1596_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1596_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(118), ack => WPIPE_Block0_starting_645_inst_req_1); -- 
    -- CP-element group 119:  transition  input  output  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	118 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	120 
    -- CP-element group 119:  members (6) 
      -- CP-element group 119: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_645_Update/$exit
      -- CP-element group 119: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_645_Update/ack
      -- CP-element group 119: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_648_sample_start_
      -- CP-element group 119: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_648_Sample/$entry
      -- CP-element group 119: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_645_update_completed_
      -- CP-element group 119: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_648_Sample/req
      -- 
    ack_1597_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_starting_645_inst_ack_1, ack => zeropad3D_CP_676_elements(119)); -- 
    req_1605_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1605_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(119), ack => WPIPE_Block0_starting_648_inst_req_0); -- 
    -- CP-element group 120:  transition  input  output  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	119 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120:  members (6) 
      -- CP-element group 120: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_648_sample_completed_
      -- CP-element group 120: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_648_update_start_
      -- CP-element group 120: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_648_Sample/$exit
      -- CP-element group 120: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_648_Update/req
      -- CP-element group 120: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_648_Update/$entry
      -- CP-element group 120: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_648_Sample/ack
      -- 
    ack_1606_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_starting_648_inst_ack_0, ack => zeropad3D_CP_676_elements(120)); -- 
    req_1610_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1610_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(120), ack => WPIPE_Block0_starting_648_inst_req_1); -- 
    -- CP-element group 121:  transition  input  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	124 
    -- CP-element group 121:  members (3) 
      -- CP-element group 121: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_648_update_completed_
      -- CP-element group 121: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_648_Update/ack
      -- CP-element group 121: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_648_Update/$exit
      -- 
    ack_1611_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_starting_648_inst_ack_1, ack => zeropad3D_CP_676_elements(121)); -- 
    -- CP-element group 122:  transition  input  output  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	176 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	123 
    -- CP-element group 122:  members (6) 
      -- CP-element group 122: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/RPIPE_Block0_complete_652_Update/cr
      -- CP-element group 122: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/RPIPE_Block0_complete_652_Update/$entry
      -- CP-element group 122: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/RPIPE_Block0_complete_652_Sample/ra
      -- CP-element group 122: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/RPIPE_Block0_complete_652_Sample/$exit
      -- CP-element group 122: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/RPIPE_Block0_complete_652_update_start_
      -- CP-element group 122: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/RPIPE_Block0_complete_652_sample_completed_
      -- 
    ra_1620_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_complete_652_inst_ack_0, ack => zeropad3D_CP_676_elements(122)); -- 
    cr_1624_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1624_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(122), ack => RPIPE_Block0_complete_652_inst_req_1); -- 
    -- CP-element group 123:  transition  input  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	122 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	124 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/RPIPE_Block0_complete_652_Update/ca
      -- CP-element group 123: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/RPIPE_Block0_complete_652_Update/$exit
      -- CP-element group 123: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/RPIPE_Block0_complete_652_update_completed_
      -- 
    ca_1625_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_complete_652_inst_ack_1, ack => zeropad3D_CP_676_elements(123)); -- 
    -- CP-element group 124:  join  fork  transition  place  output  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	107 
    -- CP-element group 124: 	121 
    -- CP-element group 124: 	123 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	125 
    -- CP-element group 124: 	126 
    -- CP-element group 124: 	128 
    -- CP-element group 124: 	130 
    -- CP-element group 124: 	132 
    -- CP-element group 124: 	134 
    -- CP-element group 124: 	136 
    -- CP-element group 124: 	138 
    -- CP-element group 124: 	140 
    -- CP-element group 124: 	142 
    -- CP-element group 124: 	144 
    -- CP-element group 124:  members (37) 
      -- CP-element group 124: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653__exit__
      -- CP-element group 124: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764__entry__
      -- CP-element group 124: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_679_Update/cr
      -- CP-element group 124: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/$exit
      -- CP-element group 124: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_689_Update/$entry
      -- CP-element group 124: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_689_update_start_
      -- CP-element group 124: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_729_Update/$entry
      -- CP-element group 124: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_719_update_start_
      -- CP-element group 124: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_729_Update/cr
      -- CP-element group 124: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_679_update_start_
      -- CP-element group 124: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_709_Update/cr
      -- CP-element group 124: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_709_Update/$entry
      -- CP-element group 124: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_669_Update/cr
      -- CP-element group 124: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_669_Update/$entry
      -- CP-element group 124: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_679_Update/$entry
      -- CP-element group 124: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_729_update_start_
      -- CP-element group 124: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_669_update_start_
      -- CP-element group 124: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_709_update_start_
      -- CP-element group 124: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_660_Update/cr
      -- CP-element group 124: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_739_Update/cr
      -- CP-element group 124: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_660_Update/$entry
      -- CP-element group 124: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_739_Update/$entry
      -- CP-element group 124: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_689_Update/cr
      -- CP-element group 124: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_719_Update/cr
      -- CP-element group 124: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_660_update_start_
      -- CP-element group 124: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_719_Update/$entry
      -- CP-element group 124: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/call_stmt_656_Update/ccr
      -- CP-element group 124: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_699_Update/cr
      -- CP-element group 124: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_699_Update/$entry
      -- CP-element group 124: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/call_stmt_656_Update/$entry
      -- CP-element group 124: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/call_stmt_656_Sample/crr
      -- CP-element group 124: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/call_stmt_656_Sample/$entry
      -- CP-element group 124: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/call_stmt_656_update_start_
      -- CP-element group 124: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/call_stmt_656_sample_start_
      -- CP-element group 124: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/$entry
      -- CP-element group 124: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_739_update_start_
      -- CP-element group 124: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_699_update_start_
      -- 
    cr_1683_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1683_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(124), ack => type_cast_679_inst_req_1); -- 
    cr_1753_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1753_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(124), ack => type_cast_729_inst_req_1); -- 
    cr_1725_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1725_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(124), ack => type_cast_709_inst_req_1); -- 
    cr_1669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(124), ack => type_cast_669_inst_req_1); -- 
    cr_1655_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1655_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(124), ack => type_cast_660_inst_req_1); -- 
    cr_1767_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1767_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(124), ack => type_cast_739_inst_req_1); -- 
    cr_1697_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1697_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(124), ack => type_cast_689_inst_req_1); -- 
    cr_1739_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1739_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(124), ack => type_cast_719_inst_req_1); -- 
    ccr_1641_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1641_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(124), ack => call_stmt_656_call_req_1); -- 
    cr_1711_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1711_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(124), ack => type_cast_699_inst_req_1); -- 
    crr_1636_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1636_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(124), ack => call_stmt_656_call_req_0); -- 
    zeropad3D_cp_element_group_124: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_124"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(107) & zeropad3D_CP_676_elements(121) & zeropad3D_CP_676_elements(123);
      gj_zeropad3D_cp_element_group_124 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(124), clk => clk, reset => reset); --
    end block;
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	124 
    -- CP-element group 125: successors 
    -- CP-element group 125:  members (3) 
      -- CP-element group 125: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/call_stmt_656_Sample/cra
      -- CP-element group 125: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/call_stmt_656_Sample/$exit
      -- CP-element group 125: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/call_stmt_656_sample_completed_
      -- 
    cra_1637_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_656_call_ack_0, ack => zeropad3D_CP_676_elements(125)); -- 
    -- CP-element group 126:  transition  input  output  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	124 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126:  members (6) 
      -- CP-element group 126: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_660_Sample/rr
      -- CP-element group 126: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_660_Sample/$entry
      -- CP-element group 126: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_660_sample_start_
      -- CP-element group 126: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/call_stmt_656_Update/cca
      -- CP-element group 126: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/call_stmt_656_Update/$exit
      -- CP-element group 126: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/call_stmt_656_update_completed_
      -- 
    cca_1642_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_656_call_ack_1, ack => zeropad3D_CP_676_elements(126)); -- 
    rr_1650_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1650_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(126), ack => type_cast_660_inst_req_0); -- 
    -- CP-element group 127:  transition  input  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_660_Sample/ra
      -- CP-element group 127: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_660_Sample/$exit
      -- CP-element group 127: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_660_sample_completed_
      -- 
    ra_1651_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_660_inst_ack_0, ack => zeropad3D_CP_676_elements(127)); -- 
    -- CP-element group 128:  fork  transition  input  output  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	124 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	129 
    -- CP-element group 128: 	131 
    -- CP-element group 128: 	133 
    -- CP-element group 128: 	135 
    -- CP-element group 128: 	137 
    -- CP-element group 128: 	139 
    -- CP-element group 128: 	141 
    -- CP-element group 128: 	143 
    -- CP-element group 128:  members (27) 
      -- CP-element group 128: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_679_sample_start_
      -- CP-element group 128: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_719_sample_start_
      -- CP-element group 128: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_679_Sample/rr
      -- CP-element group 128: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_689_Sample/$entry
      -- CP-element group 128: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_709_Sample/rr
      -- CP-element group 128: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_689_sample_start_
      -- CP-element group 128: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_729_Sample/rr
      -- CP-element group 128: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_729_Sample/$entry
      -- CP-element group 128: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_699_sample_start_
      -- CP-element group 128: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_679_Sample/$entry
      -- CP-element group 128: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_689_Sample/rr
      -- CP-element group 128: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_669_Sample/rr
      -- CP-element group 128: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_669_Sample/$entry
      -- CP-element group 128: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_709_Sample/$entry
      -- CP-element group 128: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_729_sample_start_
      -- CP-element group 128: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_669_sample_start_
      -- CP-element group 128: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_660_Update/ca
      -- CP-element group 128: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_660_Update/$exit
      -- CP-element group 128: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_709_sample_start_
      -- CP-element group 128: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_660_update_completed_
      -- CP-element group 128: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_739_Sample/rr
      -- CP-element group 128: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_739_Sample/$entry
      -- CP-element group 128: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_699_Sample/rr
      -- CP-element group 128: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_719_Sample/rr
      -- CP-element group 128: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_699_Sample/$entry
      -- CP-element group 128: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_719_Sample/$entry
      -- CP-element group 128: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_739_sample_start_
      -- 
    ca_1656_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_660_inst_ack_1, ack => zeropad3D_CP_676_elements(128)); -- 
    rr_1664_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1664_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(128), ack => type_cast_669_inst_req_0); -- 
    rr_1678_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1678_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(128), ack => type_cast_679_inst_req_0); -- 
    rr_1692_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1692_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(128), ack => type_cast_689_inst_req_0); -- 
    rr_1706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(128), ack => type_cast_699_inst_req_0); -- 
    rr_1720_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1720_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(128), ack => type_cast_709_inst_req_0); -- 
    rr_1734_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1734_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(128), ack => type_cast_719_inst_req_0); -- 
    rr_1748_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1748_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(128), ack => type_cast_729_inst_req_0); -- 
    rr_1762_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1762_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(128), ack => type_cast_739_inst_req_0); -- 
    -- CP-element group 129:  transition  input  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	128 
    -- CP-element group 129: successors 
    -- CP-element group 129:  members (3) 
      -- CP-element group 129: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_669_Sample/ra
      -- CP-element group 129: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_669_Sample/$exit
      -- CP-element group 129: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_669_sample_completed_
      -- 
    ra_1665_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_669_inst_ack_0, ack => zeropad3D_CP_676_elements(129)); -- 
    -- CP-element group 130:  transition  input  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	124 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	165 
    -- CP-element group 130:  members (3) 
      -- CP-element group 130: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_669_Update/$exit
      -- CP-element group 130: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_669_Update/ca
      -- CP-element group 130: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_669_update_completed_
      -- 
    ca_1670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_669_inst_ack_1, ack => zeropad3D_CP_676_elements(130)); -- 
    -- CP-element group 131:  transition  input  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	128 
    -- CP-element group 131: successors 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_679_Sample/ra
      -- CP-element group 131: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_679_Sample/$exit
      -- CP-element group 131: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_679_sample_completed_
      -- 
    ra_1679_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_679_inst_ack_0, ack => zeropad3D_CP_676_elements(131)); -- 
    -- CP-element group 132:  transition  input  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	124 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	162 
    -- CP-element group 132:  members (3) 
      -- CP-element group 132: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_679_Update/$exit
      -- CP-element group 132: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_679_Update/ca
      -- CP-element group 132: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_679_update_completed_
      -- 
    ca_1684_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_679_inst_ack_1, ack => zeropad3D_CP_676_elements(132)); -- 
    -- CP-element group 133:  transition  input  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	128 
    -- CP-element group 133: successors 
    -- CP-element group 133:  members (3) 
      -- CP-element group 133: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_689_Sample/ra
      -- CP-element group 133: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_689_sample_completed_
      -- CP-element group 133: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_689_Sample/$exit
      -- 
    ra_1693_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_689_inst_ack_0, ack => zeropad3D_CP_676_elements(133)); -- 
    -- CP-element group 134:  transition  input  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	124 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	159 
    -- CP-element group 134:  members (3) 
      -- CP-element group 134: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_689_update_completed_
      -- CP-element group 134: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_689_Update/$exit
      -- CP-element group 134: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_689_Update/ca
      -- 
    ca_1698_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_689_inst_ack_1, ack => zeropad3D_CP_676_elements(134)); -- 
    -- CP-element group 135:  transition  input  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	128 
    -- CP-element group 135: successors 
    -- CP-element group 135:  members (3) 
      -- CP-element group 135: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_699_Sample/ra
      -- CP-element group 135: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_699_Sample/$exit
      -- CP-element group 135: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_699_sample_completed_
      -- 
    ra_1707_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_699_inst_ack_0, ack => zeropad3D_CP_676_elements(135)); -- 
    -- CP-element group 136:  transition  input  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	124 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	156 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_699_Update/ca
      -- CP-element group 136: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_699_Update/$exit
      -- CP-element group 136: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_699_update_completed_
      -- 
    ca_1712_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_699_inst_ack_1, ack => zeropad3D_CP_676_elements(136)); -- 
    -- CP-element group 137:  transition  input  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	128 
    -- CP-element group 137: successors 
    -- CP-element group 137:  members (3) 
      -- CP-element group 137: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_709_Sample/ra
      -- CP-element group 137: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_709_Sample/$exit
      -- CP-element group 137: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_709_sample_completed_
      -- 
    ra_1721_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_709_inst_ack_0, ack => zeropad3D_CP_676_elements(137)); -- 
    -- CP-element group 138:  transition  input  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	124 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	153 
    -- CP-element group 138:  members (3) 
      -- CP-element group 138: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_709_Update/ca
      -- CP-element group 138: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_709_Update/$exit
      -- CP-element group 138: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_709_update_completed_
      -- 
    ca_1726_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_709_inst_ack_1, ack => zeropad3D_CP_676_elements(138)); -- 
    -- CP-element group 139:  transition  input  bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	128 
    -- CP-element group 139: successors 
    -- CP-element group 139:  members (3) 
      -- CP-element group 139: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_719_sample_completed_
      -- CP-element group 139: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_719_Sample/ra
      -- CP-element group 139: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_719_Sample/$exit
      -- 
    ra_1735_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_719_inst_ack_0, ack => zeropad3D_CP_676_elements(139)); -- 
    -- CP-element group 140:  transition  input  bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	124 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	150 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_719_update_completed_
      -- CP-element group 140: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_719_Update/ca
      -- CP-element group 140: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_719_Update/$exit
      -- 
    ca_1740_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_719_inst_ack_1, ack => zeropad3D_CP_676_elements(140)); -- 
    -- CP-element group 141:  transition  input  bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	128 
    -- CP-element group 141: successors 
    -- CP-element group 141:  members (3) 
      -- CP-element group 141: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_729_Sample/$exit
      -- CP-element group 141: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_729_Sample/ra
      -- CP-element group 141: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_729_sample_completed_
      -- 
    ra_1749_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_729_inst_ack_0, ack => zeropad3D_CP_676_elements(141)); -- 
    -- CP-element group 142:  transition  input  bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	124 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	147 
    -- CP-element group 142:  members (3) 
      -- CP-element group 142: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_729_Update/ca
      -- CP-element group 142: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_729_Update/$exit
      -- CP-element group 142: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_729_update_completed_
      -- 
    ca_1754_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_729_inst_ack_1, ack => zeropad3D_CP_676_elements(142)); -- 
    -- CP-element group 143:  transition  input  bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	128 
    -- CP-element group 143: successors 
    -- CP-element group 143:  members (3) 
      -- CP-element group 143: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_739_Sample/ra
      -- CP-element group 143: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_739_Sample/$exit
      -- CP-element group 143: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_739_sample_completed_
      -- 
    ra_1763_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_739_inst_ack_0, ack => zeropad3D_CP_676_elements(143)); -- 
    -- CP-element group 144:  transition  input  output  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	124 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	145 
    -- CP-element group 144:  members (6) 
      -- CP-element group 144: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_741_Sample/$entry
      -- CP-element group 144: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_741_Sample/req
      -- CP-element group 144: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_741_sample_start_
      -- CP-element group 144: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_739_Update/ca
      -- CP-element group 144: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_739_Update/$exit
      -- CP-element group 144: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/type_cast_739_update_completed_
      -- 
    ca_1768_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_739_inst_ack_1, ack => zeropad3D_CP_676_elements(144)); -- 
    req_1776_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1776_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(144), ack => WPIPE_zeropad_output_pipe_741_inst_req_0); -- 
    -- CP-element group 145:  transition  input  output  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	144 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	146 
    -- CP-element group 145:  members (6) 
      -- CP-element group 145: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_741_sample_completed_
      -- CP-element group 145: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_741_Sample/ack
      -- CP-element group 145: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_741_Update/req
      -- CP-element group 145: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_741_Update/$entry
      -- CP-element group 145: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_741_Sample/$exit
      -- CP-element group 145: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_741_update_start_
      -- 
    ack_1777_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_741_inst_ack_0, ack => zeropad3D_CP_676_elements(145)); -- 
    req_1781_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1781_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(145), ack => WPIPE_zeropad_output_pipe_741_inst_req_1); -- 
    -- CP-element group 146:  transition  input  bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	145 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	147 
    -- CP-element group 146:  members (3) 
      -- CP-element group 146: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_741_Update/$exit
      -- CP-element group 146: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_741_Update/ack
      -- CP-element group 146: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_741_update_completed_
      -- 
    ack_1782_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_741_inst_ack_1, ack => zeropad3D_CP_676_elements(146)); -- 
    -- CP-element group 147:  join  transition  output  bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	142 
    -- CP-element group 147: 	146 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	148 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_744_sample_start_
      -- CP-element group 147: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_744_Sample/req
      -- CP-element group 147: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_744_Sample/$entry
      -- 
    req_1790_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1790_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(147), ack => WPIPE_zeropad_output_pipe_744_inst_req_0); -- 
    zeropad3D_cp_element_group_147: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_147"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(142) & zeropad3D_CP_676_elements(146);
      gj_zeropad3D_cp_element_group_147 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(147), clk => clk, reset => reset); --
    end block;
    -- CP-element group 148:  transition  input  output  bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	147 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	149 
    -- CP-element group 148:  members (6) 
      -- CP-element group 148: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_744_sample_completed_
      -- CP-element group 148: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_744_Update/req
      -- CP-element group 148: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_744_Update/$entry
      -- CP-element group 148: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_744_Sample/ack
      -- CP-element group 148: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_744_Sample/$exit
      -- CP-element group 148: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_744_update_start_
      -- 
    ack_1791_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_744_inst_ack_0, ack => zeropad3D_CP_676_elements(148)); -- 
    req_1795_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1795_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(148), ack => WPIPE_zeropad_output_pipe_744_inst_req_1); -- 
    -- CP-element group 149:  transition  input  bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	148 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	150 
    -- CP-element group 149:  members (3) 
      -- CP-element group 149: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_744_Update/ack
      -- CP-element group 149: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_744_Update/$exit
      -- CP-element group 149: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_744_update_completed_
      -- 
    ack_1796_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_744_inst_ack_1, ack => zeropad3D_CP_676_elements(149)); -- 
    -- CP-element group 150:  join  transition  output  bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	140 
    -- CP-element group 150: 	149 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	151 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_747_Sample/req
      -- CP-element group 150: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_747_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_747_sample_start_
      -- 
    req_1804_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1804_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(150), ack => WPIPE_zeropad_output_pipe_747_inst_req_0); -- 
    zeropad3D_cp_element_group_150: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_150"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(140) & zeropad3D_CP_676_elements(149);
      gj_zeropad3D_cp_element_group_150 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(150), clk => clk, reset => reset); --
    end block;
    -- CP-element group 151:  transition  input  output  bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	150 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	152 
    -- CP-element group 151:  members (6) 
      -- CP-element group 151: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_747_Sample/$exit
      -- CP-element group 151: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_747_Sample/ack
      -- CP-element group 151: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_747_sample_completed_
      -- CP-element group 151: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_747_Update/$entry
      -- CP-element group 151: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_747_Update/req
      -- CP-element group 151: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_747_update_start_
      -- 
    ack_1805_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_747_inst_ack_0, ack => zeropad3D_CP_676_elements(151)); -- 
    req_1809_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1809_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(151), ack => WPIPE_zeropad_output_pipe_747_inst_req_1); -- 
    -- CP-element group 152:  transition  input  bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	151 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	153 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_747_Update/$exit
      -- CP-element group 152: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_747_Update/ack
      -- CP-element group 152: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_747_update_completed_
      -- 
    ack_1810_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_747_inst_ack_1, ack => zeropad3D_CP_676_elements(152)); -- 
    -- CP-element group 153:  join  transition  output  bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	138 
    -- CP-element group 153: 	152 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	154 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_750_Sample/req
      -- CP-element group 153: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_750_Sample/$entry
      -- CP-element group 153: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_750_sample_start_
      -- 
    req_1818_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1818_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(153), ack => WPIPE_zeropad_output_pipe_750_inst_req_0); -- 
    zeropad3D_cp_element_group_153: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_153"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(138) & zeropad3D_CP_676_elements(152);
      gj_zeropad3D_cp_element_group_153 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(153), clk => clk, reset => reset); --
    end block;
    -- CP-element group 154:  transition  input  output  bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	153 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	155 
    -- CP-element group 154:  members (6) 
      -- CP-element group 154: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_750_Update/req
      -- CP-element group 154: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_750_Update/$entry
      -- CP-element group 154: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_750_Sample/ack
      -- CP-element group 154: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_750_Sample/$exit
      -- CP-element group 154: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_750_update_start_
      -- CP-element group 154: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_750_sample_completed_
      -- 
    ack_1819_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_750_inst_ack_0, ack => zeropad3D_CP_676_elements(154)); -- 
    req_1823_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1823_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(154), ack => WPIPE_zeropad_output_pipe_750_inst_req_1); -- 
    -- CP-element group 155:  transition  input  bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	154 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	156 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_750_Update/ack
      -- CP-element group 155: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_750_Update/$exit
      -- CP-element group 155: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_750_update_completed_
      -- 
    ack_1824_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_750_inst_ack_1, ack => zeropad3D_CP_676_elements(155)); -- 
    -- CP-element group 156:  join  transition  output  bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	136 
    -- CP-element group 156: 	155 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	157 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_753_sample_start_
      -- CP-element group 156: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_753_Sample/req
      -- CP-element group 156: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_753_Sample/$entry
      -- 
    req_1832_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1832_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(156), ack => WPIPE_zeropad_output_pipe_753_inst_req_0); -- 
    zeropad3D_cp_element_group_156: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_156"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(136) & zeropad3D_CP_676_elements(155);
      gj_zeropad3D_cp_element_group_156 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(156), clk => clk, reset => reset); --
    end block;
    -- CP-element group 157:  transition  input  output  bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	156 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	158 
    -- CP-element group 157:  members (6) 
      -- CP-element group 157: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_753_Sample/$exit
      -- CP-element group 157: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_753_Update/req
      -- CP-element group 157: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_753_Update/$entry
      -- CP-element group 157: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_753_Sample/ack
      -- CP-element group 157: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_753_sample_completed_
      -- CP-element group 157: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_753_update_start_
      -- 
    ack_1833_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_753_inst_ack_0, ack => zeropad3D_CP_676_elements(157)); -- 
    req_1837_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1837_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(157), ack => WPIPE_zeropad_output_pipe_753_inst_req_1); -- 
    -- CP-element group 158:  transition  input  bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	157 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	159 
    -- CP-element group 158:  members (3) 
      -- CP-element group 158: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_753_Update/ack
      -- CP-element group 158: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_753_Update/$exit
      -- CP-element group 158: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_753_update_completed_
      -- 
    ack_1838_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_753_inst_ack_1, ack => zeropad3D_CP_676_elements(158)); -- 
    -- CP-element group 159:  join  transition  output  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	134 
    -- CP-element group 159: 	158 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	160 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_756_sample_start_
      -- CP-element group 159: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_756_Sample/req
      -- CP-element group 159: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_756_Sample/$entry
      -- 
    req_1846_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1846_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(159), ack => WPIPE_zeropad_output_pipe_756_inst_req_0); -- 
    zeropad3D_cp_element_group_159: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_159"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(134) & zeropad3D_CP_676_elements(158);
      gj_zeropad3D_cp_element_group_159 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(159), clk => clk, reset => reset); --
    end block;
    -- CP-element group 160:  transition  input  output  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	159 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	161 
    -- CP-element group 160:  members (6) 
      -- CP-element group 160: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_756_Update/req
      -- CP-element group 160: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_756_Update/$entry
      -- CP-element group 160: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_756_Sample/ack
      -- CP-element group 160: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_756_Sample/$exit
      -- CP-element group 160: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_756_update_start_
      -- CP-element group 160: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_756_sample_completed_
      -- 
    ack_1847_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_756_inst_ack_0, ack => zeropad3D_CP_676_elements(160)); -- 
    req_1851_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1851_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(160), ack => WPIPE_zeropad_output_pipe_756_inst_req_1); -- 
    -- CP-element group 161:  transition  input  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	160 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	162 
    -- CP-element group 161:  members (3) 
      -- CP-element group 161: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_756_Update/ack
      -- CP-element group 161: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_756_Update/$exit
      -- CP-element group 161: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_756_update_completed_
      -- 
    ack_1852_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_756_inst_ack_1, ack => zeropad3D_CP_676_elements(161)); -- 
    -- CP-element group 162:  join  transition  output  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	132 
    -- CP-element group 162: 	161 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	163 
    -- CP-element group 162:  members (3) 
      -- CP-element group 162: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_759_Sample/req
      -- CP-element group 162: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_759_Sample/$entry
      -- CP-element group 162: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_759_sample_start_
      -- 
    req_1860_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1860_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(162), ack => WPIPE_zeropad_output_pipe_759_inst_req_0); -- 
    zeropad3D_cp_element_group_162: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_162"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(132) & zeropad3D_CP_676_elements(161);
      gj_zeropad3D_cp_element_group_162 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(162), clk => clk, reset => reset); --
    end block;
    -- CP-element group 163:  transition  input  output  bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	162 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	164 
    -- CP-element group 163:  members (6) 
      -- CP-element group 163: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_759_Update/req
      -- CP-element group 163: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_759_Update/$entry
      -- CP-element group 163: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_759_Sample/ack
      -- CP-element group 163: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_759_Sample/$exit
      -- CP-element group 163: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_759_update_start_
      -- CP-element group 163: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_759_sample_completed_
      -- 
    ack_1861_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_759_inst_ack_0, ack => zeropad3D_CP_676_elements(163)); -- 
    req_1865_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1865_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(163), ack => WPIPE_zeropad_output_pipe_759_inst_req_1); -- 
    -- CP-element group 164:  transition  input  bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	163 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	165 
    -- CP-element group 164:  members (3) 
      -- CP-element group 164: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_759_Update/ack
      -- CP-element group 164: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_759_Update/$exit
      -- CP-element group 164: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_759_update_completed_
      -- 
    ack_1866_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_759_inst_ack_1, ack => zeropad3D_CP_676_elements(164)); -- 
    -- CP-element group 165:  join  transition  output  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	130 
    -- CP-element group 165: 	164 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	166 
    -- CP-element group 165:  members (3) 
      -- CP-element group 165: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_762_sample_start_
      -- CP-element group 165: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_762_Sample/req
      -- CP-element group 165: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_762_Sample/$entry
      -- 
    req_1874_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1874_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(165), ack => WPIPE_zeropad_output_pipe_762_inst_req_0); -- 
    zeropad3D_cp_element_group_165: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_165"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(130) & zeropad3D_CP_676_elements(164);
      gj_zeropad3D_cp_element_group_165 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(165), clk => clk, reset => reset); --
    end block;
    -- CP-element group 166:  transition  input  output  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	165 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	167 
    -- CP-element group 166:  members (6) 
      -- CP-element group 166: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_762_sample_completed_
      -- CP-element group 166: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_762_Update/$entry
      -- CP-element group 166: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_762_Sample/ack
      -- CP-element group 166: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_762_Sample/$exit
      -- CP-element group 166: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_762_Update/req
      -- CP-element group 166: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_762_update_start_
      -- 
    ack_1875_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_762_inst_ack_0, ack => zeropad3D_CP_676_elements(166)); -- 
    req_1879_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1879_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(166), ack => WPIPE_zeropad_output_pipe_762_inst_req_1); -- 
    -- CP-element group 167:  fork  transition  place  input  output  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	166 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	168 
    -- CP-element group 167: 	169 
    -- CP-element group 167:  members (13) 
      -- CP-element group 167: 	 branch_block_stmt_224/assign_stmt_770_to_call_stmt_777__entry__
      -- CP-element group 167: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764__exit__
      -- CP-element group 167: 	 branch_block_stmt_224/assign_stmt_770_to_call_stmt_777/call_stmt_777_Update/ccr
      -- CP-element group 167: 	 branch_block_stmt_224/assign_stmt_770_to_call_stmt_777/$entry
      -- CP-element group 167: 	 branch_block_stmt_224/assign_stmt_770_to_call_stmt_777/call_stmt_777_Update/$entry
      -- CP-element group 167: 	 branch_block_stmt_224/assign_stmt_770_to_call_stmt_777/call_stmt_777_sample_start_
      -- CP-element group 167: 	 branch_block_stmt_224/assign_stmt_770_to_call_stmt_777/call_stmt_777_Sample/crr
      -- CP-element group 167: 	 branch_block_stmt_224/assign_stmt_770_to_call_stmt_777/call_stmt_777_Sample/$entry
      -- CP-element group 167: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_762_Update/ack
      -- CP-element group 167: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_762_Update/$exit
      -- CP-element group 167: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/WPIPE_zeropad_output_pipe_762_update_completed_
      -- CP-element group 167: 	 branch_block_stmt_224/assign_stmt_770_to_call_stmt_777/call_stmt_777_update_start_
      -- CP-element group 167: 	 branch_block_stmt_224/call_stmt_656_to_assign_stmt_764/$exit
      -- 
    ack_1880_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_zeropad_output_pipe_762_inst_ack_1, ack => zeropad3D_CP_676_elements(167)); -- 
    ccr_1896_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1896_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(167), ack => call_stmt_777_call_req_1); -- 
    crr_1891_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1891_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(167), ack => call_stmt_777_call_req_0); -- 
    -- CP-element group 168:  transition  input  bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	167 
    -- CP-element group 168: successors 
    -- CP-element group 168:  members (3) 
      -- CP-element group 168: 	 branch_block_stmt_224/assign_stmt_770_to_call_stmt_777/call_stmt_777_Sample/cra
      -- CP-element group 168: 	 branch_block_stmt_224/assign_stmt_770_to_call_stmt_777/call_stmt_777_Sample/$exit
      -- CP-element group 168: 	 branch_block_stmt_224/assign_stmt_770_to_call_stmt_777/call_stmt_777_sample_completed_
      -- 
    cra_1892_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_777_call_ack_0, ack => zeropad3D_CP_676_elements(168)); -- 
    -- CP-element group 169:  transition  place  input  bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	167 
    -- CP-element group 169: successors 
    -- CP-element group 169:  members (16) 
      -- CP-element group 169: 	 branch_block_stmt_224/assign_stmt_770_to_call_stmt_777__exit__
      -- CP-element group 169: 	 $exit
      -- CP-element group 169: 	 branch_block_stmt_224/branch_block_stmt_224__exit__
      -- CP-element group 169: 	 branch_block_stmt_224/$exit
      -- CP-element group 169: 	 branch_block_stmt_224/merge_stmt_779__exit__
      -- CP-element group 169: 	 branch_block_stmt_224/assign_stmt_770_to_call_stmt_777/call_stmt_777_Update/$exit
      -- CP-element group 169: 	 branch_block_stmt_224/return__
      -- CP-element group 169: 	 branch_block_stmt_224/assign_stmt_770_to_call_stmt_777/$exit
      -- CP-element group 169: 	 branch_block_stmt_224/assign_stmt_770_to_call_stmt_777/call_stmt_777_Update/cca
      -- CP-element group 169: 	 branch_block_stmt_224/assign_stmt_770_to_call_stmt_777/call_stmt_777_update_completed_
      -- CP-element group 169: 	 branch_block_stmt_224/return___PhiReq/$entry
      -- CP-element group 169: 	 branch_block_stmt_224/return___PhiReq/$exit
      -- CP-element group 169: 	 branch_block_stmt_224/merge_stmt_779_PhiReqMerge
      -- CP-element group 169: 	 branch_block_stmt_224/merge_stmt_779_PhiAck/$entry
      -- CP-element group 169: 	 branch_block_stmt_224/merge_stmt_779_PhiAck/$exit
      -- CP-element group 169: 	 branch_block_stmt_224/merge_stmt_779_PhiAck/dummy
      -- 
    cca_1897_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_777_call_ack_1, ack => zeropad3D_CP_676_elements(169)); -- 
    -- CP-element group 170:  transition  output  delay-element  bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	60 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	174 
    -- CP-element group 170:  members (5) 
      -- CP-element group 170: 	 branch_block_stmt_224/bbx_xnph_forx_xbody_PhiReq/$exit
      -- CP-element group 170: 	 branch_block_stmt_224/bbx_xnph_forx_xbody_PhiReq/phi_stmt_450/$exit
      -- CP-element group 170: 	 branch_block_stmt_224/bbx_xnph_forx_xbody_PhiReq/phi_stmt_450/phi_stmt_450_sources/$exit
      -- CP-element group 170: 	 branch_block_stmt_224/bbx_xnph_forx_xbody_PhiReq/phi_stmt_450/phi_stmt_450_sources/type_cast_454_konst_delay_trans
      -- CP-element group 170: 	 branch_block_stmt_224/bbx_xnph_forx_xbody_PhiReq/phi_stmt_450/phi_stmt_450_req
      -- 
    phi_stmt_450_req_1920_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_450_req_1920_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(170), ack => phi_stmt_450_req_0); -- 
    -- Element group zeropad3D_CP_676_elements(170) is a control-delay.
    cp_element_170_delay: control_delay_element  generic map(name => " 170_delay", delay_value => 1)  port map(req => zeropad3D_CP_676_elements(60), ack => zeropad3D_CP_676_elements(170), clk => clk, reset =>reset);
    -- CP-element group 171:  transition  input  bypass 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	103 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	173 
    -- CP-element group 171:  members (2) 
      -- CP-element group 171: 	 branch_block_stmt_224/forx_xbody_forx_xbody_PhiReq/phi_stmt_450/phi_stmt_450_sources/type_cast_456/SplitProtocol/Sample/$exit
      -- CP-element group 171: 	 branch_block_stmt_224/forx_xbody_forx_xbody_PhiReq/phi_stmt_450/phi_stmt_450_sources/type_cast_456/SplitProtocol/Sample/ra
      -- 
    ra_1940_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_456_inst_ack_0, ack => zeropad3D_CP_676_elements(171)); -- 
    -- CP-element group 172:  transition  input  bypass 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	103 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	173 
    -- CP-element group 172:  members (2) 
      -- CP-element group 172: 	 branch_block_stmt_224/forx_xbody_forx_xbody_PhiReq/phi_stmt_450/phi_stmt_450_sources/type_cast_456/SplitProtocol/Update/$exit
      -- CP-element group 172: 	 branch_block_stmt_224/forx_xbody_forx_xbody_PhiReq/phi_stmt_450/phi_stmt_450_sources/type_cast_456/SplitProtocol/Update/ca
      -- 
    ca_1945_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_456_inst_ack_1, ack => zeropad3D_CP_676_elements(172)); -- 
    -- CP-element group 173:  join  transition  output  bypass 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	171 
    -- CP-element group 173: 	172 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	174 
    -- CP-element group 173:  members (6) 
      -- CP-element group 173: 	 branch_block_stmt_224/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 173: 	 branch_block_stmt_224/forx_xbody_forx_xbody_PhiReq/phi_stmt_450/$exit
      -- CP-element group 173: 	 branch_block_stmt_224/forx_xbody_forx_xbody_PhiReq/phi_stmt_450/phi_stmt_450_sources/$exit
      -- CP-element group 173: 	 branch_block_stmt_224/forx_xbody_forx_xbody_PhiReq/phi_stmt_450/phi_stmt_450_sources/type_cast_456/$exit
      -- CP-element group 173: 	 branch_block_stmt_224/forx_xbody_forx_xbody_PhiReq/phi_stmt_450/phi_stmt_450_sources/type_cast_456/SplitProtocol/$exit
      -- CP-element group 173: 	 branch_block_stmt_224/forx_xbody_forx_xbody_PhiReq/phi_stmt_450/phi_stmt_450_req
      -- 
    phi_stmt_450_req_1946_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_450_req_1946_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(173), ack => phi_stmt_450_req_1); -- 
    zeropad3D_cp_element_group_173: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "zeropad3D_cp_element_group_173"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_CP_676_elements(171) & zeropad3D_CP_676_elements(172);
      gj_zeropad3D_cp_element_group_173 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_CP_676_elements(173), clk => clk, reset => reset); --
    end block;
    -- CP-element group 174:  merge  transition  place  bypass 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	170 
    -- CP-element group 174: 	173 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	175 
    -- CP-element group 174:  members (2) 
      -- CP-element group 174: 	 branch_block_stmt_224/merge_stmt_449_PhiReqMerge
      -- CP-element group 174: 	 branch_block_stmt_224/merge_stmt_449_PhiAck/$entry
      -- 
    zeropad3D_CP_676_elements(174) <= OrReduce(zeropad3D_CP_676_elements(170) & zeropad3D_CP_676_elements(173));
    -- CP-element group 175:  fork  transition  place  input  output  bypass 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	174 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	62 
    -- CP-element group 175: 	63 
    -- CP-element group 175: 	65 
    -- CP-element group 175: 	66 
    -- CP-element group 175: 	69 
    -- CP-element group 175: 	73 
    -- CP-element group 175: 	77 
    -- CP-element group 175: 	81 
    -- CP-element group 175: 	85 
    -- CP-element group 175: 	89 
    -- CP-element group 175: 	93 
    -- CP-element group 175: 	97 
    -- CP-element group 175: 	100 
    -- CP-element group 175:  members (56) 
      -- CP-element group 175: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612__entry__
      -- CP-element group 175: 	 branch_block_stmt_224/merge_stmt_449__exit__
      -- CP-element group 175: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/$entry
      -- CP-element group 175: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/addr_of_463_update_start_
      -- CP-element group 175: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/array_obj_ref_462_index_resized_1
      -- CP-element group 175: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/array_obj_ref_462_index_scaled_1
      -- CP-element group 175: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/array_obj_ref_462_index_computed_1
      -- CP-element group 175: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/array_obj_ref_462_index_resize_1/$entry
      -- CP-element group 175: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/array_obj_ref_462_index_resize_1/$exit
      -- CP-element group 175: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/array_obj_ref_462_index_resize_1/index_resize_req
      -- CP-element group 175: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/array_obj_ref_462_index_resize_1/index_resize_ack
      -- CP-element group 175: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/array_obj_ref_462_index_scale_1/$entry
      -- CP-element group 175: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/array_obj_ref_462_index_scale_1/$exit
      -- CP-element group 175: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/array_obj_ref_462_index_scale_1/scale_rename_req
      -- CP-element group 175: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/array_obj_ref_462_index_scale_1/scale_rename_ack
      -- CP-element group 175: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/array_obj_ref_462_final_index_sum_regn_update_start
      -- CP-element group 175: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/array_obj_ref_462_final_index_sum_regn_Sample/$entry
      -- CP-element group 175: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/array_obj_ref_462_final_index_sum_regn_Sample/req
      -- CP-element group 175: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/array_obj_ref_462_final_index_sum_regn_Update/$entry
      -- CP-element group 175: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/array_obj_ref_462_final_index_sum_regn_Update/req
      -- CP-element group 175: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/addr_of_463_complete/$entry
      -- CP-element group 175: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/addr_of_463_complete/req
      -- CP-element group 175: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_466_sample_start_
      -- CP-element group 175: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_466_Sample/$entry
      -- CP-element group 175: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/RPIPE_zeropad_input_pipe_466_Sample/rr
      -- CP-element group 175: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_470_update_start_
      -- CP-element group 175: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_470_Update/$entry
      -- CP-element group 175: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_470_Update/cr
      -- CP-element group 175: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_483_update_start_
      -- CP-element group 175: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_483_Update/$entry
      -- CP-element group 175: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_483_Update/cr
      -- CP-element group 175: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_501_update_start_
      -- CP-element group 175: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_501_Update/$entry
      -- CP-element group 175: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_501_Update/cr
      -- CP-element group 175: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_519_update_start_
      -- CP-element group 175: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_519_Update/$entry
      -- CP-element group 175: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_519_Update/cr
      -- CP-element group 175: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_537_update_start_
      -- CP-element group 175: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_537_Update/$entry
      -- CP-element group 175: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_537_Update/cr
      -- CP-element group 175: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_555_update_start_
      -- CP-element group 175: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_555_Update/$entry
      -- CP-element group 175: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_555_Update/cr
      -- CP-element group 175: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_573_update_start_
      -- CP-element group 175: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_573_Update/$entry
      -- CP-element group 175: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_573_Update/cr
      -- CP-element group 175: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_591_update_start_
      -- CP-element group 175: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_591_Update/$entry
      -- CP-element group 175: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/type_cast_591_Update/cr
      -- CP-element group 175: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/ptr_deref_599_update_start_
      -- CP-element group 175: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/ptr_deref_599_Update/$entry
      -- CP-element group 175: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/ptr_deref_599_Update/word_access_complete/$entry
      -- CP-element group 175: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/ptr_deref_599_Update/word_access_complete/word_0/$entry
      -- CP-element group 175: 	 branch_block_stmt_224/assign_stmt_464_to_assign_stmt_612/ptr_deref_599_Update/word_access_complete/word_0/cr
      -- CP-element group 175: 	 branch_block_stmt_224/merge_stmt_449_PhiAck/$exit
      -- CP-element group 175: 	 branch_block_stmt_224/merge_stmt_449_PhiAck/phi_stmt_450_ack
      -- 
    phi_stmt_450_ack_1951_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_450_ack_0, ack => zeropad3D_CP_676_elements(175)); -- 
    req_1168_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1168_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(175), ack => array_obj_ref_462_index_offset_req_0); -- 
    req_1173_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1173_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(175), ack => array_obj_ref_462_index_offset_req_1); -- 
    req_1188_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1188_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(175), ack => addr_of_463_final_reg_req_1); -- 
    rr_1197_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1197_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(175), ack => RPIPE_zeropad_input_pipe_466_inst_req_0); -- 
    cr_1216_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1216_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(175), ack => type_cast_470_inst_req_1); -- 
    cr_1244_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1244_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(175), ack => type_cast_483_inst_req_1); -- 
    cr_1272_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1272_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(175), ack => type_cast_501_inst_req_1); -- 
    cr_1300_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1300_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(175), ack => type_cast_519_inst_req_1); -- 
    cr_1328_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1328_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(175), ack => type_cast_537_inst_req_1); -- 
    cr_1356_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1356_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(175), ack => type_cast_555_inst_req_1); -- 
    cr_1384_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1384_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(175), ack => type_cast_573_inst_req_1); -- 
    cr_1412_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1412_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(175), ack => type_cast_591_inst_req_1); -- 
    cr_1462_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1462_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(175), ack => ptr_deref_599_store_0_req_1); -- 
    -- CP-element group 176:  merge  fork  transition  place  output  bypass 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	61 
    -- CP-element group 176: 	102 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	104 
    -- CP-element group 176: 	105 
    -- CP-element group 176: 	107 
    -- CP-element group 176: 	108 
    -- CP-element group 176: 	122 
    -- CP-element group 176:  members (22) 
      -- CP-element group 176: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_630_sample_start_
      -- CP-element group 176: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653__entry__
      -- CP-element group 176: 	 branch_block_stmt_224/merge_stmt_621__exit__
      -- CP-element group 176: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/call_stmt_624_Update/$entry
      -- CP-element group 176: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_630_Sample/$entry
      -- CP-element group 176: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/WPIPE_Block0_starting_630_Sample/req
      -- CP-element group 176: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/call_stmt_624_Update/ccr
      -- CP-element group 176: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/type_cast_628_update_start_
      -- CP-element group 176: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/call_stmt_624_Sample/crr
      -- CP-element group 176: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/call_stmt_624_sample_start_
      -- CP-element group 176: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/call_stmt_624_Sample/$entry
      -- CP-element group 176: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/$entry
      -- CP-element group 176: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/call_stmt_624_update_start_
      -- CP-element group 176: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/type_cast_628_Update/cr
      -- CP-element group 176: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/type_cast_628_Update/$entry
      -- CP-element group 176: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/RPIPE_Block0_complete_652_Sample/rr
      -- CP-element group 176: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/RPIPE_Block0_complete_652_Sample/$entry
      -- CP-element group 176: 	 branch_block_stmt_224/call_stmt_624_to_assign_stmt_653/RPIPE_Block0_complete_652_sample_start_
      -- CP-element group 176: 	 branch_block_stmt_224/merge_stmt_621_PhiReqMerge
      -- CP-element group 176: 	 branch_block_stmt_224/merge_stmt_621_PhiAck/$entry
      -- CP-element group 176: 	 branch_block_stmt_224/merge_stmt_621_PhiAck/$exit
      -- CP-element group 176: 	 branch_block_stmt_224/merge_stmt_621_PhiAck/dummy
      -- 
    req_1521_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1521_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(176), ack => WPIPE_Block0_starting_630_inst_req_0); -- 
    ccr_1498_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1498_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(176), ack => call_stmt_624_call_req_1); -- 
    crr_1493_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1493_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(176), ack => call_stmt_624_call_req_0); -- 
    cr_1512_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1512_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(176), ack => type_cast_628_inst_req_1); -- 
    rr_1619_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1619_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_CP_676_elements(176), ack => RPIPE_Block0_complete_652_inst_req_0); -- 
    zeropad3D_CP_676_elements(176) <= OrReduce(zeropad3D_CP_676_elements(61) & zeropad3D_CP_676_elements(102));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i64_i64_413_wire : std_logic_vector(63 downto 0);
    signal R_indvar_461_resized : std_logic_vector(13 downto 0);
    signal R_indvar_461_scaled : std_logic_vector(13 downto 0);
    signal add104_525 : std_logic_vector(63 downto 0);
    signal add110_543 : std_logic_vector(63 downto 0);
    signal add116_561 : std_logic_vector(63 downto 0);
    signal add122_579 : std_logic_vector(63 downto 0);
    signal add128_597 : std_logic_vector(63 downto 0);
    signal add23_261 : std_logic_vector(63 downto 0);
    signal add32_286 : std_logic_vector(63 downto 0);
    signal add41_311 : std_logic_vector(63 downto 0);
    signal add51_339 : std_logic_vector(31 downto 0);
    signal add60_364 : std_logic_vector(31 downto 0);
    signal add69_389 : std_logic_vector(31 downto 0);
    signal add92_489 : std_logic_vector(63 downto 0);
    signal add98_507 : std_logic_vector(63 downto 0);
    signal array_obj_ref_462_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_462_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_462_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_462_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_462_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_462_root_address : std_logic_vector(13 downto 0);
    signal arrayidx_464 : std_logic_vector(31 downto 0);
    signal call101_516 : std_logic_vector(7 downto 0);
    signal call107_534 : std_logic_vector(7 downto 0);
    signal call113_552 : std_logic_vector(7 downto 0);
    signal call119_570 : std_logic_vector(7 downto 0);
    signal call11_236 : std_logic_vector(7 downto 0);
    signal call125_588 : std_logic_vector(7 downto 0);
    signal call133_624 : std_logic_vector(63 downto 0);
    signal call149_653 : std_logic_vector(7 downto 0);
    signal call152_656 : std_logic_vector(63 downto 0);
    signal call16_239 : std_logic_vector(7 downto 0);
    signal call21_252 : std_logic_vector(7 downto 0);
    signal call25_264 : std_logic_vector(7 downto 0);
    signal call2_230 : std_logic_vector(7 downto 0);
    signal call30_277 : std_logic_vector(7 downto 0);
    signal call34_289 : std_logic_vector(7 downto 0);
    signal call39_302 : std_logic_vector(7 downto 0);
    signal call43_314 : std_logic_vector(7 downto 0);
    signal call44_317 : std_logic_vector(7 downto 0);
    signal call49_330 : std_logic_vector(7 downto 0);
    signal call53_342 : std_logic_vector(7 downto 0);
    signal call58_355 : std_logic_vector(7 downto 0);
    signal call62_367 : std_logic_vector(7 downto 0);
    signal call67_380 : std_logic_vector(7 downto 0);
    signal call6_233 : std_logic_vector(7 downto 0);
    signal call85_467 : std_logic_vector(7 downto 0);
    signal call89_480 : std_logic_vector(7 downto 0);
    signal call95_498 : std_logic_vector(7 downto 0);
    signal call_227 : std_logic_vector(7 downto 0);
    signal cmp229_421 : std_logic_vector(0 downto 0);
    signal conv103_520 : std_logic_vector(63 downto 0);
    signal conv109_538 : std_logic_vector(63 downto 0);
    signal conv115_556 : std_logic_vector(63 downto 0);
    signal conv121_574 : std_logic_vector(63 downto 0);
    signal conv127_592 : std_logic_vector(63 downto 0);
    signal conv134_629 : std_logic_vector(63 downto 0);
    signal conv153_661 : std_logic_vector(63 downto 0);
    signal conv159_670 : std_logic_vector(7 downto 0);
    signal conv165_680 : std_logic_vector(7 downto 0);
    signal conv171_690 : std_logic_vector(7 downto 0);
    signal conv177_700 : std_logic_vector(7 downto 0);
    signal conv183_710 : std_logic_vector(7 downto 0);
    signal conv189_720 : std_logic_vector(7 downto 0);
    signal conv195_730 : std_logic_vector(7 downto 0);
    signal conv19_243 : std_logic_vector(63 downto 0);
    signal conv201_740 : std_logic_vector(7 downto 0);
    signal conv22_256 : std_logic_vector(63 downto 0);
    signal conv28_268 : std_logic_vector(63 downto 0);
    signal conv31_281 : std_logic_vector(63 downto 0);
    signal conv37_293 : std_logic_vector(63 downto 0);
    signal conv40_306 : std_logic_vector(63 downto 0);
    signal conv47_321 : std_logic_vector(31 downto 0);
    signal conv50_334 : std_logic_vector(31 downto 0);
    signal conv56_346 : std_logic_vector(31 downto 0);
    signal conv59_359 : std_logic_vector(31 downto 0);
    signal conv65_371 : std_logic_vector(31 downto 0);
    signal conv68_384 : std_logic_vector(31 downto 0);
    signal conv79_415 : std_logic_vector(63 downto 0);
    signal conv86_471 : std_logic_vector(63 downto 0);
    signal conv91_484 : std_logic_vector(63 downto 0);
    signal conv97_502 : std_logic_vector(63 downto 0);
    signal exitcond3_612 : std_logic_vector(0 downto 0);
    signal indvar_450 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_607 : std_logic_vector(63 downto 0);
    signal mul223_770 : std_logic_vector(31 downto 0);
    signal mul226_775 : std_logic_vector(31 downto 0);
    signal mul78_400 : std_logic_vector(63 downto 0);
    signal mul_395 : std_logic_vector(63 downto 0);
    signal ptr_deref_599_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_599_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_599_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_599_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_599_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_599_word_offset_0 : std_logic_vector(13 downto 0);
    signal sext_405 : std_logic_vector(63 downto 0);
    signal shl100_513 : std_logic_vector(63 downto 0);
    signal shl106_531 : std_logic_vector(63 downto 0);
    signal shl112_549 : std_logic_vector(63 downto 0);
    signal shl118_567 : std_logic_vector(63 downto 0);
    signal shl124_585 : std_logic_vector(63 downto 0);
    signal shl20_249 : std_logic_vector(63 downto 0);
    signal shl29_274 : std_logic_vector(63 downto 0);
    signal shl38_299 : std_logic_vector(63 downto 0);
    signal shl48_327 : std_logic_vector(31 downto 0);
    signal shl57_352 : std_logic_vector(31 downto 0);
    signal shl66_377 : std_logic_vector(31 downto 0);
    signal shl88_477 : std_logic_vector(63 downto 0);
    signal shl94_495 : std_logic_vector(63 downto 0);
    signal shr162_676 : std_logic_vector(63 downto 0);
    signal shr168_686 : std_logic_vector(63 downto 0);
    signal shr174_696 : std_logic_vector(63 downto 0);
    signal shr180_706 : std_logic_vector(63 downto 0);
    signal shr186_716 : std_logic_vector(63 downto 0);
    signal shr192_726 : std_logic_vector(63 downto 0);
    signal shr198_736 : std_logic_vector(63 downto 0);
    signal shr_434 : std_logic_vector(63 downto 0);
    signal sub_666 : std_logic_vector(63 downto 0);
    signal tmp1_440 : std_logic_vector(0 downto 0);
    signal type_cast_247_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_272_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_297_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_325_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_350_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_375_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_393_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_409_wire : std_logic_vector(63 downto 0);
    signal type_cast_412_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_419_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_432_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_438_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_445_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_454_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_456_wire : std_logic_vector(63 downto 0);
    signal type_cast_475_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_493_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_511_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_529_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_547_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_565_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_583_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_605_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_627_wire : std_logic_vector(63 downto 0);
    signal type_cast_659_wire : std_logic_vector(63 downto 0);
    signal type_cast_674_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_684_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_694_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_704_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_714_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_724_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_734_wire_constant : std_logic_vector(63 downto 0);
    signal umax2_447 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    array_obj_ref_462_constant_part_of_offset <= "00000000000000";
    array_obj_ref_462_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_462_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_462_resized_base_address <= "00000000000000";
    ptr_deref_599_word_offset_0 <= "00000000000000";
    type_cast_247_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_272_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_297_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_325_wire_constant <= "00000000000000000000000000001000";
    type_cast_350_wire_constant <= "00000000000000000000000000001000";
    type_cast_375_wire_constant <= "00000000000000000000000000001000";
    type_cast_393_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_412_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_419_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000111";
    type_cast_432_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    type_cast_438_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_445_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_454_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_475_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_493_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_511_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_529_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_547_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_565_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_583_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_605_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_674_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_684_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_694_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_704_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_714_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_724_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_734_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    phi_stmt_450: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_454_wire_constant & type_cast_456_wire;
      req <= phi_stmt_450_req_0 & phi_stmt_450_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_450",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_450_ack_0,
          idata => idata,
          odata => indvar_450,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_450
    -- flow-through select operator MUX_446_inst
    umax2_447 <= shr_434 when (tmp1_440(0) /=  '0') else type_cast_445_wire_constant;
    addr_of_463_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_463_final_reg_req_0;
      addr_of_463_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_463_final_reg_req_1;
      addr_of_463_final_reg_ack_1<= rack(0);
      addr_of_463_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_463_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_462_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_464,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_242_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_242_inst_req_0;
      type_cast_242_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_242_inst_req_1;
      type_cast_242_inst_ack_1<= rack(0);
      type_cast_242_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_242_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call16_239,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv19_243,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_255_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_255_inst_req_0;
      type_cast_255_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_255_inst_req_1;
      type_cast_255_inst_ack_1<= rack(0);
      type_cast_255_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_255_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call21_252,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv22_256,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_267_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_267_inst_req_0;
      type_cast_267_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_267_inst_req_1;
      type_cast_267_inst_ack_1<= rack(0);
      type_cast_267_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_267_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call25_264,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv28_268,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_280_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_280_inst_req_0;
      type_cast_280_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_280_inst_req_1;
      type_cast_280_inst_ack_1<= rack(0);
      type_cast_280_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_280_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call30_277,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv31_281,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_292_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_292_inst_req_0;
      type_cast_292_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_292_inst_req_1;
      type_cast_292_inst_ack_1<= rack(0);
      type_cast_292_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_292_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call34_289,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv37_293,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_305_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_305_inst_req_0;
      type_cast_305_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_305_inst_req_1;
      type_cast_305_inst_ack_1<= rack(0);
      type_cast_305_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_305_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call39_302,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv40_306,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_320_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_320_inst_req_0;
      type_cast_320_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_320_inst_req_1;
      type_cast_320_inst_ack_1<= rack(0);
      type_cast_320_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_320_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call44_317,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv47_321,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_333_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_333_inst_req_0;
      type_cast_333_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_333_inst_req_1;
      type_cast_333_inst_ack_1<= rack(0);
      type_cast_333_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_333_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call49_330,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv50_334,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_345_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_345_inst_req_0;
      type_cast_345_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_345_inst_req_1;
      type_cast_345_inst_ack_1<= rack(0);
      type_cast_345_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_345_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call53_342,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv56_346,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_358_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_358_inst_req_0;
      type_cast_358_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_358_inst_req_1;
      type_cast_358_inst_ack_1<= rack(0);
      type_cast_358_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_358_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call58_355,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv59_359,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_370_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_370_inst_req_0;
      type_cast_370_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_370_inst_req_1;
      type_cast_370_inst_ack_1<= rack(0);
      type_cast_370_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_370_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call62_367,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv65_371,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_383_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_383_inst_req_0;
      type_cast_383_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_383_inst_req_1;
      type_cast_383_inst_ack_1<= rack(0);
      type_cast_383_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_383_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call67_380,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv68_384,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_409_inst
    process(sext_405) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := sext_405(63 downto 0);
      type_cast_409_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_414_inst
    process(ASHR_i64_i64_413_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := ASHR_i64_i64_413_wire(63 downto 0);
      conv79_415 <= tmp_var; -- 
    end process;
    type_cast_456_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_456_inst_req_0;
      type_cast_456_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_456_inst_req_1;
      type_cast_456_inst_ack_1<= rack(0);
      type_cast_456_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_456_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_607,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_456_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_470_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_470_inst_req_0;
      type_cast_470_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_470_inst_req_1;
      type_cast_470_inst_ack_1<= rack(0);
      type_cast_470_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_470_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call85_467,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv86_471,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_483_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_483_inst_req_0;
      type_cast_483_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_483_inst_req_1;
      type_cast_483_inst_ack_1<= rack(0);
      type_cast_483_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_483_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call89_480,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv91_484,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_501_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_501_inst_req_0;
      type_cast_501_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_501_inst_req_1;
      type_cast_501_inst_ack_1<= rack(0);
      type_cast_501_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_501_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call95_498,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv97_502,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_519_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_519_inst_req_0;
      type_cast_519_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_519_inst_req_1;
      type_cast_519_inst_ack_1<= rack(0);
      type_cast_519_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_519_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call101_516,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv103_520,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_537_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_537_inst_req_0;
      type_cast_537_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_537_inst_req_1;
      type_cast_537_inst_ack_1<= rack(0);
      type_cast_537_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_537_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call107_534,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv109_538,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_555_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_555_inst_req_0;
      type_cast_555_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_555_inst_req_1;
      type_cast_555_inst_ack_1<= rack(0);
      type_cast_555_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_555_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call113_552,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv115_556,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_573_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_573_inst_req_0;
      type_cast_573_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_573_inst_req_1;
      type_cast_573_inst_ack_1<= rack(0);
      type_cast_573_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_573_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call119_570,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv121_574,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_591_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_591_inst_req_0;
      type_cast_591_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_591_inst_req_1;
      type_cast_591_inst_ack_1<= rack(0);
      type_cast_591_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_591_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call125_588,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv127_592,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_628_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_628_inst_req_0;
      type_cast_628_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_628_inst_req_1;
      type_cast_628_inst_ack_1<= rack(0);
      type_cast_628_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_628_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_627_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv134_629,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_660_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_660_inst_req_0;
      type_cast_660_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_660_inst_req_1;
      type_cast_660_inst_ack_1<= rack(0);
      type_cast_660_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_660_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_659_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv153_661,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_669_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_669_inst_req_0;
      type_cast_669_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_669_inst_req_1;
      type_cast_669_inst_ack_1<= rack(0);
      type_cast_669_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_669_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub_666,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv159_670,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_679_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_679_inst_req_0;
      type_cast_679_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_679_inst_req_1;
      type_cast_679_inst_ack_1<= rack(0);
      type_cast_679_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_679_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr162_676,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv165_680,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_689_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_689_inst_req_0;
      type_cast_689_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_689_inst_req_1;
      type_cast_689_inst_ack_1<= rack(0);
      type_cast_689_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_689_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr168_686,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv171_690,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_699_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_699_inst_req_0;
      type_cast_699_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_699_inst_req_1;
      type_cast_699_inst_ack_1<= rack(0);
      type_cast_699_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_699_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr174_696,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv177_700,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_709_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_709_inst_req_0;
      type_cast_709_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_709_inst_req_1;
      type_cast_709_inst_ack_1<= rack(0);
      type_cast_709_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_709_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr180_706,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv183_710,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_719_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_719_inst_req_0;
      type_cast_719_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_719_inst_req_1;
      type_cast_719_inst_ack_1<= rack(0);
      type_cast_719_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_719_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr186_716,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv189_720,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_729_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_729_inst_req_0;
      type_cast_729_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_729_inst_req_1;
      type_cast_729_inst_ack_1<= rack(0);
      type_cast_729_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_729_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr192_726,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv195_730,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_739_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_739_inst_req_0;
      type_cast_739_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_739_inst_req_1;
      type_cast_739_inst_ack_1<= rack(0);
      type_cast_739_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_739_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr198_736,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv201_740,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_462_index_1_rename
    process(R_indvar_461_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_461_resized;
      ov(13 downto 0) := iv;
      R_indvar_461_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_462_index_1_resize
    process(indvar_450) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_450;
      ov := iv(13 downto 0);
      R_indvar_461_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_462_root_address_inst
    process(array_obj_ref_462_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_462_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_462_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_599_addr_0
    process(ptr_deref_599_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_599_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_599_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_599_base_resize
    process(arrayidx_464) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_464;
      ov := iv(13 downto 0);
      ptr_deref_599_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_599_gather_scatter
    process(add128_597) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add128_597;
      ov(63 downto 0) := iv;
      ptr_deref_599_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_599_root_address_inst
    process(ptr_deref_599_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_599_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_599_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_422_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp229_421;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_422_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_422_branch_req_0,
          ack0 => if_stmt_422_branch_ack_0,
          ack1 => if_stmt_422_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_613_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond3_612;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_613_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_613_branch_req_0,
          ack0 => if_stmt_613_branch_ack_0,
          ack1 => if_stmt_613_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u64_u64_606_inst
    process(indvar_450) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_450, type_cast_605_wire_constant, tmp_var);
      indvarx_xnext_607 <= tmp_var; --
    end process;
    -- binary operator ASHR_i64_i64_413_inst
    process(type_cast_409_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_409_wire, type_cast_412_wire_constant, tmp_var);
      ASHR_i64_i64_413_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_611_inst
    process(indvarx_xnext_607, umax2_447) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_607, umax2_447, tmp_var);
      exitcond3_612 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_433_inst
    process(conv79_415) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv79_415, type_cast_432_wire_constant, tmp_var);
      shr_434 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_675_inst
    process(sub_666) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_666, type_cast_674_wire_constant, tmp_var);
      shr162_676 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_685_inst
    process(sub_666) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_666, type_cast_684_wire_constant, tmp_var);
      shr168_686 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_695_inst
    process(sub_666) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_666, type_cast_694_wire_constant, tmp_var);
      shr174_696 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_705_inst
    process(sub_666) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_666, type_cast_704_wire_constant, tmp_var);
      shr180_706 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_715_inst
    process(sub_666) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_666, type_cast_714_wire_constant, tmp_var);
      shr186_716 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_725_inst
    process(sub_666) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_666, type_cast_724_wire_constant, tmp_var);
      shr192_726 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_735_inst
    process(sub_666) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_666, type_cast_734_wire_constant, tmp_var);
      shr198_736 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_769_inst
    process(add60_364, add51_339) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add60_364, add51_339, tmp_var);
      mul223_770 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_774_inst
    process(mul223_770, add69_389) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul223_770, add69_389, tmp_var);
      mul226_775 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_399_inst
    process(mul_395, add32_286) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_395, add32_286, tmp_var);
      mul78_400 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_404_inst
    process(mul78_400, add41_311) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul78_400, add41_311, tmp_var);
      sext_405 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_338_inst
    process(shl48_327, conv50_334) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl48_327, conv50_334, tmp_var);
      add51_339 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_363_inst
    process(shl57_352, conv59_359) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl57_352, conv59_359, tmp_var);
      add60_364 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_388_inst
    process(shl66_377, conv68_384) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl66_377, conv68_384, tmp_var);
      add69_389 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_260_inst
    process(shl20_249, conv22_256) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl20_249, conv22_256, tmp_var);
      add23_261 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_285_inst
    process(shl29_274, conv31_281) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl29_274, conv31_281, tmp_var);
      add32_286 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_310_inst
    process(shl38_299, conv40_306) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl38_299, conv40_306, tmp_var);
      add41_311 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_488_inst
    process(shl88_477, conv91_484) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl88_477, conv91_484, tmp_var);
      add92_489 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_506_inst
    process(shl94_495, conv97_502) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl94_495, conv97_502, tmp_var);
      add98_507 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_524_inst
    process(shl100_513, conv103_520) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl100_513, conv103_520, tmp_var);
      add104_525 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_542_inst
    process(shl106_531, conv109_538) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl106_531, conv109_538, tmp_var);
      add110_543 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_560_inst
    process(shl112_549, conv115_556) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl112_549, conv115_556, tmp_var);
      add116_561 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_578_inst
    process(shl118_567, conv121_574) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl118_567, conv121_574, tmp_var);
      add122_579 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_596_inst
    process(shl124_585, conv127_592) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl124_585, conv127_592, tmp_var);
      add128_597 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_326_inst
    process(conv47_321) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv47_321, type_cast_325_wire_constant, tmp_var);
      shl48_327 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_351_inst
    process(conv56_346) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv56_346, type_cast_350_wire_constant, tmp_var);
      shl57_352 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_376_inst
    process(conv65_371) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv65_371, type_cast_375_wire_constant, tmp_var);
      shl66_377 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_248_inst
    process(conv19_243) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv19_243, type_cast_247_wire_constant, tmp_var);
      shl20_249 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_273_inst
    process(conv28_268) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv28_268, type_cast_272_wire_constant, tmp_var);
      shl29_274 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_298_inst
    process(conv37_293) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv37_293, type_cast_297_wire_constant, tmp_var);
      shl38_299 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_394_inst
    process(add23_261) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add23_261, type_cast_393_wire_constant, tmp_var);
      mul_395 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_476_inst
    process(conv86_471) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv86_471, type_cast_475_wire_constant, tmp_var);
      shl88_477 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_494_inst
    process(add92_489) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add92_489, type_cast_493_wire_constant, tmp_var);
      shl94_495 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_512_inst
    process(add98_507) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add98_507, type_cast_511_wire_constant, tmp_var);
      shl100_513 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_530_inst
    process(add104_525) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add104_525, type_cast_529_wire_constant, tmp_var);
      shl106_531 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_548_inst
    process(add110_543) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add110_543, type_cast_547_wire_constant, tmp_var);
      shl112_549 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_566_inst
    process(add116_561) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add116_561, type_cast_565_wire_constant, tmp_var);
      shl118_567 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_584_inst
    process(add122_579) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add122_579, type_cast_583_wire_constant, tmp_var);
      shl124_585 <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_665_inst
    process(conv153_661, conv134_629) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv153_661, conv134_629, tmp_var);
      sub_666 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_420_inst
    process(conv79_415) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(conv79_415, type_cast_419_wire_constant, tmp_var);
      cmp229_421 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_439_inst
    process(shr_434) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(shr_434, type_cast_438_wire_constant, tmp_var);
      tmp1_440 <= tmp_var; --
    end process;
    -- shared split operator group (45) : array_obj_ref_462_index_offset 
    ApIntAdd_group_45: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_461_scaled;
      array_obj_ref_462_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_462_index_offset_req_0;
      array_obj_ref_462_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_462_index_offset_req_1;
      array_obj_ref_462_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_45_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_45_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_45",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 45
    -- unary operator type_cast_627_inst
    process(call133_624) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call133_624, tmp_var);
      type_cast_627_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_659_inst
    process(call152_656) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call152_656, tmp_var);
      type_cast_659_wire <= tmp_var; -- 
    end process;
    -- shared store operator group (0) : ptr_deref_599_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_599_store_0_req_0;
      ptr_deref_599_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_599_store_0_req_1;
      ptr_deref_599_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_599_word_address_0;
      data_in <= ptr_deref_599_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(13 downto 0),
          mdata => memory_space_1_sr_data(63 downto 0),
          mtag => memory_space_1_sr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block0_complete_652_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(7 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block0_complete_652_inst_req_0;
      RPIPE_Block0_complete_652_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block0_complete_652_inst_req_1;
      RPIPE_Block0_complete_652_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call149_653 <= data_out(7 downto 0);
      Block0_complete_read_0_gI: SplitGuardInterface generic map(name => "Block0_complete_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block0_complete_read_0: InputPortRevised -- 
        generic map ( name => "Block0_complete_read_0", data_width => 8,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block0_complete_pipe_read_req(0),
          oack => Block0_complete_pipe_read_ack(0),
          odata => Block0_complete_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_zeropad_input_pipe_587_inst RPIPE_zeropad_input_pipe_569_inst RPIPE_zeropad_input_pipe_551_inst RPIPE_zeropad_input_pipe_533_inst RPIPE_zeropad_input_pipe_515_inst RPIPE_zeropad_input_pipe_226_inst RPIPE_zeropad_input_pipe_229_inst RPIPE_zeropad_input_pipe_497_inst RPIPE_zeropad_input_pipe_232_inst RPIPE_zeropad_input_pipe_235_inst RPIPE_zeropad_input_pipe_479_inst RPIPE_zeropad_input_pipe_238_inst RPIPE_zeropad_input_pipe_466_inst RPIPE_zeropad_input_pipe_251_inst RPIPE_zeropad_input_pipe_263_inst RPIPE_zeropad_input_pipe_276_inst RPIPE_zeropad_input_pipe_288_inst RPIPE_zeropad_input_pipe_379_inst RPIPE_zeropad_input_pipe_301_inst RPIPE_zeropad_input_pipe_366_inst RPIPE_zeropad_input_pipe_313_inst RPIPE_zeropad_input_pipe_316_inst RPIPE_zeropad_input_pipe_354_inst RPIPE_zeropad_input_pipe_329_inst RPIPE_zeropad_input_pipe_341_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(199 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 24 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 24 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 24 downto 0);
      signal guard_vector : std_logic_vector( 24 downto 0);
      constant outBUFs : IntegerArray(24 downto 0) := (24 => 1, 23 => 1, 22 => 1, 21 => 1, 20 => 1, 19 => 1, 18 => 1, 17 => 1, 16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(24 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false, 17 => false, 18 => false, 19 => false, 20 => false, 21 => false, 22 => false, 23 => false, 24 => false);
      constant guardBuffering: IntegerArray(24 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2, 17 => 2, 18 => 2, 19 => 2, 20 => 2, 21 => 2, 22 => 2, 23 => 2, 24 => 2);
      -- 
    begin -- 
      reqL_unguarded(24) <= RPIPE_zeropad_input_pipe_587_inst_req_0;
      reqL_unguarded(23) <= RPIPE_zeropad_input_pipe_569_inst_req_0;
      reqL_unguarded(22) <= RPIPE_zeropad_input_pipe_551_inst_req_0;
      reqL_unguarded(21) <= RPIPE_zeropad_input_pipe_533_inst_req_0;
      reqL_unguarded(20) <= RPIPE_zeropad_input_pipe_515_inst_req_0;
      reqL_unguarded(19) <= RPIPE_zeropad_input_pipe_226_inst_req_0;
      reqL_unguarded(18) <= RPIPE_zeropad_input_pipe_229_inst_req_0;
      reqL_unguarded(17) <= RPIPE_zeropad_input_pipe_497_inst_req_0;
      reqL_unguarded(16) <= RPIPE_zeropad_input_pipe_232_inst_req_0;
      reqL_unguarded(15) <= RPIPE_zeropad_input_pipe_235_inst_req_0;
      reqL_unguarded(14) <= RPIPE_zeropad_input_pipe_479_inst_req_0;
      reqL_unguarded(13) <= RPIPE_zeropad_input_pipe_238_inst_req_0;
      reqL_unguarded(12) <= RPIPE_zeropad_input_pipe_466_inst_req_0;
      reqL_unguarded(11) <= RPIPE_zeropad_input_pipe_251_inst_req_0;
      reqL_unguarded(10) <= RPIPE_zeropad_input_pipe_263_inst_req_0;
      reqL_unguarded(9) <= RPIPE_zeropad_input_pipe_276_inst_req_0;
      reqL_unguarded(8) <= RPIPE_zeropad_input_pipe_288_inst_req_0;
      reqL_unguarded(7) <= RPIPE_zeropad_input_pipe_379_inst_req_0;
      reqL_unguarded(6) <= RPIPE_zeropad_input_pipe_301_inst_req_0;
      reqL_unguarded(5) <= RPIPE_zeropad_input_pipe_366_inst_req_0;
      reqL_unguarded(4) <= RPIPE_zeropad_input_pipe_313_inst_req_0;
      reqL_unguarded(3) <= RPIPE_zeropad_input_pipe_316_inst_req_0;
      reqL_unguarded(2) <= RPIPE_zeropad_input_pipe_354_inst_req_0;
      reqL_unguarded(1) <= RPIPE_zeropad_input_pipe_329_inst_req_0;
      reqL_unguarded(0) <= RPIPE_zeropad_input_pipe_341_inst_req_0;
      RPIPE_zeropad_input_pipe_587_inst_ack_0 <= ackL_unguarded(24);
      RPIPE_zeropad_input_pipe_569_inst_ack_0 <= ackL_unguarded(23);
      RPIPE_zeropad_input_pipe_551_inst_ack_0 <= ackL_unguarded(22);
      RPIPE_zeropad_input_pipe_533_inst_ack_0 <= ackL_unguarded(21);
      RPIPE_zeropad_input_pipe_515_inst_ack_0 <= ackL_unguarded(20);
      RPIPE_zeropad_input_pipe_226_inst_ack_0 <= ackL_unguarded(19);
      RPIPE_zeropad_input_pipe_229_inst_ack_0 <= ackL_unguarded(18);
      RPIPE_zeropad_input_pipe_497_inst_ack_0 <= ackL_unguarded(17);
      RPIPE_zeropad_input_pipe_232_inst_ack_0 <= ackL_unguarded(16);
      RPIPE_zeropad_input_pipe_235_inst_ack_0 <= ackL_unguarded(15);
      RPIPE_zeropad_input_pipe_479_inst_ack_0 <= ackL_unguarded(14);
      RPIPE_zeropad_input_pipe_238_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_zeropad_input_pipe_466_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_zeropad_input_pipe_251_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_zeropad_input_pipe_263_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_zeropad_input_pipe_276_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_zeropad_input_pipe_288_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_zeropad_input_pipe_379_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_zeropad_input_pipe_301_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_zeropad_input_pipe_366_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_zeropad_input_pipe_313_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_zeropad_input_pipe_316_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_zeropad_input_pipe_354_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_zeropad_input_pipe_329_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_zeropad_input_pipe_341_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(24) <= RPIPE_zeropad_input_pipe_587_inst_req_1;
      reqR_unguarded(23) <= RPIPE_zeropad_input_pipe_569_inst_req_1;
      reqR_unguarded(22) <= RPIPE_zeropad_input_pipe_551_inst_req_1;
      reqR_unguarded(21) <= RPIPE_zeropad_input_pipe_533_inst_req_1;
      reqR_unguarded(20) <= RPIPE_zeropad_input_pipe_515_inst_req_1;
      reqR_unguarded(19) <= RPIPE_zeropad_input_pipe_226_inst_req_1;
      reqR_unguarded(18) <= RPIPE_zeropad_input_pipe_229_inst_req_1;
      reqR_unguarded(17) <= RPIPE_zeropad_input_pipe_497_inst_req_1;
      reqR_unguarded(16) <= RPIPE_zeropad_input_pipe_232_inst_req_1;
      reqR_unguarded(15) <= RPIPE_zeropad_input_pipe_235_inst_req_1;
      reqR_unguarded(14) <= RPIPE_zeropad_input_pipe_479_inst_req_1;
      reqR_unguarded(13) <= RPIPE_zeropad_input_pipe_238_inst_req_1;
      reqR_unguarded(12) <= RPIPE_zeropad_input_pipe_466_inst_req_1;
      reqR_unguarded(11) <= RPIPE_zeropad_input_pipe_251_inst_req_1;
      reqR_unguarded(10) <= RPIPE_zeropad_input_pipe_263_inst_req_1;
      reqR_unguarded(9) <= RPIPE_zeropad_input_pipe_276_inst_req_1;
      reqR_unguarded(8) <= RPIPE_zeropad_input_pipe_288_inst_req_1;
      reqR_unguarded(7) <= RPIPE_zeropad_input_pipe_379_inst_req_1;
      reqR_unguarded(6) <= RPIPE_zeropad_input_pipe_301_inst_req_1;
      reqR_unguarded(5) <= RPIPE_zeropad_input_pipe_366_inst_req_1;
      reqR_unguarded(4) <= RPIPE_zeropad_input_pipe_313_inst_req_1;
      reqR_unguarded(3) <= RPIPE_zeropad_input_pipe_316_inst_req_1;
      reqR_unguarded(2) <= RPIPE_zeropad_input_pipe_354_inst_req_1;
      reqR_unguarded(1) <= RPIPE_zeropad_input_pipe_329_inst_req_1;
      reqR_unguarded(0) <= RPIPE_zeropad_input_pipe_341_inst_req_1;
      RPIPE_zeropad_input_pipe_587_inst_ack_1 <= ackR_unguarded(24);
      RPIPE_zeropad_input_pipe_569_inst_ack_1 <= ackR_unguarded(23);
      RPIPE_zeropad_input_pipe_551_inst_ack_1 <= ackR_unguarded(22);
      RPIPE_zeropad_input_pipe_533_inst_ack_1 <= ackR_unguarded(21);
      RPIPE_zeropad_input_pipe_515_inst_ack_1 <= ackR_unguarded(20);
      RPIPE_zeropad_input_pipe_226_inst_ack_1 <= ackR_unguarded(19);
      RPIPE_zeropad_input_pipe_229_inst_ack_1 <= ackR_unguarded(18);
      RPIPE_zeropad_input_pipe_497_inst_ack_1 <= ackR_unguarded(17);
      RPIPE_zeropad_input_pipe_232_inst_ack_1 <= ackR_unguarded(16);
      RPIPE_zeropad_input_pipe_235_inst_ack_1 <= ackR_unguarded(15);
      RPIPE_zeropad_input_pipe_479_inst_ack_1 <= ackR_unguarded(14);
      RPIPE_zeropad_input_pipe_238_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_zeropad_input_pipe_466_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_zeropad_input_pipe_251_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_zeropad_input_pipe_263_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_zeropad_input_pipe_276_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_zeropad_input_pipe_288_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_zeropad_input_pipe_379_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_zeropad_input_pipe_301_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_zeropad_input_pipe_366_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_zeropad_input_pipe_313_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_zeropad_input_pipe_316_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_zeropad_input_pipe_354_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_zeropad_input_pipe_329_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_zeropad_input_pipe_341_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      guard_vector(18)  <=  '1';
      guard_vector(19)  <=  '1';
      guard_vector(20)  <=  '1';
      guard_vector(21)  <=  '1';
      guard_vector(22)  <=  '1';
      guard_vector(23)  <=  '1';
      guard_vector(24)  <=  '1';
      call125_588 <= data_out(199 downto 192);
      call119_570 <= data_out(191 downto 184);
      call113_552 <= data_out(183 downto 176);
      call107_534 <= data_out(175 downto 168);
      call101_516 <= data_out(167 downto 160);
      call_227 <= data_out(159 downto 152);
      call2_230 <= data_out(151 downto 144);
      call95_498 <= data_out(143 downto 136);
      call6_233 <= data_out(135 downto 128);
      call11_236 <= data_out(127 downto 120);
      call89_480 <= data_out(119 downto 112);
      call16_239 <= data_out(111 downto 104);
      call85_467 <= data_out(103 downto 96);
      call21_252 <= data_out(95 downto 88);
      call25_264 <= data_out(87 downto 80);
      call30_277 <= data_out(79 downto 72);
      call34_289 <= data_out(71 downto 64);
      call67_380 <= data_out(63 downto 56);
      call39_302 <= data_out(55 downto 48);
      call62_367 <= data_out(47 downto 40);
      call43_314 <= data_out(39 downto 32);
      call44_317 <= data_out(31 downto 24);
      call58_355 <= data_out(23 downto 16);
      call49_330 <= data_out(15 downto 8);
      call53_342 <= data_out(7 downto 0);
      zeropad_input_pipe_read_1_gI: SplitGuardInterface generic map(name => "zeropad_input_pipe_read_1_gI", nreqs => 25, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      zeropad_input_pipe_read_1: InputPortRevised -- 
        generic map ( name => "zeropad_input_pipe_read_1", data_width => 8,  num_reqs => 25,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => zeropad_input_pipe_pipe_read_req(0),
          oack => zeropad_input_pipe_pipe_read_ack(0),
          odata => zeropad_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared outport operator group (0) : WPIPE_Block0_starting_633_inst WPIPE_Block0_starting_630_inst WPIPE_Block0_starting_636_inst WPIPE_Block0_starting_639_inst WPIPE_Block0_starting_642_inst WPIPE_Block0_starting_645_inst WPIPE_Block0_starting_648_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(55 downto 0);
      signal sample_req, sample_ack : BooleanArray( 6 downto 0);
      signal update_req, update_ack : BooleanArray( 6 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 6 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 6 downto 0);
      signal guard_vector : std_logic_vector( 6 downto 0);
      constant inBUFs : IntegerArray(6 downto 0) := (6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(6 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false);
      constant guardBuffering: IntegerArray(6 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2);
      -- 
    begin -- 
      sample_req_unguarded(6) <= WPIPE_Block0_starting_633_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Block0_starting_630_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Block0_starting_636_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Block0_starting_639_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Block0_starting_642_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Block0_starting_645_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Block0_starting_648_inst_req_0;
      WPIPE_Block0_starting_633_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Block0_starting_630_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Block0_starting_636_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Block0_starting_639_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Block0_starting_642_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Block0_starting_645_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Block0_starting_648_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(6) <= WPIPE_Block0_starting_633_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Block0_starting_630_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Block0_starting_636_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Block0_starting_639_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Block0_starting_642_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Block0_starting_645_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Block0_starting_648_inst_req_1;
      WPIPE_Block0_starting_633_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Block0_starting_630_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Block0_starting_636_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Block0_starting_639_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Block0_starting_642_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Block0_starting_645_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Block0_starting_648_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      data_in <= call30_277 & call21_252 & call39_302 & call49_330 & call58_355 & call67_380 & call43_314;
      Block0_starting_write_0_gI: SplitGuardInterface generic map(name => "Block0_starting_write_0_gI", nreqs => 7, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block0_starting_write_0: OutputPortRevised -- 
        generic map ( name => "Block0_starting", data_width => 8, num_reqs => 7, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block0_starting_pipe_write_req(0),
          oack => Block0_starting_pipe_write_ack(0),
          odata => Block0_starting_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_zeropad_output_pipe_741_inst WPIPE_zeropad_output_pipe_750_inst WPIPE_zeropad_output_pipe_759_inst WPIPE_zeropad_output_pipe_744_inst WPIPE_zeropad_output_pipe_753_inst WPIPE_zeropad_output_pipe_756_inst WPIPE_zeropad_output_pipe_747_inst WPIPE_zeropad_output_pipe_762_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 7 downto 0);
      signal update_req, update_ack : BooleanArray( 7 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 7 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 7 downto 0);
      signal guard_vector : std_logic_vector( 7 downto 0);
      constant inBUFs : IntegerArray(7 downto 0) := (7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(7 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false);
      constant guardBuffering: IntegerArray(7 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2);
      -- 
    begin -- 
      sample_req_unguarded(7) <= WPIPE_zeropad_output_pipe_741_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_zeropad_output_pipe_750_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_zeropad_output_pipe_759_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_zeropad_output_pipe_744_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_zeropad_output_pipe_753_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_zeropad_output_pipe_756_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_zeropad_output_pipe_747_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_zeropad_output_pipe_762_inst_req_0;
      WPIPE_zeropad_output_pipe_741_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_zeropad_output_pipe_750_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_zeropad_output_pipe_759_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_zeropad_output_pipe_744_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_zeropad_output_pipe_753_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_zeropad_output_pipe_756_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_zeropad_output_pipe_747_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_zeropad_output_pipe_762_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(7) <= WPIPE_zeropad_output_pipe_741_inst_req_1;
      update_req_unguarded(6) <= WPIPE_zeropad_output_pipe_750_inst_req_1;
      update_req_unguarded(5) <= WPIPE_zeropad_output_pipe_759_inst_req_1;
      update_req_unguarded(4) <= WPIPE_zeropad_output_pipe_744_inst_req_1;
      update_req_unguarded(3) <= WPIPE_zeropad_output_pipe_753_inst_req_1;
      update_req_unguarded(2) <= WPIPE_zeropad_output_pipe_756_inst_req_1;
      update_req_unguarded(1) <= WPIPE_zeropad_output_pipe_747_inst_req_1;
      update_req_unguarded(0) <= WPIPE_zeropad_output_pipe_762_inst_req_1;
      WPIPE_zeropad_output_pipe_741_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_zeropad_output_pipe_750_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_zeropad_output_pipe_759_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_zeropad_output_pipe_744_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_zeropad_output_pipe_753_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_zeropad_output_pipe_756_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_zeropad_output_pipe_747_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_zeropad_output_pipe_762_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      data_in <= conv201_740 & conv183_710 & conv165_680 & conv195_730 & conv177_700 & conv171_690 & conv189_720 & conv159_670;
      zeropad_output_pipe_write_1_gI: SplitGuardInterface generic map(name => "zeropad_output_pipe_write_1_gI", nreqs => 8, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      zeropad_output_pipe_write_1: OutputPortRevised -- 
        generic map ( name => "zeropad_output_pipe", data_width => 8, num_reqs => 8, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => zeropad_output_pipe_pipe_write_req(0),
          oack => zeropad_output_pipe_pipe_write_ack(0),
          odata => zeropad_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared call operator group (0) : call_stmt_656_call call_stmt_624_call 
    timer_call_group_0: Block -- 
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_656_call_req_0;
      reqL_unguarded(0) <= call_stmt_624_call_req_0;
      call_stmt_656_call_ack_0 <= ackL_unguarded(1);
      call_stmt_624_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_656_call_req_1;
      reqR_unguarded(0) <= call_stmt_624_call_req_1;
      call_stmt_656_call_ack_1 <= ackR_unguarded(1);
      call_stmt_624_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      timer_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      timer_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      timer_call_group_0_gI: SplitGuardInterface generic map(name => "timer_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      call152_656 <= data_out(127 downto 64);
      call133_624 <= data_out(63 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 2,
        nreqs => 2,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => timer_call_reqs(0),
          ackR => timer_call_acks(0),
          tagR => timer_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => timer_return_acks(0), -- cross-over
          ackL => timer_return_reqs(0), -- cross-over
          dataL => timer_return_data(63 downto 0),
          tagL => timer_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_777_call 
    sendOutput_call_group_1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_777_call_req_0;
      call_stmt_777_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_777_call_req_1;
      call_stmt_777_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      sendOutput_call_group_1_gI: SplitGuardInterface generic map(name => "sendOutput_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= mul226_775;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 32,
        owidth => 32,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => sendOutput_call_reqs(0),
          ackR => sendOutput_call_acks(0),
          dataR => sendOutput_call_data(31 downto 0),
          tagR => sendOutput_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => sendOutput_return_acks(0), -- cross-over
          ackL => sendOutput_return_reqs(0), -- cross-over
          tagL => sendOutput_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- 
  end Block; -- data_path
  -- 
end zeropad3D_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity zeropad3D_A is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
    Block0_starting_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block0_starting_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block0_starting_pipe_read_data : in   std_logic_vector(7 downto 0);
    Block0_complete_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block0_complete_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block0_complete_pipe_write_data : out  std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity zeropad3D_A;
architecture zeropad3D_A_arch of zeropad3D_A is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal zeropad3D_A_CP_1983_start: Boolean;
  signal zeropad3D_A_CP_1983_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal phi_stmt_915_req_1 : boolean;
  signal phi_stmt_910_req_1 : boolean;
  signal type_cast_923_inst_ack_0 : boolean;
  signal phi_stmt_905_req_0 : boolean;
  signal type_cast_854_inst_ack_1 : boolean;
  signal type_cast_868_inst_ack_1 : boolean;
  signal W_ifx_xthen_ifx_xend80_taken_1078_delayed_3_0_1149_inst_req_1 : boolean;
  signal W_ifx_xend80_exec_guard_1189_delayed_1_0_1278_inst_ack_0 : boolean;
  signal type_cast_854_inst_req_1 : boolean;
  signal type_cast_918_inst_ack_1 : boolean;
  signal phi_stmt_915_ack_0 : boolean;
  signal phi_stmt_910_ack_0 : boolean;
  signal phi_stmt_915_req_0 : boolean;
  signal W_ifx_xend80_exec_guard_1161_delayed_1_0_1236_inst_req_0 : boolean;
  signal W_kx_x1_944_delayed_1_0_945_inst_ack_0 : boolean;
  signal W_kx_x1_944_delayed_1_0_945_inst_req_0 : boolean;
  signal W_jx_x1_957_delayed_1_0_961_inst_ack_0 : boolean;
  signal type_cast_913_inst_ack_1 : boolean;
  signal W_jx_x1_957_delayed_1_0_961_inst_req_0 : boolean;
  signal type_cast_854_inst_ack_0 : boolean;
  signal type_cast_913_inst_req_1 : boolean;
  signal type_cast_854_inst_req_0 : boolean;
  signal W_kx_x1_944_delayed_1_0_945_inst_req_1 : boolean;
  signal W_kx_x1_944_delayed_1_0_945_inst_ack_1 : boolean;
  signal type_cast_908_inst_ack_1 : boolean;
  signal type_cast_923_inst_req_1 : boolean;
  signal type_cast_923_inst_ack_1 : boolean;
  signal type_cast_1304_inst_ack_0 : boolean;
  signal type_cast_1260_inst_req_0 : boolean;
  signal W_ifx_xelse_exec_guard_973_delayed_1_0_985_inst_req_0 : boolean;
  signal type_cast_1260_inst_req_1 : boolean;
  signal type_cast_913_inst_ack_0 : boolean;
  signal type_cast_974_inst_req_0 : boolean;
  signal W_ifx_xelse_exec_guard_978_delayed_2_0_993_inst_req_0 : boolean;
  signal type_cast_1304_inst_req_0 : boolean;
  signal type_cast_868_inst_ack_0 : boolean;
  signal W_ifx_xelse_exec_guard_967_delayed_1_0_976_inst_ack_0 : boolean;
  signal W_ifx_xelse_exec_guard_978_delayed_2_0_993_inst_ack_1 : boolean;
  signal type_cast_1330_inst_req_0 : boolean;
  signal type_cast_991_inst_ack_1 : boolean;
  signal W_ifx_xelse_exec_guard_978_delayed_2_0_993_inst_req_1 : boolean;
  signal W_ifx_xelse_exec_guard_973_delayed_1_0_985_inst_ack_0 : boolean;
  signal addr_of_1502_final_reg_ack_0 : boolean;
  signal type_cast_974_inst_ack_0 : boolean;
  signal W_ifx_xelse_exec_guard_973_delayed_1_0_985_inst_req_1 : boolean;
  signal W_ifx_xelse_exec_guard_973_delayed_1_0_985_inst_ack_1 : boolean;
  signal W_jx_x1_957_delayed_1_0_961_inst_req_1 : boolean;
  signal type_cast_918_inst_req_0 : boolean;
  signal W_ifx_xend80_exec_guard_1189_delayed_1_0_1278_inst_req_0 : boolean;
  signal type_cast_918_inst_ack_0 : boolean;
  signal W_ifx_xelse_exec_guard_967_delayed_1_0_976_inst_req_0 : boolean;
  signal W_ifx_xthen_ifx_xend80_taken_1078_delayed_3_0_1149_inst_ack_0 : boolean;
  signal type_cast_908_inst_req_0 : boolean;
  signal W_ifx_xthen_ifx_xend80_taken_1078_delayed_3_0_1149_inst_req_0 : boolean;
  signal type_cast_839_inst_ack_1 : boolean;
  signal phi_stmt_905_ack_0 : boolean;
  signal type_cast_868_inst_req_0 : boolean;
  signal W_lorx_xlhsx_xfalse135_exec_guard_1240_delayed_1_0_1356_inst_ack_0 : boolean;
  signal type_cast_908_inst_ack_0 : boolean;
  signal type_cast_913_inst_req_0 : boolean;
  signal W_ifx_xend80_exec_guard_1167_delayed_1_0_1245_inst_req_0 : boolean;
  signal W_jx_x1_957_delayed_1_0_961_inst_ack_1 : boolean;
  signal type_cast_839_inst_req_1 : boolean;
  signal type_cast_1234_inst_req_0 : boolean;
  signal W_ifx_xelse_exec_guard_967_delayed_1_0_976_inst_req_1 : boolean;
  signal W_ifx_xelse_exec_guard_967_delayed_1_0_976_inst_ack_1 : boolean;
  signal type_cast_908_inst_req_1 : boolean;
  signal type_cast_991_inst_req_0 : boolean;
  signal type_cast_991_inst_ack_0 : boolean;
  signal type_cast_991_inst_req_1 : boolean;
  signal phi_stmt_910_req_0 : boolean;
  signal W_add96_1252_delayed_2_0_1373_inst_ack_0 : boolean;
  signal type_cast_974_inst_req_1 : boolean;
  signal type_cast_923_inst_req_0 : boolean;
  signal W_ifx_xelse_exec_guard_978_delayed_2_0_993_inst_ack_0 : boolean;
  signal type_cast_868_inst_req_1 : boolean;
  signal type_cast_1260_inst_ack_1 : boolean;
  signal type_cast_1234_inst_ack_0 : boolean;
  signal type_cast_918_inst_req_1 : boolean;
  signal type_cast_1260_inst_ack_0 : boolean;
  signal W_ifx_xend80_exec_guard_1167_delayed_1_0_1245_inst_ack_0 : boolean;
  signal phi_stmt_905_req_1 : boolean;
  signal type_cast_974_inst_ack_1 : boolean;
  signal W_lorx_xlhsx_xfalse135_exec_guard_1220_delayed_1_0_1325_inst_req_1 : boolean;
  signal W_ifx_xend80_exec_guard_1161_delayed_1_0_1236_inst_ack_0 : boolean;
  signal W_lorx_xlhsx_xfalse135_exec_guard_1220_delayed_1_0_1325_inst_ack_1 : boolean;
  signal type_cast_1330_inst_ack_0 : boolean;
  signal W_ifx_xthen_ifx_xend80_taken_1078_delayed_3_0_1149_inst_ack_1 : boolean;
  signal type_cast_927_inst_ack_1 : boolean;
  signal type_cast_927_inst_req_1 : boolean;
  signal W_ifx_xelse155_exec_guard_1328_delayed_1_0_1475_inst_ack_1 : boolean;
  signal type_cast_927_inst_ack_0 : boolean;
  signal type_cast_927_inst_req_0 : boolean;
  signal do_while_stmt_903_branch_req_0 : boolean;
  signal type_cast_1495_inst_ack_0 : boolean;
  signal if_stmt_1527_branch_ack_0 : boolean;
  signal type_cast_1234_inst_req_1 : boolean;
  signal type_cast_1330_inst_req_1 : boolean;
  signal addr_of_1502_final_reg_req_0 : boolean;
  signal type_cast_1234_inst_ack_1 : boolean;
  signal RPIPE_Block0_starting_785_inst_req_0 : boolean;
  signal RPIPE_Block0_starting_785_inst_ack_0 : boolean;
  signal type_cast_1304_inst_req_1 : boolean;
  signal RPIPE_Block0_starting_785_inst_req_1 : boolean;
  signal RPIPE_Block0_starting_785_inst_ack_1 : boolean;
  signal W_ifx_xend80_exec_guard_1161_delayed_1_0_1236_inst_req_1 : boolean;
  signal W_add96_1324_delayed_2_0_1466_inst_req_0 : boolean;
  signal type_cast_1304_inst_ack_1 : boolean;
  signal RPIPE_Block0_starting_788_inst_req_0 : boolean;
  signal RPIPE_Block0_starting_788_inst_ack_0 : boolean;
  signal W_ifx_xend80_exec_guard_1161_delayed_1_0_1236_inst_ack_1 : boolean;
  signal RPIPE_Block0_starting_788_inst_req_1 : boolean;
  signal RPIPE_Block0_starting_788_inst_ack_1 : boolean;
  signal RPIPE_Block0_starting_791_inst_req_0 : boolean;
  signal RPIPE_Block0_starting_791_inst_ack_0 : boolean;
  signal RPIPE_Block0_starting_791_inst_req_1 : boolean;
  signal RPIPE_Block0_starting_791_inst_ack_1 : boolean;
  signal W_ifx_xend80_exec_guard_1182_delayed_1_0_1269_inst_req_0 : boolean;
  signal RPIPE_Block0_starting_794_inst_req_0 : boolean;
  signal RPIPE_Block0_starting_794_inst_ack_0 : boolean;
  signal RPIPE_Block0_starting_794_inst_req_1 : boolean;
  signal RPIPE_Block0_starting_794_inst_ack_1 : boolean;
  signal W_ifx_xend80_exec_guard_1182_delayed_1_0_1269_inst_ack_0 : boolean;
  signal W_ifx_xend80_exec_guard_1189_delayed_1_0_1278_inst_req_1 : boolean;
  signal RPIPE_Block0_starting_797_inst_req_0 : boolean;
  signal RPIPE_Block0_starting_797_inst_ack_0 : boolean;
  signal RPIPE_Block0_starting_797_inst_req_1 : boolean;
  signal RPIPE_Block0_starting_797_inst_ack_1 : boolean;
  signal W_ifx_xend80_exec_guard_1182_delayed_1_0_1269_inst_req_1 : boolean;
  signal RPIPE_Block0_starting_800_inst_req_0 : boolean;
  signal RPIPE_Block0_starting_800_inst_ack_0 : boolean;
  signal RPIPE_Block0_starting_800_inst_req_1 : boolean;
  signal RPIPE_Block0_starting_800_inst_ack_1 : boolean;
  signal RPIPE_Block0_starting_803_inst_req_0 : boolean;
  signal RPIPE_Block0_starting_803_inst_ack_0 : boolean;
  signal RPIPE_Block0_starting_803_inst_req_1 : boolean;
  signal RPIPE_Block0_starting_803_inst_ack_1 : boolean;
  signal type_cast_809_inst_req_0 : boolean;
  signal type_cast_809_inst_ack_0 : boolean;
  signal type_cast_809_inst_req_1 : boolean;
  signal type_cast_809_inst_ack_1 : boolean;
  signal type_cast_813_inst_req_0 : boolean;
  signal type_cast_813_inst_ack_0 : boolean;
  signal type_cast_813_inst_req_1 : boolean;
  signal type_cast_813_inst_ack_1 : boolean;
  signal type_cast_817_inst_req_0 : boolean;
  signal type_cast_817_inst_ack_0 : boolean;
  signal type_cast_817_inst_req_1 : boolean;
  signal type_cast_817_inst_ack_1 : boolean;
  signal type_cast_821_inst_req_0 : boolean;
  signal type_cast_821_inst_ack_0 : boolean;
  signal type_cast_821_inst_req_1 : boolean;
  signal type_cast_821_inst_ack_1 : boolean;
  signal type_cast_825_inst_req_0 : boolean;
  signal type_cast_825_inst_ack_0 : boolean;
  signal type_cast_825_inst_req_1 : boolean;
  signal type_cast_825_inst_ack_1 : boolean;
  signal type_cast_835_inst_req_0 : boolean;
  signal type_cast_835_inst_ack_0 : boolean;
  signal type_cast_835_inst_req_1 : boolean;
  signal type_cast_835_inst_ack_1 : boolean;
  signal type_cast_839_inst_req_0 : boolean;
  signal type_cast_839_inst_ack_0 : boolean;
  signal W_ix_x2_981_delayed_3_0_996_inst_req_0 : boolean;
  signal W_ix_x2_981_delayed_3_0_996_inst_ack_0 : boolean;
  signal W_ix_x2_981_delayed_3_0_996_inst_req_1 : boolean;
  signal W_ix_x2_981_delayed_3_0_996_inst_ack_1 : boolean;
  signal ptr_deref_1512_store_0_ack_0 : boolean;
  signal W_add96_1252_delayed_2_0_1373_inst_ack_1 : boolean;
  signal W_ifx_xelse_exec_guard_984_delayed_1_0_1005_inst_req_0 : boolean;
  signal W_ifx_xelse_exec_guard_984_delayed_1_0_1005_inst_ack_0 : boolean;
  signal W_ifx_xelse_exec_guard_984_delayed_1_0_1005_inst_req_1 : boolean;
  signal W_ifx_xelse_exec_guard_984_delayed_1_0_1005_inst_ack_1 : boolean;
  signal W_add96_1252_delayed_2_0_1373_inst_req_1 : boolean;
  signal W_add96_1252_delayed_2_0_1373_inst_req_0 : boolean;
  signal type_cast_1380_inst_req_0 : boolean;
  signal W_lorx_xlhsx_xfalse135_exec_guard_1220_delayed_1_0_1325_inst_ack_0 : boolean;
  signal W_lorx_xlhsx_xfalse135_exec_guard_1220_delayed_1_0_1325_inst_req_0 : boolean;
  signal W_inc_989_delayed_1_0_1008_inst_req_0 : boolean;
  signal W_inc_989_delayed_1_0_1008_inst_ack_0 : boolean;
  signal W_inc_989_delayed_1_0_1008_inst_req_1 : boolean;
  signal W_inc_989_delayed_1_0_1008_inst_ack_1 : boolean;
  signal W_ifx_xelse_exec_guard_992_delayed_2_0_1019_inst_req_0 : boolean;
  signal W_ifx_xelse_exec_guard_992_delayed_2_0_1019_inst_ack_0 : boolean;
  signal W_ifx_xelse_exec_guard_992_delayed_2_0_1019_inst_req_1 : boolean;
  signal W_jx_x0_1204_delayed_1_0_1298_inst_ack_1 : boolean;
  signal W_ifx_xelse_exec_guard_992_delayed_2_0_1019_inst_ack_1 : boolean;
  signal W_ifx_xend80_ifx_xthen152_taken_1246_delayed_1_0_1365_inst_ack_1 : boolean;
  signal W_ifx_xend80_ifx_xthen152_taken_1246_delayed_1_0_1365_inst_req_1 : boolean;
  signal W_lorx_xlhsx_xfalse135_exec_guard_1228_delayed_1_0_1339_inst_ack_1 : boolean;
  signal W_jx_x0_1204_delayed_1_0_1298_inst_req_1 : boolean;
  signal W_lorx_xlhsx_xfalse135_exec_guard_1228_delayed_1_0_1339_inst_req_1 : boolean;
  signal type_cast_1025_inst_req_0 : boolean;
  signal type_cast_1025_inst_ack_0 : boolean;
  signal type_cast_1025_inst_req_1 : boolean;
  signal type_cast_1025_inst_ack_1 : boolean;
  signal W_lorx_xlhsx_xfalse135_exec_guard_1213_delayed_1_0_1315_inst_ack_1 : boolean;
  signal W_ifx_xelse_exec_guard_997_delayed_3_0_1027_inst_req_0 : boolean;
  signal W_jx_x0_1204_delayed_1_0_1298_inst_ack_0 : boolean;
  signal W_ifx_xelse_exec_guard_997_delayed_3_0_1027_inst_ack_0 : boolean;
  signal W_ifx_xelse_exec_guard_997_delayed_3_0_1027_inst_req_1 : boolean;
  signal W_jx_x0_1204_delayed_1_0_1298_inst_req_0 : boolean;
  signal W_ifx_xelse_exec_guard_997_delayed_3_0_1027_inst_ack_1 : boolean;
  signal W_lorx_xlhsx_xfalse135_exec_guard_1213_delayed_1_0_1315_inst_req_1 : boolean;
  signal W_ifx_xend80_exec_guard_1174_delayed_1_0_1255_inst_ack_1 : boolean;
  signal W_lorx_xlhsx_xfalse135_exec_guard_1228_delayed_1_0_1339_inst_ack_0 : boolean;
  signal W_ifx_xelse_exec_guard_1004_delayed_3_0_1036_inst_req_0 : boolean;
  signal W_ifx_xelse_exec_guard_1004_delayed_3_0_1036_inst_ack_0 : boolean;
  signal ptr_deref_1512_store_0_req_1 : boolean;
  signal W_lorx_xlhsx_xfalse135_exec_guard_1235_delayed_1_0_1348_inst_ack_1 : boolean;
  signal W_ifx_xelse_exec_guard_1004_delayed_3_0_1036_inst_req_1 : boolean;
  signal W_ifx_xelse_exec_guard_1004_delayed_3_0_1036_inst_ack_1 : boolean;
  signal W_lorx_xlhsx_xfalse135_exec_guard_1240_delayed_1_0_1356_inst_req_0 : boolean;
  signal W_lorx_xlhsx_xfalse135_exec_guard_1235_delayed_1_0_1348_inst_req_1 : boolean;
  signal if_stmt_1527_branch_ack_1 : boolean;
  signal W_ifx_xend80_exec_guard_1174_delayed_1_0_1255_inst_req_1 : boolean;
  signal W_lorx_xlhsx_xfalse135_exec_guard_1213_delayed_1_0_1315_inst_ack_0 : boolean;
  signal W_ifx_xelse_exec_guard_1009_delayed_3_0_1044_inst_req_0 : boolean;
  signal W_ifx_xelse_exec_guard_1009_delayed_3_0_1044_inst_ack_0 : boolean;
  signal W_lorx_xlhsx_xfalse135_exec_guard_1228_delayed_1_0_1339_inst_req_0 : boolean;
  signal W_ifx_xelse_exec_guard_1009_delayed_3_0_1044_inst_req_1 : boolean;
  signal W_ifx_xelse_exec_guard_1009_delayed_3_0_1044_inst_ack_1 : boolean;
  signal W_ifx_xend80_ifx_xthen152_taken_1246_delayed_1_0_1365_inst_ack_0 : boolean;
  signal W_lorx_xlhsx_xfalse135_exec_guard_1213_delayed_1_0_1315_inst_req_0 : boolean;
  signal W_ifx_xthen_ifx_xend80_taken_1022_delayed_3_0_1059_inst_req_0 : boolean;
  signal W_ifx_xthen_ifx_xend80_taken_1022_delayed_3_0_1059_inst_ack_0 : boolean;
  signal W_ifx_xthen_ifx_xend80_taken_1022_delayed_3_0_1059_inst_req_1 : boolean;
  signal W_ifx_xthen_ifx_xend80_taken_1022_delayed_3_0_1059_inst_ack_1 : boolean;
  signal W_ifx_xend80_ifx_xthen152_taken_1246_delayed_1_0_1365_inst_req_0 : boolean;
  signal W_lorx_xlhsx_xfalse135_exec_guard_1235_delayed_1_0_1348_inst_ack_0 : boolean;
  signal W_lorx_xlhsx_xfalse135_exec_guard_1235_delayed_1_0_1348_inst_req_0 : boolean;
  signal W_ifx_xthen_ifx_xend80_taken_1028_delayed_3_0_1069_inst_req_0 : boolean;
  signal W_ifx_xend80_exec_guard_1194_delayed_1_0_1286_inst_ack_1 : boolean;
  signal W_ifx_xthen_ifx_xend80_taken_1028_delayed_3_0_1069_inst_ack_0 : boolean;
  signal W_ifx_xthen_ifx_xend80_taken_1028_delayed_3_0_1069_inst_req_1 : boolean;
  signal W_ifx_xend80_exec_guard_1194_delayed_1_0_1286_inst_req_1 : boolean;
  signal W_ifx_xthen_ifx_xend80_taken_1028_delayed_3_0_1069_inst_ack_1 : boolean;
  signal W_ifx_xelse155_exec_guard_1328_delayed_1_0_1475_inst_req_1 : boolean;
  signal W_ifx_xend80_exec_guard_1174_delayed_1_0_1255_inst_ack_0 : boolean;
  signal type_cast_1074_inst_req_0 : boolean;
  signal type_cast_1074_inst_ack_0 : boolean;
  signal type_cast_1074_inst_req_1 : boolean;
  signal W_ifx_xend80_exec_guard_1194_delayed_1_0_1286_inst_ack_0 : boolean;
  signal type_cast_1074_inst_ack_1 : boolean;
  signal W_lorx_xlhsx_xfalse135_exec_guard_1207_delayed_1_0_1306_inst_ack_1 : boolean;
  signal type_cast_1380_inst_req_1 : boolean;
  signal type_cast_1380_inst_ack_1 : boolean;
  signal W_ifx_xend80_exec_guard_1174_delayed_1_0_1255_inst_req_0 : boolean;
  signal W_lorx_xlhsx_xfalse135_exec_guard_1207_delayed_1_0_1306_inst_req_1 : boolean;
  signal W_ifx_xthen_ifx_xend80_taken_1046_delayed_3_0_1093_inst_req_0 : boolean;
  signal W_ifx_xend80_exec_guard_1194_delayed_1_0_1286_inst_req_0 : boolean;
  signal W_ifx_xthen_ifx_xend80_taken_1046_delayed_3_0_1093_inst_ack_0 : boolean;
  signal W_ifx_xthen_ifx_xend80_taken_1046_delayed_3_0_1093_inst_req_1 : boolean;
  signal W_ifx_xthen_ifx_xend80_taken_1046_delayed_3_0_1093_inst_ack_1 : boolean;
  signal W_lorx_xlhsx_xfalse135_exec_guard_1240_delayed_1_0_1356_inst_ack_1 : boolean;
  signal type_cast_1098_inst_req_0 : boolean;
  signal type_cast_1098_inst_ack_0 : boolean;
  signal addr_of_1502_final_reg_req_1 : boolean;
  signal type_cast_1098_inst_req_1 : boolean;
  signal type_cast_1098_inst_ack_1 : boolean;
  signal W_lorx_xlhsx_xfalse135_exec_guard_1207_delayed_1_0_1306_inst_ack_0 : boolean;
  signal type_cast_1102_inst_req_0 : boolean;
  signal type_cast_1102_inst_ack_0 : boolean;
  signal type_cast_1102_inst_req_1 : boolean;
  signal type_cast_1102_inst_ack_1 : boolean;
  signal W_lorx_xlhsx_xfalse135_exec_guard_1240_delayed_1_0_1356_inst_req_1 : boolean;
  signal type_cast_1380_inst_ack_0 : boolean;
  signal W_lorx_xlhsx_xfalse135_exec_guard_1207_delayed_1_0_1306_inst_req_0 : boolean;
  signal W_ifx_xend80_exec_guard_1182_delayed_1_0_1269_inst_ack_1 : boolean;
  signal type_cast_1106_inst_req_0 : boolean;
  signal type_cast_1106_inst_ack_0 : boolean;
  signal type_cast_1106_inst_req_1 : boolean;
  signal W_ifx_xend80_exec_guard_1189_delayed_1_0_1278_inst_ack_1 : boolean;
  signal type_cast_1106_inst_ack_1 : boolean;
  signal addr_of_1502_final_reg_ack_1 : boolean;
  signal W_ifx_xend80_exec_guard_1167_delayed_1_0_1245_inst_ack_1 : boolean;
  signal W_ifx_xend80_exec_guard_1167_delayed_1_0_1245_inst_req_1 : boolean;
  signal type_cast_1495_inst_req_0 : boolean;
  signal type_cast_1330_inst_ack_1 : boolean;
  signal W_ifx_xthen_ifx_xend80_taken_1062_delayed_3_0_1121_inst_req_0 : boolean;
  signal W_ifx_xthen_ifx_xend80_taken_1062_delayed_3_0_1121_inst_ack_0 : boolean;
  signal W_ifx_xthen_ifx_xend80_taken_1062_delayed_3_0_1121_inst_req_1 : boolean;
  signal W_ifx_xthen_ifx_xend80_taken_1062_delayed_3_0_1121_inst_ack_1 : boolean;
  signal ptr_deref_1512_store_0_ack_1 : boolean;
  signal ptr_deref_1464_load_0_req_1 : boolean;
  signal type_cast_1126_inst_req_0 : boolean;
  signal W_ifx_xelse155_exec_guard_1338_delayed_1_0_1488_inst_req_0 : boolean;
  signal type_cast_1126_inst_ack_0 : boolean;
  signal type_cast_1126_inst_req_1 : boolean;
  signal type_cast_1126_inst_ack_1 : boolean;
  signal ptr_deref_1464_load_0_ack_1 : boolean;
  signal type_cast_1130_inst_req_0 : boolean;
  signal type_cast_1130_inst_ack_0 : boolean;
  signal type_cast_1130_inst_req_1 : boolean;
  signal type_cast_1130_inst_ack_1 : boolean;
  signal type_cast_1134_inst_req_0 : boolean;
  signal type_cast_1134_inst_ack_0 : boolean;
  signal type_cast_1134_inst_req_1 : boolean;
  signal type_cast_1134_inst_ack_1 : boolean;
  signal W_ifx_xthen152_exec_guard_1256_delayed_1_0_1382_inst_req_0 : boolean;
  signal W_ifx_xthen152_exec_guard_1256_delayed_1_0_1382_inst_ack_0 : boolean;
  signal W_ifx_xthen152_exec_guard_1256_delayed_1_0_1382_inst_req_1 : boolean;
  signal W_ifx_xthen152_exec_guard_1256_delayed_1_0_1382_inst_ack_1 : boolean;
  signal if_stmt_1527_branch_req_0 : boolean;
  signal W_ifx_xthen152_exec_guard_1266_delayed_1_0_1395_inst_req_0 : boolean;
  signal W_ifx_xthen152_exec_guard_1266_delayed_1_0_1395_inst_ack_0 : boolean;
  signal W_ifx_xthen152_exec_guard_1266_delayed_1_0_1395_inst_req_1 : boolean;
  signal array_obj_ref_1501_index_offset_ack_1 : boolean;
  signal W_ifx_xthen152_exec_guard_1266_delayed_1_0_1395_inst_ack_1 : boolean;
  signal W_ifx_xelse155_exec_guard_1328_delayed_1_0_1475_inst_ack_0 : boolean;
  signal array_obj_ref_1501_index_offset_req_1 : boolean;
  signal type_cast_1402_inst_req_0 : boolean;
  signal type_cast_1402_inst_ack_0 : boolean;
  signal type_cast_1402_inst_req_1 : boolean;
  signal type_cast_1402_inst_ack_1 : boolean;
  signal W_ifx_xelse155_exec_guard_1328_delayed_1_0_1475_inst_req_0 : boolean;
  signal array_obj_ref_1408_index_offset_req_0 : boolean;
  signal array_obj_ref_1501_index_offset_ack_0 : boolean;
  signal array_obj_ref_1408_index_offset_ack_0 : boolean;
  signal array_obj_ref_1408_index_offset_req_1 : boolean;
  signal array_obj_ref_1408_index_offset_ack_1 : boolean;
  signal array_obj_ref_1501_index_offset_req_0 : boolean;
  signal addr_of_1409_final_reg_req_0 : boolean;
  signal addr_of_1409_final_reg_ack_0 : boolean;
  signal W_ifx_xelse155_exec_guard_1338_delayed_1_0_1488_inst_ack_1 : boolean;
  signal addr_of_1409_final_reg_req_1 : boolean;
  signal addr_of_1409_final_reg_ack_1 : boolean;
  signal W_arrayidx166_1352_delayed_6_0_1507_inst_ack_1 : boolean;
  signal W_arrayidx166_1352_delayed_6_0_1507_inst_req_1 : boolean;
  signal W_arrayidx166_1352_delayed_6_0_1507_inst_ack_0 : boolean;
  signal W_arrayidx166_1352_delayed_6_0_1507_inst_req_0 : boolean;
  signal type_cast_1473_inst_ack_1 : boolean;
  signal type_cast_1473_inst_req_1 : boolean;
  signal W_ifx_xelse155_exec_guard_1338_delayed_1_0_1488_inst_req_1 : boolean;
  signal ptr_deref_1512_store_0_req_0 : boolean;
  signal ptr_deref_1413_store_0_req_0 : boolean;
  signal ptr_deref_1413_store_0_ack_0 : boolean;
  signal ptr_deref_1413_store_0_req_1 : boolean;
  signal ptr_deref_1413_store_0_ack_1 : boolean;
  signal type_cast_1473_inst_ack_0 : boolean;
  signal W_add118_1290_delayed_2_0_1420_inst_req_0 : boolean;
  signal W_add118_1290_delayed_2_0_1420_inst_ack_0 : boolean;
  signal W_add118_1290_delayed_2_0_1420_inst_req_1 : boolean;
  signal W_add118_1290_delayed_2_0_1420_inst_ack_1 : boolean;
  signal do_while_stmt_903_branch_ack_1 : boolean;
  signal type_cast_1427_inst_req_0 : boolean;
  signal type_cast_1427_inst_ack_0 : boolean;
  signal type_cast_1427_inst_req_1 : boolean;
  signal type_cast_1427_inst_ack_1 : boolean;
  signal type_cast_1473_inst_req_0 : boolean;
  signal W_ifx_xelse155_exec_guard_1351_delayed_15_0_1504_inst_ack_1 : boolean;
  signal W_ifx_xelse155_exec_guard_1294_delayed_1_0_1429_inst_req_0 : boolean;
  signal W_ifx_xelse155_exec_guard_1294_delayed_1_0_1429_inst_ack_0 : boolean;
  signal W_ifx_xelse155_exec_guard_1294_delayed_1_0_1429_inst_req_1 : boolean;
  signal W_ifx_xelse155_exec_guard_1294_delayed_1_0_1429_inst_ack_1 : boolean;
  signal do_while_stmt_903_branch_ack_0 : boolean;
  signal W_ifx_xelse155_exec_guard_1351_delayed_15_0_1504_inst_req_1 : boolean;
  signal WPIPE_Block0_complete_1533_inst_ack_1 : boolean;
  signal W_ifx_xelse155_exec_guard_1304_delayed_1_0_1442_inst_req_0 : boolean;
  signal W_ifx_xelse155_exec_guard_1304_delayed_1_0_1442_inst_ack_0 : boolean;
  signal WPIPE_Block0_complete_1533_inst_req_1 : boolean;
  signal W_ifx_xelse155_exec_guard_1304_delayed_1_0_1442_inst_req_1 : boolean;
  signal W_ifx_xelse155_exec_guard_1304_delayed_1_0_1442_inst_ack_1 : boolean;
  signal W_ifx_xelse155_exec_guard_1351_delayed_15_0_1504_inst_ack_0 : boolean;
  signal WPIPE_Block0_complete_1533_inst_ack_0 : boolean;
  signal type_cast_1449_inst_req_0 : boolean;
  signal type_cast_1449_inst_ack_0 : boolean;
  signal WPIPE_Block0_complete_1533_inst_req_0 : boolean;
  signal type_cast_1449_inst_req_1 : boolean;
  signal type_cast_1449_inst_ack_1 : boolean;
  signal W_ifx_xelse155_exec_guard_1351_delayed_15_0_1504_inst_req_0 : boolean;
  signal W_add96_1324_delayed_2_0_1466_inst_ack_1 : boolean;
  signal W_add96_1324_delayed_2_0_1466_inst_req_1 : boolean;
  signal W_add96_1324_delayed_2_0_1466_inst_ack_0 : boolean;
  signal array_obj_ref_1455_index_offset_req_0 : boolean;
  signal array_obj_ref_1455_index_offset_ack_0 : boolean;
  signal array_obj_ref_1455_index_offset_req_1 : boolean;
  signal array_obj_ref_1455_index_offset_ack_1 : boolean;
  signal ptr_deref_1464_load_0_ack_0 : boolean;
  signal W_ifx_xelse155_exec_guard_1338_delayed_1_0_1488_inst_ack_0 : boolean;
  signal ptr_deref_1464_load_0_req_0 : boolean;
  signal type_cast_1495_inst_ack_1 : boolean;
  signal addr_of_1456_final_reg_req_0 : boolean;
  signal type_cast_1495_inst_req_1 : boolean;
  signal addr_of_1456_final_reg_ack_0 : boolean;
  signal addr_of_1456_final_reg_req_1 : boolean;
  signal addr_of_1456_final_reg_ack_1 : boolean;
  signal W_ifx_xelse155_exec_guard_1317_delayed_9_0_1458_inst_req_0 : boolean;
  signal W_ifx_xelse155_exec_guard_1317_delayed_9_0_1458_inst_ack_0 : boolean;
  signal W_ifx_xelse155_exec_guard_1317_delayed_9_0_1458_inst_req_1 : boolean;
  signal W_ifx_xelse155_exec_guard_1317_delayed_9_0_1458_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "zeropad3D_A_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  zeropad3D_A_CP_1983_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "zeropad3D_A_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= zeropad3D_A_CP_1983_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= zeropad3D_A_CP_1983_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= zeropad3D_A_CP_1983_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  zeropad3D_A_CP_1983: Block -- control-path 
    signal zeropad3D_A_CP_1983_elements: BooleanArray(411 downto 0);
    -- 
  begin -- 
    zeropad3D_A_CP_1983_elements(0) <= zeropad3D_A_CP_1983_start;
    zeropad3D_A_CP_1983_symbol <= zeropad3D_A_CP_1983_elements(411);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_783/$entry
      -- CP-element group 0: 	 branch_block_stmt_783/branch_block_stmt_783__entry__
      -- CP-element group 0: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804__entry__
      -- CP-element group 0: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/$entry
      -- CP-element group 0: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_785_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_785_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_785_Sample/rr
      -- 
    rr_2017_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2017_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(0), ack => RPIPE_Block0_starting_785_inst_req_0); -- 
    -- CP-element group 1:  branch  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	407 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	408 
    -- CP-element group 1: 	409 
    -- CP-element group 1:  members (9) 
      -- CP-element group 1: 	 branch_block_stmt_783/do_while_stmt_903__exit__
      -- CP-element group 1: 	 branch_block_stmt_783/if_stmt_1527__entry__
      -- CP-element group 1: 	 branch_block_stmt_783/if_stmt_1527_else_link/$entry
      -- CP-element group 1: 	 branch_block_stmt_783/if_stmt_1527_if_link/$entry
      -- CP-element group 1: 	 branch_block_stmt_783/if_stmt_1527_eval_test/branch_req
      -- CP-element group 1: 	 branch_block_stmt_783/if_stmt_1527_eval_test/$exit
      -- CP-element group 1: 	 branch_block_stmt_783/if_stmt_1527_eval_test/$entry
      -- CP-element group 1: 	 branch_block_stmt_783/if_stmt_1527_dead_link/$entry
      -- CP-element group 1: 	 branch_block_stmt_783/R_ifx_xend167_whilex_xend_taken_1528_place
      -- 
    branch_req_3606_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3606_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(1), ack => if_stmt_1527_branch_req_0); -- 
    zeropad3D_A_CP_1983_elements(1) <= zeropad3D_A_CP_1983_elements(407);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_785_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_785_update_start_
      -- CP-element group 2: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_785_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_785_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_785_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_785_Update/cr
      -- 
    ra_2018_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_starting_785_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(2)); -- 
    cr_2022_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2022_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(2), ack => RPIPE_Block0_starting_785_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_785_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_785_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_785_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_788_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_788_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_788_Sample/rr
      -- 
    ca_2023_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_starting_785_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(3)); -- 
    rr_2031_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2031_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(3), ack => RPIPE_Block0_starting_788_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_788_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_788_update_start_
      -- CP-element group 4: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_788_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_788_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_788_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_788_Update/cr
      -- 
    ra_2032_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_starting_788_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(4)); -- 
    cr_2036_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2036_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(4), ack => RPIPE_Block0_starting_788_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_788_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_788_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_788_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_791_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_791_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_791_Sample/rr
      -- 
    ca_2037_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_starting_788_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(5)); -- 
    rr_2045_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2045_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(5), ack => RPIPE_Block0_starting_791_inst_req_0); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_791_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_791_update_start_
      -- CP-element group 6: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_791_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_791_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_791_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_791_Update/cr
      -- 
    ra_2046_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_starting_791_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(6)); -- 
    cr_2050_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2050_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(6), ack => RPIPE_Block0_starting_791_inst_req_1); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_791_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_791_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_791_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_794_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_794_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_794_Sample/rr
      -- 
    ca_2051_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_starting_791_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(7)); -- 
    rr_2059_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2059_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(7), ack => RPIPE_Block0_starting_794_inst_req_0); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_794_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_794_update_start_
      -- CP-element group 8: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_794_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_794_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_794_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_794_Update/cr
      -- 
    ra_2060_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_starting_794_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(8)); -- 
    cr_2064_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2064_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(8), ack => RPIPE_Block0_starting_794_inst_req_1); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_794_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_794_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_794_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_797_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_797_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_797_Sample/rr
      -- 
    ca_2065_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_starting_794_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(9)); -- 
    rr_2073_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2073_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(9), ack => RPIPE_Block0_starting_797_inst_req_0); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_797_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_797_update_start_
      -- CP-element group 10: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_797_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_797_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_797_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_797_Update/cr
      -- 
    ra_2074_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_starting_797_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(10)); -- 
    cr_2078_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2078_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(10), ack => RPIPE_Block0_starting_797_inst_req_1); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_797_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_797_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_797_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_800_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_800_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_800_Sample/rr
      -- 
    ca_2079_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_starting_797_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(11)); -- 
    rr_2087_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2087_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(11), ack => RPIPE_Block0_starting_800_inst_req_0); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_800_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_800_update_start_
      -- CP-element group 12: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_800_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_800_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_800_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_800_Update/cr
      -- 
    ra_2088_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_starting_800_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(12)); -- 
    cr_2092_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2092_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(12), ack => RPIPE_Block0_starting_800_inst_req_1); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_800_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_800_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_800_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_803_sample_start_
      -- CP-element group 13: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_803_Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_803_Sample/rr
      -- 
    ca_2093_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_starting_800_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(13)); -- 
    rr_2101_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2101_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(13), ack => RPIPE_Block0_starting_803_inst_req_0); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_803_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_803_update_start_
      -- CP-element group 14: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_803_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_803_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_803_Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_803_Update/cr
      -- 
    ra_2102_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_starting_803_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(14)); -- 
    cr_2106_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2106_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(14), ack => RPIPE_Block0_starting_803_inst_req_1); -- 
    -- CP-element group 15:  fork  transition  place  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15: 	17 
    -- CP-element group 15: 	18 
    -- CP-element group 15: 	19 
    -- CP-element group 15: 	20 
    -- CP-element group 15: 	21 
    -- CP-element group 15: 	22 
    -- CP-element group 15: 	23 
    -- CP-element group 15: 	24 
    -- CP-element group 15: 	25 
    -- CP-element group 15: 	26 
    -- CP-element group 15: 	27 
    -- CP-element group 15: 	28 
    -- CP-element group 15: 	29 
    -- CP-element group 15: 	30 
    -- CP-element group 15: 	31 
    -- CP-element group 15: 	32 
    -- CP-element group 15: 	33 
    -- CP-element group 15:  members (61) 
      -- CP-element group 15: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_854_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_854_update_start_
      -- CP-element group 15: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_868_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_854_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_854_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_854_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_868_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_868_update_start_
      -- CP-element group 15: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_854_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_868_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_839_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_868_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_839_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_868_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804__exit__
      -- CP-element group 15: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884__entry__
      -- CP-element group 15: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/$exit
      -- CP-element group 15: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_803_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_803_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_783/assign_stmt_786_to_assign_stmt_804/RPIPE_Block0_starting_803_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/$entry
      -- CP-element group 15: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_809_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_809_update_start_
      -- CP-element group 15: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_809_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_809_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_809_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_809_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_813_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_813_update_start_
      -- CP-element group 15: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_813_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_813_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_813_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_813_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_817_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_817_update_start_
      -- CP-element group 15: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_817_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_817_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_817_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_817_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_821_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_821_update_start_
      -- CP-element group 15: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_821_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_821_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_821_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_821_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_825_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_825_update_start_
      -- CP-element group 15: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_825_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_825_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_825_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_825_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_835_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_835_update_start_
      -- CP-element group 15: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_835_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_835_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_835_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_835_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_839_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_839_update_start_
      -- CP-element group 15: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_839_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_839_Sample/rr
      -- 
    ca_2107_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_starting_803_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(15)); -- 
    cr_2221_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2221_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(15), ack => type_cast_854_inst_req_1); -- 
    rr_2216_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2216_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(15), ack => type_cast_854_inst_req_0); -- 
    rr_2230_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2230_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(15), ack => type_cast_868_inst_req_0); -- 
    cr_2207_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2207_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(15), ack => type_cast_839_inst_req_1); -- 
    cr_2235_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2235_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(15), ack => type_cast_868_inst_req_1); -- 
    rr_2118_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2118_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(15), ack => type_cast_809_inst_req_0); -- 
    cr_2123_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2123_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(15), ack => type_cast_809_inst_req_1); -- 
    rr_2132_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2132_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(15), ack => type_cast_813_inst_req_0); -- 
    cr_2137_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2137_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(15), ack => type_cast_813_inst_req_1); -- 
    rr_2146_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2146_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(15), ack => type_cast_817_inst_req_0); -- 
    cr_2151_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2151_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(15), ack => type_cast_817_inst_req_1); -- 
    rr_2160_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2160_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(15), ack => type_cast_821_inst_req_0); -- 
    cr_2165_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2165_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(15), ack => type_cast_821_inst_req_1); -- 
    rr_2174_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2174_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(15), ack => type_cast_825_inst_req_0); -- 
    cr_2179_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2179_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(15), ack => type_cast_825_inst_req_1); -- 
    rr_2188_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2188_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(15), ack => type_cast_835_inst_req_0); -- 
    cr_2193_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2193_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(15), ack => type_cast_835_inst_req_1); -- 
    rr_2202_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2202_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(15), ack => type_cast_839_inst_req_0); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_809_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_809_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_809_Sample/ra
      -- 
    ra_2119_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_809_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	15 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	34 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_809_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_809_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_809_Update/ca
      -- 
    ca_2124_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_809_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(17)); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	15 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_813_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_813_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_813_Sample/ra
      -- 
    ra_2133_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_813_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	15 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	34 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_813_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_813_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_813_Update/ca
      -- 
    ca_2138_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_813_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	15 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_817_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_817_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_817_Sample/ra
      -- 
    ra_2147_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_817_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	15 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	34 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_817_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_817_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_817_Update/ca
      -- 
    ca_2152_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_817_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	15 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_821_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_821_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_821_Sample/ra
      -- 
    ra_2161_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_821_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	15 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	34 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_821_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_821_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_821_Update/ca
      -- 
    ca_2166_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_821_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	15 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_825_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_825_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_825_Sample/ra
      -- 
    ra_2175_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_825_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	15 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	34 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_825_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_825_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_825_Update/ca
      -- 
    ca_2180_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_825_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	15 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_835_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_835_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_835_Sample/ra
      -- 
    ra_2189_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_835_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	15 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	34 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_835_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_835_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_835_Update/ca
      -- 
    ca_2194_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_835_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	15 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_839_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_839_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_839_Sample/ra
      -- 
    ra_2203_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_839_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	15 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	34 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_839_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_839_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_839_update_completed_
      -- 
    ca_2208_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_839_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	15 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_854_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_854_Sample/ra
      -- CP-element group 30: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_854_sample_completed_
      -- 
    ra_2217_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_854_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	15 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	34 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_854_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_854_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_854_update_completed_
      -- 
    ca_2222_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_854_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	15 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_868_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_868_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_868_Sample/ra
      -- 
    ra_2231_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_868_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	15 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_868_Update/ca
      -- CP-element group 33: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_868_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/type_cast_868_Update/$exit
      -- 
    ca_2236_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_868_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(33)); -- 
    -- CP-element group 34:  join  transition  place  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	17 
    -- CP-element group 34: 	19 
    -- CP-element group 34: 	21 
    -- CP-element group 34: 	23 
    -- CP-element group 34: 	25 
    -- CP-element group 34: 	27 
    -- CP-element group 34: 	29 
    -- CP-element group 34: 	31 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34:  members (10) 
      -- CP-element group 34: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884__exit__
      -- CP-element group 34: 	 branch_block_stmt_783/entry_whilex_xbody
      -- CP-element group 34: 	 branch_block_stmt_783/merge_stmt_886__exit__
      -- CP-element group 34: 	 branch_block_stmt_783/do_while_stmt_903__entry__
      -- CP-element group 34: 	 branch_block_stmt_783/assign_stmt_810_to_assign_stmt_884/$exit
      -- CP-element group 34: 	 branch_block_stmt_783/merge_stmt_886_PhiReqMerge
      -- CP-element group 34: 	 branch_block_stmt_783/merge_stmt_886_PhiAck/$exit
      -- CP-element group 34: 	 branch_block_stmt_783/merge_stmt_886_PhiAck/$entry
      -- CP-element group 34: 	 branch_block_stmt_783/entry_whilex_xbody_PhiReq/$exit
      -- CP-element group 34: 	 branch_block_stmt_783/entry_whilex_xbody_PhiReq/$entry
      -- 
    zeropad3D_A_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_A_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(17) & zeropad3D_A_CP_1983_elements(19) & zeropad3D_A_CP_1983_elements(21) & zeropad3D_A_CP_1983_elements(23) & zeropad3D_A_CP_1983_elements(25) & zeropad3D_A_CP_1983_elements(27) & zeropad3D_A_CP_1983_elements(29) & zeropad3D_A_CP_1983_elements(31) & zeropad3D_A_CP_1983_elements(33);
      gj_zeropad3D_A_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  transition  place  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	41 
    -- CP-element group 35:  members (2) 
      -- CP-element group 35: 	 branch_block_stmt_783/do_while_stmt_903/$entry
      -- CP-element group 35: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903__entry__
      -- 
    zeropad3D_A_CP_1983_elements(35) <= zeropad3D_A_CP_1983_elements(34);
    -- CP-element group 36:  merge  place  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	407 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903__exit__
      -- 
    -- Element group zeropad3D_A_CP_1983_elements(36) is bound as output of CP function.
    -- CP-element group 37:  merge  place  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	40 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_783/do_while_stmt_903/loop_back
      -- 
    -- Element group zeropad3D_A_CP_1983_elements(37) is bound as output of CP function.
    -- CP-element group 38:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	43 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	405 
    -- CP-element group 38: 	406 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_783/do_while_stmt_903/condition_done
      -- CP-element group 38: 	 branch_block_stmt_783/do_while_stmt_903/loop_taken/$entry
      -- CP-element group 38: 	 branch_block_stmt_783/do_while_stmt_903/loop_exit/$entry
      -- 
    zeropad3D_A_CP_1983_elements(38) <= zeropad3D_A_CP_1983_elements(43);
    -- CP-element group 39:  branch  place  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	404 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_783/do_while_stmt_903/loop_body_done
      -- 
    zeropad3D_A_CP_1983_elements(39) <= zeropad3D_A_CP_1983_elements(404);
    -- CP-element group 40:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	37 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	52 
    -- CP-element group 40: 	73 
    -- CP-element group 40: 	94 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/back_edge_to_loop_body
      -- 
    zeropad3D_A_CP_1983_elements(40) <= zeropad3D_A_CP_1983_elements(37);
    -- CP-element group 41:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	35 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	54 
    -- CP-element group 41: 	75 
    -- CP-element group 41: 	96 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/first_time_through_loop_body
      -- 
    zeropad3D_A_CP_1983_elements(41) <= zeropad3D_A_CP_1983_elements(35);
    -- CP-element group 42:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	402 
    -- CP-element group 42: 	384 
    -- CP-element group 42: 	385 
    -- CP-element group 42: 	48 
    -- CP-element group 42: 	49 
    -- CP-element group 42: 	67 
    -- CP-element group 42: 	68 
    -- CP-element group 42: 	88 
    -- CP-element group 42: 	89 
    -- CP-element group 42: 	113 
    -- CP-element group 42: 	241 
    -- CP-element group 42: 	277 
    -- CP-element group 42: 	318 
    -- CP-element group 42: 	319 
    -- CP-element group 42: 	349 
    -- CP-element group 42: 	350 
    -- CP-element group 42:  members (2) 
      -- CP-element group 42: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/$entry
      -- CP-element group 42: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/loop_body_start
      -- 
    -- Element group zeropad3D_A_CP_1983_elements(42) is bound as output of CP function.
    -- CP-element group 43:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	402 
    -- CP-element group 43: 	47 
    -- CP-element group 43: 	164 
    -- CP-element group 43: 	172 
    -- CP-element group 43: 	176 
    -- CP-element group 43: 	224 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	38 
    -- CP-element group 43:  members (1) 
      -- CP-element group 43: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/condition_evaluated
      -- 
    condition_evaluated_2251_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_2251_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(43), ack => do_while_stmt_903_branch_req_0); -- 
    zeropad3D_A_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_A_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(402) & zeropad3D_A_CP_1983_elements(47) & zeropad3D_A_CP_1983_elements(164) & zeropad3D_A_CP_1983_elements(172) & zeropad3D_A_CP_1983_elements(176) & zeropad3D_A_CP_1983_elements(224);
      gj_zeropad3D_A_cp_element_group_43 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	48 
    -- CP-element group 44: 	67 
    -- CP-element group 44: 	88 
    -- CP-element group 44: marked-predecessors 
    -- CP-element group 44: 	47 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	69 
    -- CP-element group 44: 	90 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/phi_stmt_905_sample_start__ps
      -- CP-element group 44: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/aggregated_phi_sample_req
      -- 
    zeropad3D_A_cp_element_group_44: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_A_cp_element_group_44"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(48) & zeropad3D_A_CP_1983_elements(67) & zeropad3D_A_CP_1983_elements(88) & zeropad3D_A_CP_1983_elements(47);
      gj_zeropad3D_A_cp_element_group_44 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(44), clk => clk, reset => reset); --
    end block;
    -- CP-element group 45:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	50 
    -- CP-element group 45: 	70 
    -- CP-element group 45: 	91 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	162 
    -- CP-element group 45: 	170 
    -- CP-element group 45: 	174 
    -- CP-element group 45: 	182 
    -- CP-element group 45: 	186 
    -- CP-element group 45: 	190 
    -- CP-element group 45: 	194 
    -- CP-element group 45: 	198 
    -- CP-element group 45: 	202 
    -- CP-element group 45: 	206 
    -- CP-element group 45: 	210 
    -- CP-element group 45: 	214 
    -- CP-element group 45: 	218 
    -- CP-element group 45: marked-successors 
    -- CP-element group 45: 	48 
    -- CP-element group 45: 	67 
    -- CP-element group 45: 	88 
    -- CP-element group 45:  members (4) 
      -- CP-element group 45: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/phi_stmt_915_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/phi_stmt_905_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/phi_stmt_910_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/aggregated_phi_sample_ack
      -- 
    zeropad3D_A_cp_element_group_45: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_A_cp_element_group_45"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(50) & zeropad3D_A_CP_1983_elements(70) & zeropad3D_A_CP_1983_elements(91);
      gj_zeropad3D_A_cp_element_group_45 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(45), clk => clk, reset => reset); --
    end block;
    -- CP-element group 46:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	49 
    -- CP-element group 46: 	68 
    -- CP-element group 46: 	89 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	71 
    -- CP-element group 46: 	92 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/phi_stmt_905_update_start__ps
      -- CP-element group 46: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/aggregated_phi_update_req
      -- 
    zeropad3D_A_cp_element_group_46: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_A_cp_element_group_46"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(49) & zeropad3D_A_CP_1983_elements(68) & zeropad3D_A_CP_1983_elements(89);
      gj_zeropad3D_A_cp_element_group_46 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(46), clk => clk, reset => reset); --
    end block;
    -- CP-element group 47:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	51 
    -- CP-element group 47: 	72 
    -- CP-element group 47: 	93 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	43 
    -- CP-element group 47: marked-successors 
    -- CP-element group 47: 	44 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/aggregated_phi_update_ack
      -- 
    zeropad3D_A_cp_element_group_47: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_A_cp_element_group_47"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(51) & zeropad3D_A_CP_1983_elements(72) & zeropad3D_A_CP_1983_elements(93);
      gj_zeropad3D_A_cp_element_group_47 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(47), clk => clk, reset => reset); --
    end block;
    -- CP-element group 48:  join  transition  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	42 
    -- CP-element group 48: marked-predecessors 
    -- CP-element group 48: 	45 
    -- CP-element group 48: 	164 
    -- CP-element group 48: 	172 
    -- CP-element group 48: 	176 
    -- CP-element group 48: 	184 
    -- CP-element group 48: 	188 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	44 
    -- CP-element group 48:  members (1) 
      -- CP-element group 48: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/phi_stmt_905_sample_start_
      -- 
    zeropad3D_A_cp_element_group_48: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_A_cp_element_group_48"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(42) & zeropad3D_A_CP_1983_elements(45) & zeropad3D_A_CP_1983_elements(164) & zeropad3D_A_CP_1983_elements(172) & zeropad3D_A_CP_1983_elements(176) & zeropad3D_A_CP_1983_elements(184) & zeropad3D_A_CP_1983_elements(188);
      gj_zeropad3D_A_cp_element_group_48 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(48), clk => clk, reset => reset); --
    end block;
    -- CP-element group 49:  join  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	42 
    -- CP-element group 49: marked-predecessors 
    -- CP-element group 49: 	51 
    -- CP-element group 49: 	111 
    -- CP-element group 49: 	119 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	46 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/phi_stmt_905_update_start_
      -- 
    zeropad3D_A_cp_element_group_49: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_A_cp_element_group_49"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(42) & zeropad3D_A_CP_1983_elements(51) & zeropad3D_A_CP_1983_elements(111) & zeropad3D_A_CP_1983_elements(119);
      gj_zeropad3D_A_cp_element_group_49 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(49), clk => clk, reset => reset); --
    end block;
    -- CP-element group 50:  join  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	45 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/phi_stmt_905_sample_completed__ps
      -- 
    -- Element group zeropad3D_A_CP_1983_elements(50) is bound as output of CP function.
    -- CP-element group 51:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	47 
    -- CP-element group 51: 	109 
    -- CP-element group 51: 	117 
    -- CP-element group 51: marked-successors 
    -- CP-element group 51: 	49 
    -- CP-element group 51:  members (2) 
      -- CP-element group 51: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/phi_stmt_905_update_completed__ps
      -- CP-element group 51: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/phi_stmt_905_update_completed_
      -- 
    -- Element group zeropad3D_A_CP_1983_elements(51) is bound as output of CP function.
    -- CP-element group 52:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	40 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (1) 
      -- CP-element group 52: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/phi_stmt_905_loopback_trigger
      -- 
    zeropad3D_A_CP_1983_elements(52) <= zeropad3D_A_CP_1983_elements(40);
    -- CP-element group 53:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (2) 
      -- CP-element group 53: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/phi_stmt_905_loopback_sample_req
      -- CP-element group 53: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/phi_stmt_905_loopback_sample_req_ps
      -- 
    phi_stmt_905_loopback_sample_req_2266_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_905_loopback_sample_req_2266_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(53), ack => phi_stmt_905_req_0); -- 
    -- Element group zeropad3D_A_CP_1983_elements(53) is bound as output of CP function.
    -- CP-element group 54:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	41 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (1) 
      -- CP-element group 54: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/phi_stmt_905_entry_trigger
      -- 
    zeropad3D_A_CP_1983_elements(54) <= zeropad3D_A_CP_1983_elements(41);
    -- CP-element group 55:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (2) 
      -- CP-element group 55: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/phi_stmt_905_entry_sample_req_ps
      -- CP-element group 55: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/phi_stmt_905_entry_sample_req
      -- 
    phi_stmt_905_entry_sample_req_2269_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_905_entry_sample_req_2269_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(55), ack => phi_stmt_905_req_1); -- 
    -- Element group zeropad3D_A_CP_1983_elements(55) is bound as output of CP function.
    -- CP-element group 56:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (2) 
      -- CP-element group 56: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/phi_stmt_905_phi_mux_ack
      -- CP-element group 56: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/phi_stmt_905_phi_mux_ack_ps
      -- 
    phi_stmt_905_phi_mux_ack_2272_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_905_ack_0, ack => zeropad3D_A_CP_1983_elements(56)); -- 
    -- CP-element group 57:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	59 
    -- CP-element group 57:  members (1) 
      -- CP-element group 57: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_908_sample_start__ps
      -- 
    -- Element group zeropad3D_A_CP_1983_elements(57) is bound as output of CP function.
    -- CP-element group 58:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	60 
    -- CP-element group 58:  members (1) 
      -- CP-element group 58: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_908_update_start__ps
      -- 
    -- Element group zeropad3D_A_CP_1983_elements(58) is bound as output of CP function.
    -- CP-element group 59:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	57 
    -- CP-element group 59: marked-predecessors 
    -- CP-element group 59: 	61 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	61 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_908_sample_start_
      -- CP-element group 59: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_908_Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_908_Sample/rr
      -- 
    rr_2285_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2285_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(59), ack => type_cast_908_inst_req_0); -- 
    zeropad3D_A_cp_element_group_59: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "zeropad3D_A_cp_element_group_59"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(57) & zeropad3D_A_CP_1983_elements(61);
      gj_zeropad3D_A_cp_element_group_59 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(59), clk => clk, reset => reset); --
    end block;
    -- CP-element group 60:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	58 
    -- CP-element group 60: marked-predecessors 
    -- CP-element group 60: 	62 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	62 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_908_update_start_
      -- CP-element group 60: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_908_Update/cr
      -- CP-element group 60: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_908_Update/$entry
      -- 
    cr_2290_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2290_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(60), ack => type_cast_908_inst_req_1); -- 
    zeropad3D_A_cp_element_group_60: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_A_cp_element_group_60"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(58) & zeropad3D_A_CP_1983_elements(62);
      gj_zeropad3D_A_cp_element_group_60 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(60), clk => clk, reset => reset); --
    end block;
    -- CP-element group 61:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	59 
    -- CP-element group 61: successors 
    -- CP-element group 61: marked-successors 
    -- CP-element group 61: 	59 
    -- CP-element group 61:  members (4) 
      -- CP-element group 61: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_908_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_908_sample_completed__ps
      -- CP-element group 61: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_908_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_908_Sample/ra
      -- 
    ra_2286_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_908_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(61)); -- 
    -- CP-element group 62:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	60 
    -- CP-element group 62: successors 
    -- CP-element group 62: marked-successors 
    -- CP-element group 62: 	60 
    -- CP-element group 62:  members (4) 
      -- CP-element group 62: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_908_update_completed__ps
      -- CP-element group 62: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_908_Update/ca
      -- CP-element group 62: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_908_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_908_Update/$exit
      -- 
    ca_2291_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_908_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(62)); -- 
    -- CP-element group 63:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (4) 
      -- CP-element group 63: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/R_kx_x1_at_entry_909_sample_completed__ps
      -- CP-element group 63: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/R_kx_x1_at_entry_909_sample_start__ps
      -- CP-element group 63: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/R_kx_x1_at_entry_909_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/R_kx_x1_at_entry_909_sample_start_
      -- 
    -- Element group zeropad3D_A_CP_1983_elements(63) is bound as output of CP function.
    -- CP-element group 64:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	66 
    -- CP-element group 64:  members (2) 
      -- CP-element group 64: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/R_kx_x1_at_entry_909_update_start__ps
      -- CP-element group 64: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/R_kx_x1_at_entry_909_update_start_
      -- 
    -- Element group zeropad3D_A_CP_1983_elements(64) is bound as output of CP function.
    -- CP-element group 65:  join  transition  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	66 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (1) 
      -- CP-element group 65: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/R_kx_x1_at_entry_909_update_completed__ps
      -- 
    zeropad3D_A_CP_1983_elements(65) <= zeropad3D_A_CP_1983_elements(66);
    -- CP-element group 66:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	64 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	65 
    -- CP-element group 66:  members (1) 
      -- CP-element group 66: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/R_kx_x1_at_entry_909_update_completed_
      -- 
    -- Element group zeropad3D_A_CP_1983_elements(66) is a control-delay.
    cp_element_66_delay: control_delay_element  generic map(name => " 66_delay", delay_value => 1)  port map(req => zeropad3D_A_CP_1983_elements(64), ack => zeropad3D_A_CP_1983_elements(66), clk => clk, reset =>reset);
    -- CP-element group 67:  join  transition  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	42 
    -- CP-element group 67: marked-predecessors 
    -- CP-element group 67: 	45 
    -- CP-element group 67: 	164 
    -- CP-element group 67: 	172 
    -- CP-element group 67: 	176 
    -- CP-element group 67: 	192 
    -- CP-element group 67: 	196 
    -- CP-element group 67: 	200 
    -- CP-element group 67: 	204 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	44 
    -- CP-element group 67:  members (1) 
      -- CP-element group 67: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/phi_stmt_910_sample_start_
      -- 
    zeropad3D_A_cp_element_group_67: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_A_cp_element_group_67"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(42) & zeropad3D_A_CP_1983_elements(45) & zeropad3D_A_CP_1983_elements(164) & zeropad3D_A_CP_1983_elements(172) & zeropad3D_A_CP_1983_elements(176) & zeropad3D_A_CP_1983_elements(192) & zeropad3D_A_CP_1983_elements(196) & zeropad3D_A_CP_1983_elements(200) & zeropad3D_A_CP_1983_elements(204);
      gj_zeropad3D_A_cp_element_group_67 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(67), clk => clk, reset => reset); --
    end block;
    -- CP-element group 68:  join  transition  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	42 
    -- CP-element group 68: marked-predecessors 
    -- CP-element group 68: 	72 
    -- CP-element group 68: 	147 
    -- CP-element group 68: 	195 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	46 
    -- CP-element group 68:  members (1) 
      -- CP-element group 68: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/phi_stmt_910_update_start_
      -- 
    zeropad3D_A_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_A_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(42) & zeropad3D_A_CP_1983_elements(72) & zeropad3D_A_CP_1983_elements(147) & zeropad3D_A_CP_1983_elements(195);
      gj_zeropad3D_A_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	44 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (1) 
      -- CP-element group 69: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/phi_stmt_910_sample_start__ps
      -- 
    zeropad3D_A_CP_1983_elements(69) <= zeropad3D_A_CP_1983_elements(44);
    -- CP-element group 70:  join  transition  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	45 
    -- CP-element group 70:  members (1) 
      -- CP-element group 70: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/phi_stmt_910_sample_completed__ps
      -- 
    -- Element group zeropad3D_A_CP_1983_elements(70) is bound as output of CP function.
    -- CP-element group 71:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	46 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (1) 
      -- CP-element group 71: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/phi_stmt_910_update_start__ps
      -- 
    zeropad3D_A_CP_1983_elements(71) <= zeropad3D_A_CP_1983_elements(46);
    -- CP-element group 72:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	47 
    -- CP-element group 72: 	145 
    -- CP-element group 72: 	193 
    -- CP-element group 72: marked-successors 
    -- CP-element group 72: 	68 
    -- CP-element group 72:  members (2) 
      -- CP-element group 72: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/phi_stmt_910_update_completed__ps
      -- CP-element group 72: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/phi_stmt_910_update_completed_
      -- 
    -- Element group zeropad3D_A_CP_1983_elements(72) is bound as output of CP function.
    -- CP-element group 73:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	40 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (1) 
      -- CP-element group 73: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/phi_stmt_910_loopback_trigger
      -- 
    zeropad3D_A_CP_1983_elements(73) <= zeropad3D_A_CP_1983_elements(40);
    -- CP-element group 74:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (2) 
      -- CP-element group 74: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/phi_stmt_910_loopback_sample_req_ps
      -- CP-element group 74: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/phi_stmt_910_loopback_sample_req
      -- 
    phi_stmt_910_loopback_sample_req_2310_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_910_loopback_sample_req_2310_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(74), ack => phi_stmt_910_req_0); -- 
    -- Element group zeropad3D_A_CP_1983_elements(74) is bound as output of CP function.
    -- CP-element group 75:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	41 
    -- CP-element group 75: successors 
    -- CP-element group 75:  members (1) 
      -- CP-element group 75: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/phi_stmt_910_entry_trigger
      -- 
    zeropad3D_A_CP_1983_elements(75) <= zeropad3D_A_CP_1983_elements(41);
    -- CP-element group 76:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (2) 
      -- CP-element group 76: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/phi_stmt_910_entry_sample_req
      -- CP-element group 76: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/phi_stmt_910_entry_sample_req_ps
      -- 
    phi_stmt_910_entry_sample_req_2313_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_910_entry_sample_req_2313_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(76), ack => phi_stmt_910_req_1); -- 
    -- Element group zeropad3D_A_CP_1983_elements(76) is bound as output of CP function.
    -- CP-element group 77:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: successors 
    -- CP-element group 77:  members (2) 
      -- CP-element group 77: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/phi_stmt_910_phi_mux_ack
      -- CP-element group 77: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/phi_stmt_910_phi_mux_ack_ps
      -- 
    phi_stmt_910_phi_mux_ack_2316_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_910_ack_0, ack => zeropad3D_A_CP_1983_elements(77)); -- 
    -- CP-element group 78:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	80 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_913_sample_start__ps
      -- 
    -- Element group zeropad3D_A_CP_1983_elements(78) is bound as output of CP function.
    -- CP-element group 79:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	81 
    -- CP-element group 79:  members (1) 
      -- CP-element group 79: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_913_update_start__ps
      -- 
    -- Element group zeropad3D_A_CP_1983_elements(79) is bound as output of CP function.
    -- CP-element group 80:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: marked-predecessors 
    -- CP-element group 80: 	82 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	82 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_913_sample_start_
      -- CP-element group 80: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_913_Sample/$entry
      -- CP-element group 80: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_913_Sample/rr
      -- 
    rr_2329_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2329_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(80), ack => type_cast_913_inst_req_0); -- 
    zeropad3D_A_cp_element_group_80: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "zeropad3D_A_cp_element_group_80"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(78) & zeropad3D_A_CP_1983_elements(82);
      gj_zeropad3D_A_cp_element_group_80 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(80), clk => clk, reset => reset); --
    end block;
    -- CP-element group 81:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	79 
    -- CP-element group 81: marked-predecessors 
    -- CP-element group 81: 	83 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	83 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_913_Update/cr
      -- CP-element group 81: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_913_Update/$entry
      -- CP-element group 81: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_913_update_start_
      -- 
    cr_2334_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2334_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(81), ack => type_cast_913_inst_req_1); -- 
    zeropad3D_A_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_A_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(79) & zeropad3D_A_CP_1983_elements(83);
      gj_zeropad3D_A_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	80 
    -- CP-element group 82: successors 
    -- CP-element group 82: marked-successors 
    -- CP-element group 82: 	80 
    -- CP-element group 82:  members (4) 
      -- CP-element group 82: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_913_sample_completed_
      -- CP-element group 82: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_913_Sample/ra
      -- CP-element group 82: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_913_sample_completed__ps
      -- CP-element group 82: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_913_Sample/$exit
      -- 
    ra_2330_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_913_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(82)); -- 
    -- CP-element group 83:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	81 
    -- CP-element group 83: successors 
    -- CP-element group 83: marked-successors 
    -- CP-element group 83: 	81 
    -- CP-element group 83:  members (4) 
      -- CP-element group 83: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_913_Update/ca
      -- CP-element group 83: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_913_Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_913_update_completed_
      -- CP-element group 83: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_913_update_completed__ps
      -- 
    ca_2335_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_913_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(83)); -- 
    -- CP-element group 84:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (4) 
      -- CP-element group 84: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/R_ix_x2_at_entry_914_sample_start__ps
      -- CP-element group 84: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/R_ix_x2_at_entry_914_sample_completed_
      -- CP-element group 84: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/R_ix_x2_at_entry_914_sample_start_
      -- CP-element group 84: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/R_ix_x2_at_entry_914_sample_completed__ps
      -- 
    -- Element group zeropad3D_A_CP_1983_elements(84) is bound as output of CP function.
    -- CP-element group 85:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (2) 
      -- CP-element group 85: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/R_ix_x2_at_entry_914_update_start_
      -- CP-element group 85: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/R_ix_x2_at_entry_914_update_start__ps
      -- 
    -- Element group zeropad3D_A_CP_1983_elements(85) is bound as output of CP function.
    -- CP-element group 86:  join  transition  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	87 
    -- CP-element group 86: successors 
    -- CP-element group 86:  members (1) 
      -- CP-element group 86: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/R_ix_x2_at_entry_914_update_completed__ps
      -- 
    zeropad3D_A_CP_1983_elements(86) <= zeropad3D_A_CP_1983_elements(87);
    -- CP-element group 87:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	86 
    -- CP-element group 87:  members (1) 
      -- CP-element group 87: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/R_ix_x2_at_entry_914_update_completed_
      -- 
    -- Element group zeropad3D_A_CP_1983_elements(87) is a control-delay.
    cp_element_87_delay: control_delay_element  generic map(name => " 87_delay", delay_value => 1)  port map(req => zeropad3D_A_CP_1983_elements(85), ack => zeropad3D_A_CP_1983_elements(87), clk => clk, reset =>reset);
    -- CP-element group 88:  join  transition  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	42 
    -- CP-element group 88: marked-predecessors 
    -- CP-element group 88: 	45 
    -- CP-element group 88: 	164 
    -- CP-element group 88: 	172 
    -- CP-element group 88: 	176 
    -- CP-element group 88: 	208 
    -- CP-element group 88: 	212 
    -- CP-element group 88: 	216 
    -- CP-element group 88: 	220 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	44 
    -- CP-element group 88:  members (1) 
      -- CP-element group 88: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/phi_stmt_915_sample_start_
      -- 
    zeropad3D_A_cp_element_group_88: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_A_cp_element_group_88"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(42) & zeropad3D_A_CP_1983_elements(45) & zeropad3D_A_CP_1983_elements(164) & zeropad3D_A_CP_1983_elements(172) & zeropad3D_A_CP_1983_elements(176) & zeropad3D_A_CP_1983_elements(208) & zeropad3D_A_CP_1983_elements(212) & zeropad3D_A_CP_1983_elements(216) & zeropad3D_A_CP_1983_elements(220);
      gj_zeropad3D_A_cp_element_group_88 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(88), clk => clk, reset => reset); --
    end block;
    -- CP-element group 89:  join  transition  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	42 
    -- CP-element group 89: marked-predecessors 
    -- CP-element group 89: 	93 
    -- CP-element group 89: 	123 
    -- CP-element group 89: 	211 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	46 
    -- CP-element group 89:  members (1) 
      -- CP-element group 89: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/phi_stmt_915_update_start_
      -- 
    zeropad3D_A_cp_element_group_89: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 31) := "zeropad3D_A_cp_element_group_89"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(42) & zeropad3D_A_CP_1983_elements(93) & zeropad3D_A_CP_1983_elements(123) & zeropad3D_A_CP_1983_elements(211);
      gj_zeropad3D_A_cp_element_group_89 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(89), clk => clk, reset => reset); --
    end block;
    -- CP-element group 90:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	44 
    -- CP-element group 90: successors 
    -- CP-element group 90:  members (1) 
      -- CP-element group 90: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/phi_stmt_915_sample_start__ps
      -- 
    zeropad3D_A_CP_1983_elements(90) <= zeropad3D_A_CP_1983_elements(44);
    -- CP-element group 91:  join  transition  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	45 
    -- CP-element group 91:  members (1) 
      -- CP-element group 91: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/phi_stmt_915_sample_completed__ps
      -- 
    -- Element group zeropad3D_A_CP_1983_elements(91) is bound as output of CP function.
    -- CP-element group 92:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	46 
    -- CP-element group 92: successors 
    -- CP-element group 92:  members (1) 
      -- CP-element group 92: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/phi_stmt_915_update_start__ps
      -- 
    zeropad3D_A_CP_1983_elements(92) <= zeropad3D_A_CP_1983_elements(46);
    -- CP-element group 93:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	47 
    -- CP-element group 93: 	121 
    -- CP-element group 93: 	209 
    -- CP-element group 93: marked-successors 
    -- CP-element group 93: 	89 
    -- CP-element group 93:  members (2) 
      -- CP-element group 93: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/phi_stmt_915_update_completed__ps
      -- CP-element group 93: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/phi_stmt_915_update_completed_
      -- 
    -- Element group zeropad3D_A_CP_1983_elements(93) is bound as output of CP function.
    -- CP-element group 94:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	40 
    -- CP-element group 94: successors 
    -- CP-element group 94:  members (1) 
      -- CP-element group 94: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/phi_stmt_915_loopback_trigger
      -- 
    zeropad3D_A_CP_1983_elements(94) <= zeropad3D_A_CP_1983_elements(40);
    -- CP-element group 95:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: successors 
    -- CP-element group 95:  members (2) 
      -- CP-element group 95: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/phi_stmt_915_loopback_sample_req_ps
      -- CP-element group 95: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/phi_stmt_915_loopback_sample_req
      -- 
    phi_stmt_915_loopback_sample_req_2354_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_915_loopback_sample_req_2354_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(95), ack => phi_stmt_915_req_0); -- 
    -- Element group zeropad3D_A_CP_1983_elements(95) is bound as output of CP function.
    -- CP-element group 96:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	41 
    -- CP-element group 96: successors 
    -- CP-element group 96:  members (1) 
      -- CP-element group 96: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/phi_stmt_915_entry_trigger
      -- 
    zeropad3D_A_CP_1983_elements(96) <= zeropad3D_A_CP_1983_elements(41);
    -- CP-element group 97:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: successors 
    -- CP-element group 97:  members (2) 
      -- CP-element group 97: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/phi_stmt_915_entry_sample_req
      -- CP-element group 97: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/phi_stmt_915_entry_sample_req_ps
      -- 
    phi_stmt_915_entry_sample_req_2357_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_915_entry_sample_req_2357_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(97), ack => phi_stmt_915_req_1); -- 
    -- Element group zeropad3D_A_CP_1983_elements(97) is bound as output of CP function.
    -- CP-element group 98:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: successors 
    -- CP-element group 98:  members (2) 
      -- CP-element group 98: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/phi_stmt_915_phi_mux_ack_ps
      -- CP-element group 98: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/phi_stmt_915_phi_mux_ack
      -- 
    phi_stmt_915_phi_mux_ack_2360_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_915_ack_0, ack => zeropad3D_A_CP_1983_elements(98)); -- 
    -- CP-element group 99:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	101 
    -- CP-element group 99:  members (1) 
      -- CP-element group 99: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_918_sample_start__ps
      -- 
    -- Element group zeropad3D_A_CP_1983_elements(99) is bound as output of CP function.
    -- CP-element group 100:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	102 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_918_update_start__ps
      -- 
    -- Element group zeropad3D_A_CP_1983_elements(100) is bound as output of CP function.
    -- CP-element group 101:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	99 
    -- CP-element group 101: marked-predecessors 
    -- CP-element group 101: 	103 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	103 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_918_sample_start_
      -- CP-element group 101: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_918_Sample/$entry
      -- CP-element group 101: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_918_Sample/rr
      -- 
    rr_2373_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2373_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(101), ack => type_cast_918_inst_req_0); -- 
    zeropad3D_A_cp_element_group_101: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_101"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(99) & zeropad3D_A_CP_1983_elements(103);
      gj_zeropad3D_A_cp_element_group_101 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(101), clk => clk, reset => reset); --
    end block;
    -- CP-element group 102:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	100 
    -- CP-element group 102: marked-predecessors 
    -- CP-element group 102: 	104 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	104 
    -- CP-element group 102:  members (3) 
      -- CP-element group 102: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_918_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_918_Update/cr
      -- CP-element group 102: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_918_update_start_
      -- 
    cr_2378_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2378_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(102), ack => type_cast_918_inst_req_1); -- 
    zeropad3D_A_cp_element_group_102: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_102"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(100) & zeropad3D_A_CP_1983_elements(104);
      gj_zeropad3D_A_cp_element_group_102 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(102), clk => clk, reset => reset); --
    end block;
    -- CP-element group 103:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	101 
    -- CP-element group 103: successors 
    -- CP-element group 103: marked-successors 
    -- CP-element group 103: 	101 
    -- CP-element group 103:  members (4) 
      -- CP-element group 103: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_918_sample_completed__ps
      -- CP-element group 103: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_918_sample_completed_
      -- CP-element group 103: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_918_Sample/$exit
      -- CP-element group 103: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_918_Sample/ra
      -- 
    ra_2374_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_918_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(103)); -- 
    -- CP-element group 104:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	102 
    -- CP-element group 104: successors 
    -- CP-element group 104: marked-successors 
    -- CP-element group 104: 	102 
    -- CP-element group 104:  members (4) 
      -- CP-element group 104: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_918_Update/ca
      -- CP-element group 104: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_918_update_completed__ps
      -- CP-element group 104: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_918_Update/$exit
      -- CP-element group 104: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_918_update_completed_
      -- 
    ca_2379_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_918_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(104)); -- 
    -- CP-element group 105:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: successors 
    -- CP-element group 105:  members (4) 
      -- CP-element group 105: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/R_jx_x1_at_entry_919_sample_start__ps
      -- CP-element group 105: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/R_jx_x1_at_entry_919_sample_start_
      -- CP-element group 105: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/R_jx_x1_at_entry_919_sample_completed_
      -- CP-element group 105: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/R_jx_x1_at_entry_919_sample_completed__ps
      -- 
    -- Element group zeropad3D_A_CP_1983_elements(105) is bound as output of CP function.
    -- CP-element group 106:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	108 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/R_jx_x1_at_entry_919_update_start_
      -- CP-element group 106: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/R_jx_x1_at_entry_919_update_start__ps
      -- 
    -- Element group zeropad3D_A_CP_1983_elements(106) is bound as output of CP function.
    -- CP-element group 107:  join  transition  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	108 
    -- CP-element group 107: successors 
    -- CP-element group 107:  members (1) 
      -- CP-element group 107: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/R_jx_x1_at_entry_919_update_completed__ps
      -- 
    zeropad3D_A_CP_1983_elements(107) <= zeropad3D_A_CP_1983_elements(108);
    -- CP-element group 108:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	106 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	107 
    -- CP-element group 108:  members (1) 
      -- CP-element group 108: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/R_jx_x1_at_entry_919_update_completed_
      -- 
    -- Element group zeropad3D_A_CP_1983_elements(108) is a control-delay.
    cp_element_108_delay: control_delay_element  generic map(name => " 108_delay", delay_value => 1)  port map(req => zeropad3D_A_CP_1983_elements(106), ack => zeropad3D_A_CP_1983_elements(108), clk => clk, reset =>reset);
    -- CP-element group 109:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	51 
    -- CP-element group 109: marked-predecessors 
    -- CP-element group 109: 	111 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_923_Sample/$entry
      -- CP-element group 109: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_923_sample_start_
      -- CP-element group 109: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_923_Sample/rr
      -- 
    rr_2396_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2396_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(109), ack => type_cast_923_inst_req_0); -- 
    zeropad3D_A_cp_element_group_109: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_109"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(51) & zeropad3D_A_CP_1983_elements(111);
      gj_zeropad3D_A_cp_element_group_109 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(109), clk => clk, reset => reset); --
    end block;
    -- CP-element group 110:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: marked-predecessors 
    -- CP-element group 110: 	112 
    -- CP-element group 110: 	127 
    -- CP-element group 110: 	131 
    -- CP-element group 110: 	135 
    -- CP-element group 110: 	143 
    -- CP-element group 110: 	151 
    -- CP-element group 110: 	159 
    -- CP-element group 110: 	167 
    -- CP-element group 110: 	171 
    -- CP-element group 110: 	175 
    -- CP-element group 110: 	179 
    -- CP-element group 110: 	183 
    -- CP-element group 110: 	191 
    -- CP-element group 110: 	207 
    -- CP-element group 110: 	223 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	112 
    -- CP-element group 110:  members (3) 
      -- CP-element group 110: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_923_update_start_
      -- CP-element group 110: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_923_Update/$entry
      -- CP-element group 110: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_923_Update/cr
      -- 
    cr_2401_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2401_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(110), ack => type_cast_923_inst_req_1); -- 
    zeropad3D_A_cp_element_group_110: block -- 
      constant place_capacities: IntegerArray(0 to 14) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1);
      constant place_markings: IntegerArray(0 to 14)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1);
      constant place_delays: IntegerArray(0 to 14) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_110"; 
      signal preds: BooleanArray(1 to 15); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(112) & zeropad3D_A_CP_1983_elements(127) & zeropad3D_A_CP_1983_elements(131) & zeropad3D_A_CP_1983_elements(135) & zeropad3D_A_CP_1983_elements(143) & zeropad3D_A_CP_1983_elements(151) & zeropad3D_A_CP_1983_elements(159) & zeropad3D_A_CP_1983_elements(167) & zeropad3D_A_CP_1983_elements(171) & zeropad3D_A_CP_1983_elements(175) & zeropad3D_A_CP_1983_elements(179) & zeropad3D_A_CP_1983_elements(183) & zeropad3D_A_CP_1983_elements(191) & zeropad3D_A_CP_1983_elements(207) & zeropad3D_A_CP_1983_elements(223);
      gj_zeropad3D_A_cp_element_group_110 : generic_join generic map(name => joinName, number_of_predecessors => 15, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(110), clk => clk, reset => reset); --
    end block;
    -- CP-element group 111:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: successors 
    -- CP-element group 111: marked-successors 
    -- CP-element group 111: 	49 
    -- CP-element group 111: 	109 
    -- CP-element group 111:  members (3) 
      -- CP-element group 111: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_923_Sample/ra
      -- CP-element group 111: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_923_Sample/$exit
      -- CP-element group 111: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_923_sample_completed_
      -- 
    ra_2397_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_923_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(111)); -- 
    -- CP-element group 112:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	110 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	125 
    -- CP-element group 112: 	129 
    -- CP-element group 112: 	133 
    -- CP-element group 112: 	141 
    -- CP-element group 112: 	149 
    -- CP-element group 112: 	157 
    -- CP-element group 112: 	165 
    -- CP-element group 112: 	169 
    -- CP-element group 112: 	173 
    -- CP-element group 112: 	177 
    -- CP-element group 112: 	181 
    -- CP-element group 112: 	189 
    -- CP-element group 112: 	205 
    -- CP-element group 112: 	221 
    -- CP-element group 112: marked-successors 
    -- CP-element group 112: 	110 
    -- CP-element group 112:  members (3) 
      -- CP-element group 112: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_923_Update/$exit
      -- CP-element group 112: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_923_Update/ca
      -- CP-element group 112: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_923_update_completed_
      -- 
    ca_2402_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_923_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(112)); -- 
    -- CP-element group 113:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	42 
    -- CP-element group 113: marked-predecessors 
    -- CP-element group 113: 	115 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_927_sample_start_
      -- CP-element group 113: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_927_Sample/rr
      -- CP-element group 113: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_927_Sample/$entry
      -- 
    rr_2410_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2410_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(113), ack => type_cast_927_inst_req_0); -- 
    zeropad3D_A_cp_element_group_113: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_113"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(42) & zeropad3D_A_CP_1983_elements(115);
      gj_zeropad3D_A_cp_element_group_113 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(113), clk => clk, reset => reset); --
    end block;
    -- CP-element group 114:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: marked-predecessors 
    -- CP-element group 114: 	116 
    -- CP-element group 114: 	127 
    -- CP-element group 114: 	131 
    -- CP-element group 114: 	135 
    -- CP-element group 114: 	143 
    -- CP-element group 114: 	151 
    -- CP-element group 114: 	159 
    -- CP-element group 114: 	167 
    -- CP-element group 114: 	171 
    -- CP-element group 114: 	175 
    -- CP-element group 114: 	179 
    -- CP-element group 114: 	183 
    -- CP-element group 114: 	191 
    -- CP-element group 114: 	207 
    -- CP-element group 114: 	223 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	116 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_927_update_start_
      -- CP-element group 114: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_927_Update/cr
      -- CP-element group 114: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_927_Update/$entry
      -- 
    cr_2415_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2415_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(114), ack => type_cast_927_inst_req_1); -- 
    zeropad3D_A_cp_element_group_114: block -- 
      constant place_capacities: IntegerArray(0 to 14) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1);
      constant place_markings: IntegerArray(0 to 14)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1);
      constant place_delays: IntegerArray(0 to 14) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_114"; 
      signal preds: BooleanArray(1 to 15); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(116) & zeropad3D_A_CP_1983_elements(127) & zeropad3D_A_CP_1983_elements(131) & zeropad3D_A_CP_1983_elements(135) & zeropad3D_A_CP_1983_elements(143) & zeropad3D_A_CP_1983_elements(151) & zeropad3D_A_CP_1983_elements(159) & zeropad3D_A_CP_1983_elements(167) & zeropad3D_A_CP_1983_elements(171) & zeropad3D_A_CP_1983_elements(175) & zeropad3D_A_CP_1983_elements(179) & zeropad3D_A_CP_1983_elements(183) & zeropad3D_A_CP_1983_elements(191) & zeropad3D_A_CP_1983_elements(207) & zeropad3D_A_CP_1983_elements(223);
      gj_zeropad3D_A_cp_element_group_114 : generic_join generic map(name => joinName, number_of_predecessors => 15, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(114), clk => clk, reset => reset); --
    end block;
    -- CP-element group 115:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: successors 
    -- CP-element group 115: marked-successors 
    -- CP-element group 115: 	113 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_927_sample_completed_
      -- CP-element group 115: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_927_Sample/ra
      -- CP-element group 115: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_927_Sample/$exit
      -- 
    ra_2411_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_927_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(115)); -- 
    -- CP-element group 116:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	114 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	125 
    -- CP-element group 116: 	129 
    -- CP-element group 116: 	133 
    -- CP-element group 116: 	141 
    -- CP-element group 116: 	149 
    -- CP-element group 116: 	157 
    -- CP-element group 116: 	165 
    -- CP-element group 116: 	169 
    -- CP-element group 116: 	173 
    -- CP-element group 116: 	177 
    -- CP-element group 116: 	181 
    -- CP-element group 116: 	189 
    -- CP-element group 116: 	205 
    -- CP-element group 116: 	221 
    -- CP-element group 116: marked-successors 
    -- CP-element group 116: 	114 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_927_update_completed_
      -- CP-element group 116: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_927_Update/ca
      -- CP-element group 116: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_927_Update/$exit
      -- 
    ca_2416_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_927_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(116)); -- 
    -- CP-element group 117:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	51 
    -- CP-element group 117: marked-predecessors 
    -- CP-element group 117: 	119 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	119 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_947_Sample/req
      -- CP-element group 117: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_947_Sample/$entry
      -- CP-element group 117: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_947_sample_start_
      -- 
    req_2424_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2424_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(117), ack => W_kx_x1_944_delayed_1_0_945_inst_req_0); -- 
    zeropad3D_A_cp_element_group_117: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_117"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(51) & zeropad3D_A_CP_1983_elements(119);
      gj_zeropad3D_A_cp_element_group_117 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(117), clk => clk, reset => reset); --
    end block;
    -- CP-element group 118:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: marked-predecessors 
    -- CP-element group 118: 	120 
    -- CP-element group 118: 	187 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	120 
    -- CP-element group 118:  members (3) 
      -- CP-element group 118: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_947_Update/$entry
      -- CP-element group 118: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_947_Update/req
      -- CP-element group 118: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_947_update_start_
      -- 
    req_2429_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2429_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(118), ack => W_kx_x1_944_delayed_1_0_945_inst_req_1); -- 
    zeropad3D_A_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(120) & zeropad3D_A_CP_1983_elements(187);
      gj_zeropad3D_A_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	117 
    -- CP-element group 119: successors 
    -- CP-element group 119: marked-successors 
    -- CP-element group 119: 	49 
    -- CP-element group 119: 	117 
    -- CP-element group 119:  members (3) 
      -- CP-element group 119: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_947_Sample/ack
      -- CP-element group 119: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_947_sample_completed_
      -- CP-element group 119: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_947_Sample/$exit
      -- 
    ack_2425_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_kx_x1_944_delayed_1_0_945_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(119)); -- 
    -- CP-element group 120:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	118 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	185 
    -- CP-element group 120: marked-successors 
    -- CP-element group 120: 	118 
    -- CP-element group 120:  members (3) 
      -- CP-element group 120: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_947_Update/$exit
      -- CP-element group 120: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_947_Update/ack
      -- CP-element group 120: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_947_update_completed_
      -- 
    ack_2430_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_kx_x1_944_delayed_1_0_945_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(120)); -- 
    -- CP-element group 121:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	93 
    -- CP-element group 121: marked-predecessors 
    -- CP-element group 121: 	123 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	123 
    -- CP-element group 121:  members (3) 
      -- CP-element group 121: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_963_Sample/req
      -- CP-element group 121: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_963_Sample/$entry
      -- CP-element group 121: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_963_sample_start_
      -- 
    req_2438_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2438_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(121), ack => W_jx_x1_957_delayed_1_0_961_inst_req_0); -- 
    zeropad3D_A_cp_element_group_121: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_121"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(93) & zeropad3D_A_CP_1983_elements(123);
      gj_zeropad3D_A_cp_element_group_121 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(121), clk => clk, reset => reset); --
    end block;
    -- CP-element group 122:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: marked-predecessors 
    -- CP-element group 122: 	124 
    -- CP-element group 122: 	127 
    -- CP-element group 122: 	155 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	124 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_963_Update/$entry
      -- CP-element group 122: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_963_update_start_
      -- CP-element group 122: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_963_Update/req
      -- 
    req_2443_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2443_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(122), ack => W_jx_x1_957_delayed_1_0_961_inst_req_1); -- 
    zeropad3D_A_cp_element_group_122: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_122"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(124) & zeropad3D_A_CP_1983_elements(127) & zeropad3D_A_CP_1983_elements(155);
      gj_zeropad3D_A_cp_element_group_122 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(122), clk => clk, reset => reset); --
    end block;
    -- CP-element group 123:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	121 
    -- CP-element group 123: successors 
    -- CP-element group 123: marked-successors 
    -- CP-element group 123: 	89 
    -- CP-element group 123: 	121 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_963_Sample/ack
      -- CP-element group 123: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_963_Sample/$exit
      -- CP-element group 123: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_963_sample_completed_
      -- 
    ack_2439_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_jx_x1_957_delayed_1_0_961_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(123)); -- 
    -- CP-element group 124:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	122 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	125 
    -- CP-element group 124: 	153 
    -- CP-element group 124: marked-successors 
    -- CP-element group 124: 	122 
    -- CP-element group 124:  members (3) 
      -- CP-element group 124: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_963_Update/$exit
      -- CP-element group 124: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_963_update_completed_
      -- CP-element group 124: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_963_Update/ack
      -- 
    ack_2444_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_jx_x1_957_delayed_1_0_961_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(124)); -- 
    -- CP-element group 125:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	112 
    -- CP-element group 125: 	116 
    -- CP-element group 125: 	124 
    -- CP-element group 125: marked-predecessors 
    -- CP-element group 125: 	127 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	127 
    -- CP-element group 125:  members (3) 
      -- CP-element group 125: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_974_Sample/rr
      -- CP-element group 125: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_974_Sample/$entry
      -- CP-element group 125: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_974_sample_start_
      -- 
    rr_2452_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2452_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(125), ack => type_cast_974_inst_req_0); -- 
    zeropad3D_A_cp_element_group_125: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_125"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(112) & zeropad3D_A_CP_1983_elements(116) & zeropad3D_A_CP_1983_elements(124) & zeropad3D_A_CP_1983_elements(127);
      gj_zeropad3D_A_cp_element_group_125 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(125), clk => clk, reset => reset); --
    end block;
    -- CP-element group 126:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: marked-predecessors 
    -- CP-element group 126: 	128 
    -- CP-element group 126: 	139 
    -- CP-element group 126: 	215 
    -- CP-element group 126: 	219 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	128 
    -- CP-element group 126:  members (3) 
      -- CP-element group 126: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_974_Update/$entry
      -- CP-element group 126: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_974_Update/cr
      -- CP-element group 126: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_974_update_start_
      -- 
    cr_2457_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2457_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(126), ack => type_cast_974_inst_req_1); -- 
    zeropad3D_A_cp_element_group_126: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_126"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(128) & zeropad3D_A_CP_1983_elements(139) & zeropad3D_A_CP_1983_elements(215) & zeropad3D_A_CP_1983_elements(219);
      gj_zeropad3D_A_cp_element_group_126 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(126), clk => clk, reset => reset); --
    end block;
    -- CP-element group 127:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	125 
    -- CP-element group 127: successors 
    -- CP-element group 127: marked-successors 
    -- CP-element group 127: 	110 
    -- CP-element group 127: 	114 
    -- CP-element group 127: 	122 
    -- CP-element group 127: 	125 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_974_Sample/ra
      -- CP-element group 127: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_974_Sample/$exit
      -- CP-element group 127: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_974_sample_completed_
      -- 
    ra_2453_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_974_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(127)); -- 
    -- CP-element group 128:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	126 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	137 
    -- CP-element group 128: 	213 
    -- CP-element group 128: 	217 
    -- CP-element group 128: marked-successors 
    -- CP-element group 128: 	126 
    -- CP-element group 128:  members (3) 
      -- CP-element group 128: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_974_Update/$exit
      -- CP-element group 128: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_974_Update/ca
      -- CP-element group 128: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_974_update_completed_
      -- 
    ca_2458_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_974_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(128)); -- 
    -- CP-element group 129:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	112 
    -- CP-element group 129: 	116 
    -- CP-element group 129: marked-predecessors 
    -- CP-element group 129: 	131 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	131 
    -- CP-element group 129:  members (3) 
      -- CP-element group 129: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_978_Sample/$entry
      -- CP-element group 129: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_978_Sample/req
      -- CP-element group 129: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_978_sample_start_
      -- 
    req_2466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(129), ack => W_ifx_xelse_exec_guard_967_delayed_1_0_976_inst_req_0); -- 
    zeropad3D_A_cp_element_group_129: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_129"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(112) & zeropad3D_A_CP_1983_elements(116) & zeropad3D_A_CP_1983_elements(131);
      gj_zeropad3D_A_cp_element_group_129 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(129), clk => clk, reset => reset); --
    end block;
    -- CP-element group 130:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: marked-predecessors 
    -- CP-element group 130: 	132 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	132 
    -- CP-element group 130:  members (3) 
      -- CP-element group 130: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_978_Update/$entry
      -- CP-element group 130: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_978_update_start_
      -- CP-element group 130: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_978_Update/req
      -- 
    req_2471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(130), ack => W_ifx_xelse_exec_guard_967_delayed_1_0_976_inst_req_1); -- 
    zeropad3D_A_cp_element_group_130: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_130"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= zeropad3D_A_CP_1983_elements(132);
      gj_zeropad3D_A_cp_element_group_130 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(130), clk => clk, reset => reset); --
    end block;
    -- CP-element group 131:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	129 
    -- CP-element group 131: successors 
    -- CP-element group 131: marked-successors 
    -- CP-element group 131: 	110 
    -- CP-element group 131: 	114 
    -- CP-element group 131: 	129 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_978_Sample/ack
      -- CP-element group 131: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_978_Sample/$exit
      -- CP-element group 131: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_978_sample_completed_
      -- 
    ack_2467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xelse_exec_guard_967_delayed_1_0_976_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(131)); -- 
    -- CP-element group 132:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	130 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	404 
    -- CP-element group 132: marked-successors 
    -- CP-element group 132: 	130 
    -- CP-element group 132:  members (3) 
      -- CP-element group 132: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_978_Update/$exit
      -- CP-element group 132: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_978_Update/ack
      -- CP-element group 132: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_978_update_completed_
      -- 
    ack_2472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xelse_exec_guard_967_delayed_1_0_976_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(132)); -- 
    -- CP-element group 133:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	112 
    -- CP-element group 133: 	116 
    -- CP-element group 133: marked-predecessors 
    -- CP-element group 133: 	135 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	135 
    -- CP-element group 133:  members (3) 
      -- CP-element group 133: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_987_Sample/req
      -- CP-element group 133: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_987_Sample/$entry
      -- CP-element group 133: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_987_sample_start_
      -- 
    req_2480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(133), ack => W_ifx_xelse_exec_guard_973_delayed_1_0_985_inst_req_0); -- 
    zeropad3D_A_cp_element_group_133: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_133"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(112) & zeropad3D_A_CP_1983_elements(116) & zeropad3D_A_CP_1983_elements(135);
      gj_zeropad3D_A_cp_element_group_133 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(133), clk => clk, reset => reset); --
    end block;
    -- CP-element group 134:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: marked-predecessors 
    -- CP-element group 134: 	136 
    -- CP-element group 134: 	139 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	136 
    -- CP-element group 134:  members (3) 
      -- CP-element group 134: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_987_Update/$entry
      -- CP-element group 134: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_987_Update/req
      -- CP-element group 134: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_987_update_start_
      -- 
    req_2485_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2485_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(134), ack => W_ifx_xelse_exec_guard_973_delayed_1_0_985_inst_req_1); -- 
    zeropad3D_A_cp_element_group_134: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_134"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(136) & zeropad3D_A_CP_1983_elements(139);
      gj_zeropad3D_A_cp_element_group_134 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(134), clk => clk, reset => reset); --
    end block;
    -- CP-element group 135:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	133 
    -- CP-element group 135: successors 
    -- CP-element group 135: marked-successors 
    -- CP-element group 135: 	110 
    -- CP-element group 135: 	114 
    -- CP-element group 135: 	133 
    -- CP-element group 135:  members (3) 
      -- CP-element group 135: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_987_Sample/ack
      -- CP-element group 135: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_987_Sample/$exit
      -- CP-element group 135: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_987_sample_completed_
      -- 
    ack_2481_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xelse_exec_guard_973_delayed_1_0_985_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(135)); -- 
    -- CP-element group 136:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	134 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	137 
    -- CP-element group 136: marked-successors 
    -- CP-element group 136: 	134 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_987_Update/$exit
      -- CP-element group 136: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_987_Update/ack
      -- CP-element group 136: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_987_update_completed_
      -- 
    ack_2486_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xelse_exec_guard_973_delayed_1_0_985_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(136)); -- 
    -- CP-element group 137:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	128 
    -- CP-element group 137: 	136 
    -- CP-element group 137: marked-predecessors 
    -- CP-element group 137: 	139 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	139 
    -- CP-element group 137:  members (3) 
      -- CP-element group 137: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_991_sample_start_
      -- CP-element group 137: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_991_Sample/$entry
      -- CP-element group 137: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_991_Sample/rr
      -- 
    rr_2494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(137), ack => type_cast_991_inst_req_0); -- 
    zeropad3D_A_cp_element_group_137: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_137"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(128) & zeropad3D_A_CP_1983_elements(136) & zeropad3D_A_CP_1983_elements(139);
      gj_zeropad3D_A_cp_element_group_137 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(137), clk => clk, reset => reset); --
    end block;
    -- CP-element group 138:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: marked-predecessors 
    -- CP-element group 138: 	140 
    -- CP-element group 138: 	163 
    -- CP-element group 138: 	199 
    -- CP-element group 138: 	203 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	140 
    -- CP-element group 138:  members (3) 
      -- CP-element group 138: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_991_update_start_
      -- CP-element group 138: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_991_Update/$entry
      -- CP-element group 138: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_991_Update/cr
      -- 
    cr_2499_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2499_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(138), ack => type_cast_991_inst_req_1); -- 
    zeropad3D_A_cp_element_group_138: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_138"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(140) & zeropad3D_A_CP_1983_elements(163) & zeropad3D_A_CP_1983_elements(199) & zeropad3D_A_CP_1983_elements(203);
      gj_zeropad3D_A_cp_element_group_138 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(138), clk => clk, reset => reset); --
    end block;
    -- CP-element group 139:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	137 
    -- CP-element group 139: successors 
    -- CP-element group 139: marked-successors 
    -- CP-element group 139: 	126 
    -- CP-element group 139: 	134 
    -- CP-element group 139: 	137 
    -- CP-element group 139:  members (3) 
      -- CP-element group 139: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_991_sample_completed_
      -- CP-element group 139: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_991_Sample/$exit
      -- CP-element group 139: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_991_Sample/ra
      -- 
    ra_2495_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_991_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(139)); -- 
    -- CP-element group 140:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	138 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	161 
    -- CP-element group 140: 	197 
    -- CP-element group 140: 	201 
    -- CP-element group 140: marked-successors 
    -- CP-element group 140: 	138 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_991_Update/ca
      -- CP-element group 140: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_991_update_completed_
      -- CP-element group 140: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_991_Update/$exit
      -- 
    ca_2500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_991_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(140)); -- 
    -- CP-element group 141:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	112 
    -- CP-element group 141: 	116 
    -- CP-element group 141: marked-predecessors 
    -- CP-element group 141: 	143 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	143 
    -- CP-element group 141:  members (3) 
      -- CP-element group 141: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_995_Sample/$entry
      -- CP-element group 141: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_995_Sample/req
      -- CP-element group 141: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_995_sample_start_
      -- 
    req_2508_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2508_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(141), ack => W_ifx_xelse_exec_guard_978_delayed_2_0_993_inst_req_0); -- 
    zeropad3D_A_cp_element_group_141: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_141"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(112) & zeropad3D_A_CP_1983_elements(116) & zeropad3D_A_CP_1983_elements(143);
      gj_zeropad3D_A_cp_element_group_141 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(141), clk => clk, reset => reset); --
    end block;
    -- CP-element group 142:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: marked-predecessors 
    -- CP-element group 142: 	144 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	144 
    -- CP-element group 142:  members (3) 
      -- CP-element group 142: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_995_Update/$entry
      -- CP-element group 142: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_995_Update/req
      -- CP-element group 142: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_995_update_start_
      -- 
    req_2513_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2513_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(142), ack => W_ifx_xelse_exec_guard_978_delayed_2_0_993_inst_req_1); -- 
    zeropad3D_A_cp_element_group_142: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_142"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= zeropad3D_A_CP_1983_elements(144);
      gj_zeropad3D_A_cp_element_group_142 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(142), clk => clk, reset => reset); --
    end block;
    -- CP-element group 143:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	141 
    -- CP-element group 143: successors 
    -- CP-element group 143: marked-successors 
    -- CP-element group 143: 	110 
    -- CP-element group 143: 	114 
    -- CP-element group 143: 	141 
    -- CP-element group 143:  members (3) 
      -- CP-element group 143: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_995_sample_completed_
      -- CP-element group 143: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_995_Sample/$exit
      -- CP-element group 143: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_995_Sample/ack
      -- 
    ack_2509_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xelse_exec_guard_978_delayed_2_0_993_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(143)); -- 
    -- CP-element group 144:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	142 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	404 
    -- CP-element group 144: marked-successors 
    -- CP-element group 144: 	142 
    -- CP-element group 144:  members (3) 
      -- CP-element group 144: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_995_update_completed_
      -- CP-element group 144: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_995_Update/ack
      -- CP-element group 144: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_995_Update/$exit
      -- 
    ack_2514_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xelse_exec_guard_978_delayed_2_0_993_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(144)); -- 
    -- CP-element group 145:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	72 
    -- CP-element group 145: marked-predecessors 
    -- CP-element group 145: 	147 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	147 
    -- CP-element group 145:  members (3) 
      -- CP-element group 145: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_998_sample_start_
      -- CP-element group 145: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_998_Sample/$entry
      -- CP-element group 145: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_998_Sample/req
      -- 
    req_2522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(145), ack => W_ix_x2_981_delayed_3_0_996_inst_req_0); -- 
    zeropad3D_A_cp_element_group_145: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_145"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(72) & zeropad3D_A_CP_1983_elements(147);
      gj_zeropad3D_A_cp_element_group_145 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(145), clk => clk, reset => reset); --
    end block;
    -- CP-element group 146:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: marked-predecessors 
    -- CP-element group 146: 	148 
    -- CP-element group 146: 	163 
    -- CP-element group 146: 	199 
    -- CP-element group 146: 	203 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	148 
    -- CP-element group 146:  members (3) 
      -- CP-element group 146: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_998_update_start_
      -- CP-element group 146: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_998_Update/$entry
      -- CP-element group 146: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_998_Update/req
      -- 
    req_2527_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2527_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(146), ack => W_ix_x2_981_delayed_3_0_996_inst_req_1); -- 
    zeropad3D_A_cp_element_group_146: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_146"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(148) & zeropad3D_A_CP_1983_elements(163) & zeropad3D_A_CP_1983_elements(199) & zeropad3D_A_CP_1983_elements(203);
      gj_zeropad3D_A_cp_element_group_146 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(146), clk => clk, reset => reset); --
    end block;
    -- CP-element group 147:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	145 
    -- CP-element group 147: successors 
    -- CP-element group 147: marked-successors 
    -- CP-element group 147: 	68 
    -- CP-element group 147: 	145 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_998_sample_completed_
      -- CP-element group 147: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_998_Sample/$exit
      -- CP-element group 147: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_998_Sample/ack
      -- 
    ack_2523_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ix_x2_981_delayed_3_0_996_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(147)); -- 
    -- CP-element group 148:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	146 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	161 
    -- CP-element group 148: 	197 
    -- CP-element group 148: 	201 
    -- CP-element group 148: marked-successors 
    -- CP-element group 148: 	146 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_998_update_completed_
      -- CP-element group 148: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_998_Update/$exit
      -- CP-element group 148: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_998_Update/ack
      -- 
    ack_2528_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ix_x2_981_delayed_3_0_996_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(148)); -- 
    -- CP-element group 149:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	112 
    -- CP-element group 149: 	116 
    -- CP-element group 149: marked-predecessors 
    -- CP-element group 149: 	151 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	151 
    -- CP-element group 149:  members (3) 
      -- CP-element group 149: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1007_sample_start_
      -- CP-element group 149: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1007_Sample/$entry
      -- CP-element group 149: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1007_Sample/req
      -- 
    req_2536_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2536_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(149), ack => W_ifx_xelse_exec_guard_984_delayed_1_0_1005_inst_req_0); -- 
    zeropad3D_A_cp_element_group_149: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_149"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(112) & zeropad3D_A_CP_1983_elements(116) & zeropad3D_A_CP_1983_elements(151);
      gj_zeropad3D_A_cp_element_group_149 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(149), clk => clk, reset => reset); --
    end block;
    -- CP-element group 150:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: marked-predecessors 
    -- CP-element group 150: 	152 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	152 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1007_update_start_
      -- CP-element group 150: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1007_Update/$entry
      -- CP-element group 150: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1007_Update/req
      -- 
    req_2541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(150), ack => W_ifx_xelse_exec_guard_984_delayed_1_0_1005_inst_req_1); -- 
    zeropad3D_A_cp_element_group_150: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_150"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= zeropad3D_A_CP_1983_elements(152);
      gj_zeropad3D_A_cp_element_group_150 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(150), clk => clk, reset => reset); --
    end block;
    -- CP-element group 151:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	149 
    -- CP-element group 151: successors 
    -- CP-element group 151: marked-successors 
    -- CP-element group 151: 	110 
    -- CP-element group 151: 	114 
    -- CP-element group 151: 	149 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1007_sample_completed_
      -- CP-element group 151: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1007_Sample/$exit
      -- CP-element group 151: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1007_Sample/ack
      -- 
    ack_2537_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xelse_exec_guard_984_delayed_1_0_1005_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(151)); -- 
    -- CP-element group 152:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	150 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	404 
    -- CP-element group 152: marked-successors 
    -- CP-element group 152: 	150 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1007_update_completed_
      -- CP-element group 152: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1007_Update/$exit
      -- CP-element group 152: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1007_Update/ack
      -- 
    ack_2542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xelse_exec_guard_984_delayed_1_0_1005_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(152)); -- 
    -- CP-element group 153:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	124 
    -- CP-element group 153: marked-predecessors 
    -- CP-element group 153: 	155 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	155 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1010_sample_start_
      -- CP-element group 153: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1010_Sample/$entry
      -- CP-element group 153: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1010_Sample/req
      -- 
    req_2550_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2550_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(153), ack => W_inc_989_delayed_1_0_1008_inst_req_0); -- 
    zeropad3D_A_cp_element_group_153: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_153"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(124) & zeropad3D_A_CP_1983_elements(155);
      gj_zeropad3D_A_cp_element_group_153 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(153), clk => clk, reset => reset); --
    end block;
    -- CP-element group 154:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: marked-predecessors 
    -- CP-element group 154: 	156 
    -- CP-element group 154: 	215 
    -- CP-element group 154: 	219 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	156 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1010_update_start_
      -- CP-element group 154: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1010_Update/$entry
      -- CP-element group 154: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1010_Update/req
      -- 
    req_2555_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2555_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(154), ack => W_inc_989_delayed_1_0_1008_inst_req_1); -- 
    zeropad3D_A_cp_element_group_154: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_154"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(156) & zeropad3D_A_CP_1983_elements(215) & zeropad3D_A_CP_1983_elements(219);
      gj_zeropad3D_A_cp_element_group_154 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(154), clk => clk, reset => reset); --
    end block;
    -- CP-element group 155:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	153 
    -- CP-element group 155: successors 
    -- CP-element group 155: marked-successors 
    -- CP-element group 155: 	122 
    -- CP-element group 155: 	153 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1010_sample_completed_
      -- CP-element group 155: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1010_Sample/$exit
      -- CP-element group 155: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1010_Sample/ack
      -- 
    ack_2551_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_inc_989_delayed_1_0_1008_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(155)); -- 
    -- CP-element group 156:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	154 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	213 
    -- CP-element group 156: 	217 
    -- CP-element group 156: marked-successors 
    -- CP-element group 156: 	154 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1010_update_completed_
      -- CP-element group 156: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1010_Update/$exit
      -- CP-element group 156: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1010_Update/ack
      -- 
    ack_2556_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_inc_989_delayed_1_0_1008_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(156)); -- 
    -- CP-element group 157:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	112 
    -- CP-element group 157: 	116 
    -- CP-element group 157: marked-predecessors 
    -- CP-element group 157: 	159 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	159 
    -- CP-element group 157:  members (3) 
      -- CP-element group 157: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1021_sample_start_
      -- CP-element group 157: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1021_Sample/$entry
      -- CP-element group 157: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1021_Sample/req
      -- 
    req_2564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(157), ack => W_ifx_xelse_exec_guard_992_delayed_2_0_1019_inst_req_0); -- 
    zeropad3D_A_cp_element_group_157: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_157"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(112) & zeropad3D_A_CP_1983_elements(116) & zeropad3D_A_CP_1983_elements(159);
      gj_zeropad3D_A_cp_element_group_157 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(157), clk => clk, reset => reset); --
    end block;
    -- CP-element group 158:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: marked-predecessors 
    -- CP-element group 158: 	160 
    -- CP-element group 158: 	163 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	160 
    -- CP-element group 158:  members (3) 
      -- CP-element group 158: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1021_update_start_
      -- CP-element group 158: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1021_Update/$entry
      -- CP-element group 158: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1021_Update/req
      -- 
    req_2569_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2569_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(158), ack => W_ifx_xelse_exec_guard_992_delayed_2_0_1019_inst_req_1); -- 
    zeropad3D_A_cp_element_group_158: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_158"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(160) & zeropad3D_A_CP_1983_elements(163);
      gj_zeropad3D_A_cp_element_group_158 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(158), clk => clk, reset => reset); --
    end block;
    -- CP-element group 159:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	157 
    -- CP-element group 159: successors 
    -- CP-element group 159: marked-successors 
    -- CP-element group 159: 	110 
    -- CP-element group 159: 	114 
    -- CP-element group 159: 	157 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1021_sample_completed_
      -- CP-element group 159: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1021_Sample/$exit
      -- CP-element group 159: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1021_Sample/ack
      -- 
    ack_2565_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xelse_exec_guard_992_delayed_2_0_1019_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(159)); -- 
    -- CP-element group 160:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	158 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	161 
    -- CP-element group 160: marked-successors 
    -- CP-element group 160: 	158 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1021_update_completed_
      -- CP-element group 160: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1021_Update/$exit
      -- CP-element group 160: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1021_Update/ack
      -- 
    ack_2570_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xelse_exec_guard_992_delayed_2_0_1019_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(160)); -- 
    -- CP-element group 161:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	140 
    -- CP-element group 161: 	148 
    -- CP-element group 161: 	160 
    -- CP-element group 161: marked-predecessors 
    -- CP-element group 161: 	163 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	163 
    -- CP-element group 161:  members (3) 
      -- CP-element group 161: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1025_sample_start_
      -- CP-element group 161: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1025_Sample/$entry
      -- CP-element group 161: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1025_Sample/rr
      -- 
    rr_2578_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2578_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(161), ack => type_cast_1025_inst_req_0); -- 
    zeropad3D_A_cp_element_group_161: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_161"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(140) & zeropad3D_A_CP_1983_elements(148) & zeropad3D_A_CP_1983_elements(160) & zeropad3D_A_CP_1983_elements(163);
      gj_zeropad3D_A_cp_element_group_161 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(161), clk => clk, reset => reset); --
    end block;
    -- CP-element group 162:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	45 
    -- CP-element group 162: marked-predecessors 
    -- CP-element group 162: 	164 
    -- CP-element group 162: 	227 
    -- CP-element group 162: 	231 
    -- CP-element group 162: 	235 
    -- CP-element group 162: 	239 
    -- CP-element group 162: 	247 
    -- CP-element group 162: 	251 
    -- CP-element group 162: 	255 
    -- CP-element group 162: 	259 
    -- CP-element group 162: 	299 
    -- CP-element group 162: 	330 
    -- CP-element group 162: 	365 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	164 
    -- CP-element group 162:  members (3) 
      -- CP-element group 162: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1025_update_start_
      -- CP-element group 162: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1025_Update/$entry
      -- CP-element group 162: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1025_Update/cr
      -- 
    cr_2583_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2583_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(162), ack => type_cast_1025_inst_req_1); -- 
    zeropad3D_A_cp_element_group_162: block -- 
      constant place_capacities: IntegerArray(0 to 12) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1);
      constant place_markings: IntegerArray(0 to 12)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1);
      constant place_delays: IntegerArray(0 to 12) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_162"; 
      signal preds: BooleanArray(1 to 13); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(45) & zeropad3D_A_CP_1983_elements(164) & zeropad3D_A_CP_1983_elements(227) & zeropad3D_A_CP_1983_elements(231) & zeropad3D_A_CP_1983_elements(235) & zeropad3D_A_CP_1983_elements(239) & zeropad3D_A_CP_1983_elements(247) & zeropad3D_A_CP_1983_elements(251) & zeropad3D_A_CP_1983_elements(255) & zeropad3D_A_CP_1983_elements(259) & zeropad3D_A_CP_1983_elements(299) & zeropad3D_A_CP_1983_elements(330) & zeropad3D_A_CP_1983_elements(365);
      gj_zeropad3D_A_cp_element_group_162 : generic_join generic map(name => joinName, number_of_predecessors => 13, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(162), clk => clk, reset => reset); --
    end block;
    -- CP-element group 163:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	161 
    -- CP-element group 163: successors 
    -- CP-element group 163: marked-successors 
    -- CP-element group 163: 	138 
    -- CP-element group 163: 	146 
    -- CP-element group 163: 	158 
    -- CP-element group 163: 	161 
    -- CP-element group 163:  members (3) 
      -- CP-element group 163: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1025_sample_completed_
      -- CP-element group 163: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1025_Sample/$exit
      -- CP-element group 163: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1025_Sample/ra
      -- 
    ra_2579_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1025_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(163)); -- 
    -- CP-element group 164:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	162 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	43 
    -- CP-element group 164: 	225 
    -- CP-element group 164: 	229 
    -- CP-element group 164: 	233 
    -- CP-element group 164: 	237 
    -- CP-element group 164: 	245 
    -- CP-element group 164: 	249 
    -- CP-element group 164: 	253 
    -- CP-element group 164: 	257 
    -- CP-element group 164: 	297 
    -- CP-element group 164: 	328 
    -- CP-element group 164: 	363 
    -- CP-element group 164: marked-successors 
    -- CP-element group 164: 	48 
    -- CP-element group 164: 	67 
    -- CP-element group 164: 	88 
    -- CP-element group 164: 	162 
    -- CP-element group 164:  members (3) 
      -- CP-element group 164: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1025_update_completed_
      -- CP-element group 164: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1025_Update/$exit
      -- CP-element group 164: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1025_Update/ca
      -- 
    ca_2584_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1025_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(164)); -- 
    -- CP-element group 165:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	112 
    -- CP-element group 165: 	116 
    -- CP-element group 165: marked-predecessors 
    -- CP-element group 165: 	167 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	167 
    -- CP-element group 165:  members (3) 
      -- CP-element group 165: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1029_sample_start_
      -- CP-element group 165: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1029_Sample/$entry
      -- CP-element group 165: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1029_Sample/req
      -- 
    req_2592_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2592_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(165), ack => W_ifx_xelse_exec_guard_997_delayed_3_0_1027_inst_req_0); -- 
    zeropad3D_A_cp_element_group_165: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_165"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(112) & zeropad3D_A_CP_1983_elements(116) & zeropad3D_A_CP_1983_elements(167);
      gj_zeropad3D_A_cp_element_group_165 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(165), clk => clk, reset => reset); --
    end block;
    -- CP-element group 166:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: marked-predecessors 
    -- CP-element group 166: 	168 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	168 
    -- CP-element group 166:  members (3) 
      -- CP-element group 166: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1029_update_start_
      -- CP-element group 166: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1029_Update/$entry
      -- CP-element group 166: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1029_Update/req
      -- 
    req_2597_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2597_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(166), ack => W_ifx_xelse_exec_guard_997_delayed_3_0_1027_inst_req_1); -- 
    zeropad3D_A_cp_element_group_166: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_166"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= zeropad3D_A_CP_1983_elements(168);
      gj_zeropad3D_A_cp_element_group_166 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(166), clk => clk, reset => reset); --
    end block;
    -- CP-element group 167:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	165 
    -- CP-element group 167: successors 
    -- CP-element group 167: marked-successors 
    -- CP-element group 167: 	110 
    -- CP-element group 167: 	114 
    -- CP-element group 167: 	165 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1029_sample_completed_
      -- CP-element group 167: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1029_Sample/$exit
      -- CP-element group 167: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1029_Sample/ack
      -- 
    ack_2593_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xelse_exec_guard_997_delayed_3_0_1027_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(167)); -- 
    -- CP-element group 168:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	166 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	404 
    -- CP-element group 168: marked-successors 
    -- CP-element group 168: 	166 
    -- CP-element group 168:  members (3) 
      -- CP-element group 168: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1029_update_completed_
      -- CP-element group 168: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1029_Update/$exit
      -- CP-element group 168: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1029_Update/ack
      -- 
    ack_2598_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xelse_exec_guard_997_delayed_3_0_1027_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(168)); -- 
    -- CP-element group 169:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	112 
    -- CP-element group 169: 	116 
    -- CP-element group 169: marked-predecessors 
    -- CP-element group 169: 	171 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	171 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1038_sample_start_
      -- CP-element group 169: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1038_Sample/$entry
      -- CP-element group 169: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1038_Sample/req
      -- 
    req_2606_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2606_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(169), ack => W_ifx_xelse_exec_guard_1004_delayed_3_0_1036_inst_req_0); -- 
    zeropad3D_A_cp_element_group_169: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_169"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(112) & zeropad3D_A_CP_1983_elements(116) & zeropad3D_A_CP_1983_elements(171);
      gj_zeropad3D_A_cp_element_group_169 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(169), clk => clk, reset => reset); --
    end block;
    -- CP-element group 170:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	45 
    -- CP-element group 170: marked-predecessors 
    -- CP-element group 170: 	172 
    -- CP-element group 170: 	227 
    -- CP-element group 170: 	231 
    -- CP-element group 170: 	235 
    -- CP-element group 170: 	239 
    -- CP-element group 170: 	247 
    -- CP-element group 170: 	251 
    -- CP-element group 170: 	255 
    -- CP-element group 170: 	259 
    -- CP-element group 170: 	299 
    -- CP-element group 170: 	330 
    -- CP-element group 170: 	365 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	172 
    -- CP-element group 170:  members (3) 
      -- CP-element group 170: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1038_update_start_
      -- CP-element group 170: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1038_Update/$entry
      -- CP-element group 170: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1038_Update/req
      -- 
    req_2611_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2611_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(170), ack => W_ifx_xelse_exec_guard_1004_delayed_3_0_1036_inst_req_1); -- 
    zeropad3D_A_cp_element_group_170: block -- 
      constant place_capacities: IntegerArray(0 to 12) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1);
      constant place_markings: IntegerArray(0 to 12)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1);
      constant place_delays: IntegerArray(0 to 12) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_170"; 
      signal preds: BooleanArray(1 to 13); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(45) & zeropad3D_A_CP_1983_elements(172) & zeropad3D_A_CP_1983_elements(227) & zeropad3D_A_CP_1983_elements(231) & zeropad3D_A_CP_1983_elements(235) & zeropad3D_A_CP_1983_elements(239) & zeropad3D_A_CP_1983_elements(247) & zeropad3D_A_CP_1983_elements(251) & zeropad3D_A_CP_1983_elements(255) & zeropad3D_A_CP_1983_elements(259) & zeropad3D_A_CP_1983_elements(299) & zeropad3D_A_CP_1983_elements(330) & zeropad3D_A_CP_1983_elements(365);
      gj_zeropad3D_A_cp_element_group_170 : generic_join generic map(name => joinName, number_of_predecessors => 13, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(170), clk => clk, reset => reset); --
    end block;
    -- CP-element group 171:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	169 
    -- CP-element group 171: successors 
    -- CP-element group 171: marked-successors 
    -- CP-element group 171: 	110 
    -- CP-element group 171: 	114 
    -- CP-element group 171: 	169 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1038_sample_completed_
      -- CP-element group 171: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1038_Sample/$exit
      -- CP-element group 171: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1038_Sample/ack
      -- 
    ack_2607_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xelse_exec_guard_1004_delayed_3_0_1036_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(171)); -- 
    -- CP-element group 172:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	170 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	43 
    -- CP-element group 172: 	225 
    -- CP-element group 172: 	229 
    -- CP-element group 172: 	233 
    -- CP-element group 172: 	237 
    -- CP-element group 172: 	245 
    -- CP-element group 172: 	249 
    -- CP-element group 172: 	253 
    -- CP-element group 172: 	257 
    -- CP-element group 172: 	297 
    -- CP-element group 172: 	328 
    -- CP-element group 172: 	363 
    -- CP-element group 172: marked-successors 
    -- CP-element group 172: 	48 
    -- CP-element group 172: 	67 
    -- CP-element group 172: 	88 
    -- CP-element group 172: 	170 
    -- CP-element group 172:  members (3) 
      -- CP-element group 172: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1038_update_completed_
      -- CP-element group 172: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1038_Update/$exit
      -- CP-element group 172: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1038_Update/ack
      -- 
    ack_2612_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xelse_exec_guard_1004_delayed_3_0_1036_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(172)); -- 
    -- CP-element group 173:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	112 
    -- CP-element group 173: 	116 
    -- CP-element group 173: marked-predecessors 
    -- CP-element group 173: 	175 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	175 
    -- CP-element group 173:  members (3) 
      -- CP-element group 173: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1046_sample_start_
      -- CP-element group 173: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1046_Sample/$entry
      -- CP-element group 173: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1046_Sample/req
      -- 
    req_2620_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2620_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(173), ack => W_ifx_xelse_exec_guard_1009_delayed_3_0_1044_inst_req_0); -- 
    zeropad3D_A_cp_element_group_173: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_173"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(112) & zeropad3D_A_CP_1983_elements(116) & zeropad3D_A_CP_1983_elements(175);
      gj_zeropad3D_A_cp_element_group_173 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(173), clk => clk, reset => reset); --
    end block;
    -- CP-element group 174:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	45 
    -- CP-element group 174: marked-predecessors 
    -- CP-element group 174: 	176 
    -- CP-element group 174: 	227 
    -- CP-element group 174: 	231 
    -- CP-element group 174: 	235 
    -- CP-element group 174: 	239 
    -- CP-element group 174: 	247 
    -- CP-element group 174: 	251 
    -- CP-element group 174: 	255 
    -- CP-element group 174: 	259 
    -- CP-element group 174: 	299 
    -- CP-element group 174: 	330 
    -- CP-element group 174: 	365 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	176 
    -- CP-element group 174:  members (3) 
      -- CP-element group 174: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1046_update_start_
      -- CP-element group 174: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1046_Update/$entry
      -- CP-element group 174: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1046_Update/req
      -- 
    req_2625_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2625_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(174), ack => W_ifx_xelse_exec_guard_1009_delayed_3_0_1044_inst_req_1); -- 
    zeropad3D_A_cp_element_group_174: block -- 
      constant place_capacities: IntegerArray(0 to 12) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1);
      constant place_markings: IntegerArray(0 to 12)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1);
      constant place_delays: IntegerArray(0 to 12) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_174"; 
      signal preds: BooleanArray(1 to 13); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(45) & zeropad3D_A_CP_1983_elements(176) & zeropad3D_A_CP_1983_elements(227) & zeropad3D_A_CP_1983_elements(231) & zeropad3D_A_CP_1983_elements(235) & zeropad3D_A_CP_1983_elements(239) & zeropad3D_A_CP_1983_elements(247) & zeropad3D_A_CP_1983_elements(251) & zeropad3D_A_CP_1983_elements(255) & zeropad3D_A_CP_1983_elements(259) & zeropad3D_A_CP_1983_elements(299) & zeropad3D_A_CP_1983_elements(330) & zeropad3D_A_CP_1983_elements(365);
      gj_zeropad3D_A_cp_element_group_174 : generic_join generic map(name => joinName, number_of_predecessors => 13, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(174), clk => clk, reset => reset); --
    end block;
    -- CP-element group 175:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	173 
    -- CP-element group 175: successors 
    -- CP-element group 175: marked-successors 
    -- CP-element group 175: 	110 
    -- CP-element group 175: 	114 
    -- CP-element group 175: 	173 
    -- CP-element group 175:  members (3) 
      -- CP-element group 175: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1046_sample_completed_
      -- CP-element group 175: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1046_Sample/$exit
      -- CP-element group 175: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1046_Sample/ack
      -- 
    ack_2621_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xelse_exec_guard_1009_delayed_3_0_1044_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(175)); -- 
    -- CP-element group 176:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	174 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	43 
    -- CP-element group 176: 	225 
    -- CP-element group 176: 	229 
    -- CP-element group 176: 	233 
    -- CP-element group 176: 	237 
    -- CP-element group 176: 	245 
    -- CP-element group 176: 	249 
    -- CP-element group 176: 	253 
    -- CP-element group 176: 	257 
    -- CP-element group 176: 	297 
    -- CP-element group 176: 	328 
    -- CP-element group 176: 	363 
    -- CP-element group 176: marked-successors 
    -- CP-element group 176: 	48 
    -- CP-element group 176: 	67 
    -- CP-element group 176: 	88 
    -- CP-element group 176: 	174 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1046_update_completed_
      -- CP-element group 176: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1046_Update/$exit
      -- CP-element group 176: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1046_Update/ack
      -- 
    ack_2626_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xelse_exec_guard_1009_delayed_3_0_1044_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(176)); -- 
    -- CP-element group 177:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	112 
    -- CP-element group 177: 	116 
    -- CP-element group 177: marked-predecessors 
    -- CP-element group 177: 	179 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	179 
    -- CP-element group 177:  members (3) 
      -- CP-element group 177: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1061_sample_start_
      -- CP-element group 177: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1061_Sample/$entry
      -- CP-element group 177: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1061_Sample/req
      -- 
    req_2634_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2634_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(177), ack => W_ifx_xthen_ifx_xend80_taken_1022_delayed_3_0_1059_inst_req_0); -- 
    zeropad3D_A_cp_element_group_177: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_177"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(112) & zeropad3D_A_CP_1983_elements(116) & zeropad3D_A_CP_1983_elements(179);
      gj_zeropad3D_A_cp_element_group_177 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(177), clk => clk, reset => reset); --
    end block;
    -- CP-element group 178:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: marked-predecessors 
    -- CP-element group 178: 	180 
    -- CP-element group 178: 	227 
    -- CP-element group 178: 	231 
    -- CP-element group 178: 	235 
    -- CP-element group 178: 	239 
    -- CP-element group 178: 	247 
    -- CP-element group 178: 	251 
    -- CP-element group 178: 	255 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	180 
    -- CP-element group 178:  members (3) 
      -- CP-element group 178: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1061_update_start_
      -- CP-element group 178: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1061_Update/$entry
      -- CP-element group 178: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1061_Update/req
      -- 
    req_2639_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2639_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(178), ack => W_ifx_xthen_ifx_xend80_taken_1022_delayed_3_0_1059_inst_req_1); -- 
    zeropad3D_A_cp_element_group_178: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_178"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(180) & zeropad3D_A_CP_1983_elements(227) & zeropad3D_A_CP_1983_elements(231) & zeropad3D_A_CP_1983_elements(235) & zeropad3D_A_CP_1983_elements(239) & zeropad3D_A_CP_1983_elements(247) & zeropad3D_A_CP_1983_elements(251) & zeropad3D_A_CP_1983_elements(255);
      gj_zeropad3D_A_cp_element_group_178 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(178), clk => clk, reset => reset); --
    end block;
    -- CP-element group 179:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	177 
    -- CP-element group 179: successors 
    -- CP-element group 179: marked-successors 
    -- CP-element group 179: 	110 
    -- CP-element group 179: 	114 
    -- CP-element group 179: 	177 
    -- CP-element group 179:  members (3) 
      -- CP-element group 179: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1061_sample_completed_
      -- CP-element group 179: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1061_Sample/$exit
      -- CP-element group 179: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1061_Sample/ack
      -- 
    ack_2635_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xthen_ifx_xend80_taken_1022_delayed_3_0_1059_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(179)); -- 
    -- CP-element group 180:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	178 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	225 
    -- CP-element group 180: 	229 
    -- CP-element group 180: 	233 
    -- CP-element group 180: 	237 
    -- CP-element group 180: 	245 
    -- CP-element group 180: 	249 
    -- CP-element group 180: 	253 
    -- CP-element group 180: marked-successors 
    -- CP-element group 180: 	178 
    -- CP-element group 180:  members (3) 
      -- CP-element group 180: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1061_update_completed_
      -- CP-element group 180: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1061_Update/$exit
      -- CP-element group 180: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1061_Update/ack
      -- 
    ack_2640_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xthen_ifx_xend80_taken_1022_delayed_3_0_1059_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(180)); -- 
    -- CP-element group 181:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	112 
    -- CP-element group 181: 	116 
    -- CP-element group 181: marked-predecessors 
    -- CP-element group 181: 	183 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	183 
    -- CP-element group 181:  members (3) 
      -- CP-element group 181: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1071_sample_start_
      -- CP-element group 181: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1071_Sample/$entry
      -- CP-element group 181: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1071_Sample/req
      -- 
    req_2648_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2648_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(181), ack => W_ifx_xthen_ifx_xend80_taken_1028_delayed_3_0_1069_inst_req_0); -- 
    zeropad3D_A_cp_element_group_181: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_181"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(112) & zeropad3D_A_CP_1983_elements(116) & zeropad3D_A_CP_1983_elements(183);
      gj_zeropad3D_A_cp_element_group_181 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(181), clk => clk, reset => reset); --
    end block;
    -- CP-element group 182:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	45 
    -- CP-element group 182: marked-predecessors 
    -- CP-element group 182: 	184 
    -- CP-element group 182: 	299 
    -- CP-element group 182: 	330 
    -- CP-element group 182: 	365 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	184 
    -- CP-element group 182:  members (3) 
      -- CP-element group 182: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1071_update_start_
      -- CP-element group 182: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1071_Update/$entry
      -- CP-element group 182: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1071_Update/req
      -- 
    req_2653_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2653_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(182), ack => W_ifx_xthen_ifx_xend80_taken_1028_delayed_3_0_1069_inst_req_1); -- 
    zeropad3D_A_cp_element_group_182: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_182"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(45) & zeropad3D_A_CP_1983_elements(184) & zeropad3D_A_CP_1983_elements(299) & zeropad3D_A_CP_1983_elements(330) & zeropad3D_A_CP_1983_elements(365);
      gj_zeropad3D_A_cp_element_group_182 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(182), clk => clk, reset => reset); --
    end block;
    -- CP-element group 183:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	181 
    -- CP-element group 183: successors 
    -- CP-element group 183: marked-successors 
    -- CP-element group 183: 	110 
    -- CP-element group 183: 	114 
    -- CP-element group 183: 	181 
    -- CP-element group 183:  members (3) 
      -- CP-element group 183: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1071_sample_completed_
      -- CP-element group 183: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1071_Sample/$exit
      -- CP-element group 183: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1071_Sample/ack
      -- 
    ack_2649_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xthen_ifx_xend80_taken_1028_delayed_3_0_1069_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(183)); -- 
    -- CP-element group 184:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	182 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	297 
    -- CP-element group 184: 	328 
    -- CP-element group 184: 	363 
    -- CP-element group 184: marked-successors 
    -- CP-element group 184: 	48 
    -- CP-element group 184: 	182 
    -- CP-element group 184:  members (3) 
      -- CP-element group 184: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1071_update_completed_
      -- CP-element group 184: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1071_Update/$exit
      -- CP-element group 184: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1071_Update/ack
      -- 
    ack_2654_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xthen_ifx_xend80_taken_1028_delayed_3_0_1069_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(184)); -- 
    -- CP-element group 185:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	120 
    -- CP-element group 185: marked-predecessors 
    -- CP-element group 185: 	187 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	187 
    -- CP-element group 185:  members (3) 
      -- CP-element group 185: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1074_sample_start_
      -- CP-element group 185: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1074_Sample/$entry
      -- CP-element group 185: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1074_Sample/rr
      -- 
    rr_2662_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2662_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(185), ack => type_cast_1074_inst_req_0); -- 
    zeropad3D_A_cp_element_group_185: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_185"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(120) & zeropad3D_A_CP_1983_elements(187);
      gj_zeropad3D_A_cp_element_group_185 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(185), clk => clk, reset => reset); --
    end block;
    -- CP-element group 186:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	45 
    -- CP-element group 186: marked-predecessors 
    -- CP-element group 186: 	188 
    -- CP-element group 186: 	299 
    -- CP-element group 186: 	330 
    -- CP-element group 186: 	365 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	188 
    -- CP-element group 186:  members (3) 
      -- CP-element group 186: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1074_update_start_
      -- CP-element group 186: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1074_Update/$entry
      -- CP-element group 186: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1074_Update/cr
      -- 
    cr_2667_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2667_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(186), ack => type_cast_1074_inst_req_1); -- 
    zeropad3D_A_cp_element_group_186: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_186"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(45) & zeropad3D_A_CP_1983_elements(188) & zeropad3D_A_CP_1983_elements(299) & zeropad3D_A_CP_1983_elements(330) & zeropad3D_A_CP_1983_elements(365);
      gj_zeropad3D_A_cp_element_group_186 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(186), clk => clk, reset => reset); --
    end block;
    -- CP-element group 187:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	185 
    -- CP-element group 187: successors 
    -- CP-element group 187: marked-successors 
    -- CP-element group 187: 	118 
    -- CP-element group 187: 	185 
    -- CP-element group 187:  members (3) 
      -- CP-element group 187: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1074_sample_completed_
      -- CP-element group 187: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1074_Sample/$exit
      -- CP-element group 187: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1074_Sample/ra
      -- 
    ra_2663_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1074_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(187)); -- 
    -- CP-element group 188:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	186 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	297 
    -- CP-element group 188: 	328 
    -- CP-element group 188: 	363 
    -- CP-element group 188: marked-successors 
    -- CP-element group 188: 	48 
    -- CP-element group 188: 	186 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1074_update_completed_
      -- CP-element group 188: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1074_Update/$exit
      -- CP-element group 188: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1074_Update/ca
      -- 
    ca_2668_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1074_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(188)); -- 
    -- CP-element group 189:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	112 
    -- CP-element group 189: 	116 
    -- CP-element group 189: marked-predecessors 
    -- CP-element group 189: 	191 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	191 
    -- CP-element group 189:  members (3) 
      -- CP-element group 189: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1095_sample_start_
      -- CP-element group 189: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1095_Sample/$entry
      -- CP-element group 189: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1095_Sample/req
      -- 
    req_2676_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2676_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(189), ack => W_ifx_xthen_ifx_xend80_taken_1046_delayed_3_0_1093_inst_req_0); -- 
    zeropad3D_A_cp_element_group_189: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_189"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(112) & zeropad3D_A_CP_1983_elements(116) & zeropad3D_A_CP_1983_elements(191);
      gj_zeropad3D_A_cp_element_group_189 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(189), clk => clk, reset => reset); --
    end block;
    -- CP-element group 190:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	45 
    -- CP-element group 190: marked-predecessors 
    -- CP-element group 190: 	192 
    -- CP-element group 190: 	227 
    -- CP-element group 190: 	299 
    -- CP-element group 190: 	330 
    -- CP-element group 190: 	365 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	192 
    -- CP-element group 190:  members (3) 
      -- CP-element group 190: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1095_update_start_
      -- CP-element group 190: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1095_Update/$entry
      -- CP-element group 190: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1095_Update/req
      -- 
    req_2681_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2681_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(190), ack => W_ifx_xthen_ifx_xend80_taken_1046_delayed_3_0_1093_inst_req_1); -- 
    zeropad3D_A_cp_element_group_190: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_190"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(45) & zeropad3D_A_CP_1983_elements(192) & zeropad3D_A_CP_1983_elements(227) & zeropad3D_A_CP_1983_elements(299) & zeropad3D_A_CP_1983_elements(330) & zeropad3D_A_CP_1983_elements(365);
      gj_zeropad3D_A_cp_element_group_190 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(190), clk => clk, reset => reset); --
    end block;
    -- CP-element group 191:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	189 
    -- CP-element group 191: successors 
    -- CP-element group 191: marked-successors 
    -- CP-element group 191: 	110 
    -- CP-element group 191: 	114 
    -- CP-element group 191: 	189 
    -- CP-element group 191:  members (3) 
      -- CP-element group 191: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1095_sample_completed_
      -- CP-element group 191: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1095_Sample/$exit
      -- CP-element group 191: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1095_Sample/ack
      -- 
    ack_2677_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xthen_ifx_xend80_taken_1046_delayed_3_0_1093_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(191)); -- 
    -- CP-element group 192:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	190 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	225 
    -- CP-element group 192: 	297 
    -- CP-element group 192: 	328 
    -- CP-element group 192: 	363 
    -- CP-element group 192: marked-successors 
    -- CP-element group 192: 	67 
    -- CP-element group 192: 	190 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1095_update_completed_
      -- CP-element group 192: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1095_Update/$exit
      -- CP-element group 192: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1095_Update/ack
      -- 
    ack_2682_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xthen_ifx_xend80_taken_1046_delayed_3_0_1093_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(192)); -- 
    -- CP-element group 193:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	72 
    -- CP-element group 193: marked-predecessors 
    -- CP-element group 193: 	195 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	195 
    -- CP-element group 193:  members (3) 
      -- CP-element group 193: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1098_sample_start_
      -- CP-element group 193: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1098_Sample/$entry
      -- CP-element group 193: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1098_Sample/rr
      -- 
    rr_2690_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2690_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(193), ack => type_cast_1098_inst_req_0); -- 
    zeropad3D_A_cp_element_group_193: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_193"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(72) & zeropad3D_A_CP_1983_elements(195);
      gj_zeropad3D_A_cp_element_group_193 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(193), clk => clk, reset => reset); --
    end block;
    -- CP-element group 194:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	45 
    -- CP-element group 194: marked-predecessors 
    -- CP-element group 194: 	196 
    -- CP-element group 194: 	227 
    -- CP-element group 194: 	299 
    -- CP-element group 194: 	330 
    -- CP-element group 194: 	365 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	196 
    -- CP-element group 194:  members (3) 
      -- CP-element group 194: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1098_update_start_
      -- CP-element group 194: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1098_Update/$entry
      -- CP-element group 194: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1098_Update/cr
      -- 
    cr_2695_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2695_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(194), ack => type_cast_1098_inst_req_1); -- 
    zeropad3D_A_cp_element_group_194: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_194"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(45) & zeropad3D_A_CP_1983_elements(196) & zeropad3D_A_CP_1983_elements(227) & zeropad3D_A_CP_1983_elements(299) & zeropad3D_A_CP_1983_elements(330) & zeropad3D_A_CP_1983_elements(365);
      gj_zeropad3D_A_cp_element_group_194 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(194), clk => clk, reset => reset); --
    end block;
    -- CP-element group 195:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	193 
    -- CP-element group 195: successors 
    -- CP-element group 195: marked-successors 
    -- CP-element group 195: 	68 
    -- CP-element group 195: 	193 
    -- CP-element group 195:  members (3) 
      -- CP-element group 195: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1098_sample_completed_
      -- CP-element group 195: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1098_Sample/$exit
      -- CP-element group 195: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1098_Sample/ra
      -- 
    ra_2691_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1098_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(195)); -- 
    -- CP-element group 196:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	194 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	225 
    -- CP-element group 196: 	297 
    -- CP-element group 196: 	328 
    -- CP-element group 196: 	363 
    -- CP-element group 196: marked-successors 
    -- CP-element group 196: 	67 
    -- CP-element group 196: 	194 
    -- CP-element group 196:  members (3) 
      -- CP-element group 196: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1098_update_completed_
      -- CP-element group 196: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1098_Update/$exit
      -- CP-element group 196: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1098_Update/ca
      -- 
    ca_2696_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1098_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(196)); -- 
    -- CP-element group 197:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	140 
    -- CP-element group 197: 	148 
    -- CP-element group 197: marked-predecessors 
    -- CP-element group 197: 	199 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	199 
    -- CP-element group 197:  members (3) 
      -- CP-element group 197: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1102_sample_start_
      -- CP-element group 197: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1102_Sample/$entry
      -- CP-element group 197: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1102_Sample/rr
      -- 
    rr_2704_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2704_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(197), ack => type_cast_1102_inst_req_0); -- 
    zeropad3D_A_cp_element_group_197: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_197"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(140) & zeropad3D_A_CP_1983_elements(148) & zeropad3D_A_CP_1983_elements(199);
      gj_zeropad3D_A_cp_element_group_197 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(197), clk => clk, reset => reset); --
    end block;
    -- CP-element group 198:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	45 
    -- CP-element group 198: marked-predecessors 
    -- CP-element group 198: 	200 
    -- CP-element group 198: 	227 
    -- CP-element group 198: 	299 
    -- CP-element group 198: 	330 
    -- CP-element group 198: 	365 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	200 
    -- CP-element group 198:  members (3) 
      -- CP-element group 198: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1102_update_start_
      -- CP-element group 198: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1102_Update/$entry
      -- CP-element group 198: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1102_Update/cr
      -- 
    cr_2709_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2709_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(198), ack => type_cast_1102_inst_req_1); -- 
    zeropad3D_A_cp_element_group_198: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_198"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(45) & zeropad3D_A_CP_1983_elements(200) & zeropad3D_A_CP_1983_elements(227) & zeropad3D_A_CP_1983_elements(299) & zeropad3D_A_CP_1983_elements(330) & zeropad3D_A_CP_1983_elements(365);
      gj_zeropad3D_A_cp_element_group_198 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(198), clk => clk, reset => reset); --
    end block;
    -- CP-element group 199:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	197 
    -- CP-element group 199: successors 
    -- CP-element group 199: marked-successors 
    -- CP-element group 199: 	138 
    -- CP-element group 199: 	146 
    -- CP-element group 199: 	197 
    -- CP-element group 199:  members (3) 
      -- CP-element group 199: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1102_sample_completed_
      -- CP-element group 199: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1102_Sample/$exit
      -- CP-element group 199: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1102_Sample/ra
      -- 
    ra_2705_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1102_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(199)); -- 
    -- CP-element group 200:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	198 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	225 
    -- CP-element group 200: 	297 
    -- CP-element group 200: 	328 
    -- CP-element group 200: 	363 
    -- CP-element group 200: marked-successors 
    -- CP-element group 200: 	67 
    -- CP-element group 200: 	198 
    -- CP-element group 200:  members (3) 
      -- CP-element group 200: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1102_update_completed_
      -- CP-element group 200: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1102_Update/$exit
      -- CP-element group 200: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1102_Update/ca
      -- 
    ca_2710_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 200_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1102_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(200)); -- 
    -- CP-element group 201:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	140 
    -- CP-element group 201: 	148 
    -- CP-element group 201: marked-predecessors 
    -- CP-element group 201: 	203 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	203 
    -- CP-element group 201:  members (3) 
      -- CP-element group 201: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1106_sample_start_
      -- CP-element group 201: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1106_Sample/$entry
      -- CP-element group 201: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1106_Sample/rr
      -- 
    rr_2718_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2718_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(201), ack => type_cast_1106_inst_req_0); -- 
    zeropad3D_A_cp_element_group_201: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_201"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(140) & zeropad3D_A_CP_1983_elements(148) & zeropad3D_A_CP_1983_elements(203);
      gj_zeropad3D_A_cp_element_group_201 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(201), clk => clk, reset => reset); --
    end block;
    -- CP-element group 202:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	45 
    -- CP-element group 202: marked-predecessors 
    -- CP-element group 202: 	204 
    -- CP-element group 202: 	227 
    -- CP-element group 202: 	299 
    -- CP-element group 202: 	330 
    -- CP-element group 202: 	365 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	204 
    -- CP-element group 202:  members (3) 
      -- CP-element group 202: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1106_update_start_
      -- CP-element group 202: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1106_Update/$entry
      -- CP-element group 202: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1106_Update/cr
      -- 
    cr_2723_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2723_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(202), ack => type_cast_1106_inst_req_1); -- 
    zeropad3D_A_cp_element_group_202: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_202"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(45) & zeropad3D_A_CP_1983_elements(204) & zeropad3D_A_CP_1983_elements(227) & zeropad3D_A_CP_1983_elements(299) & zeropad3D_A_CP_1983_elements(330) & zeropad3D_A_CP_1983_elements(365);
      gj_zeropad3D_A_cp_element_group_202 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(202), clk => clk, reset => reset); --
    end block;
    -- CP-element group 203:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	201 
    -- CP-element group 203: successors 
    -- CP-element group 203: marked-successors 
    -- CP-element group 203: 	138 
    -- CP-element group 203: 	146 
    -- CP-element group 203: 	201 
    -- CP-element group 203:  members (3) 
      -- CP-element group 203: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1106_sample_completed_
      -- CP-element group 203: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1106_Sample/$exit
      -- CP-element group 203: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1106_Sample/ra
      -- 
    ra_2719_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 203_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1106_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(203)); -- 
    -- CP-element group 204:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	202 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	225 
    -- CP-element group 204: 	297 
    -- CP-element group 204: 	328 
    -- CP-element group 204: 	363 
    -- CP-element group 204: marked-successors 
    -- CP-element group 204: 	67 
    -- CP-element group 204: 	202 
    -- CP-element group 204:  members (3) 
      -- CP-element group 204: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1106_update_completed_
      -- CP-element group 204: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1106_Update/$exit
      -- CP-element group 204: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1106_Update/ca
      -- 
    ca_2724_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 204_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1106_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(204)); -- 
    -- CP-element group 205:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	112 
    -- CP-element group 205: 	116 
    -- CP-element group 205: marked-predecessors 
    -- CP-element group 205: 	207 
    -- CP-element group 205: successors 
    -- CP-element group 205: 	207 
    -- CP-element group 205:  members (3) 
      -- CP-element group 205: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1123_sample_start_
      -- CP-element group 205: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1123_Sample/$entry
      -- CP-element group 205: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1123_Sample/req
      -- 
    req_2732_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2732_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(205), ack => W_ifx_xthen_ifx_xend80_taken_1062_delayed_3_0_1121_inst_req_0); -- 
    zeropad3D_A_cp_element_group_205: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_205"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(112) & zeropad3D_A_CP_1983_elements(116) & zeropad3D_A_CP_1983_elements(207);
      gj_zeropad3D_A_cp_element_group_205 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(205), clk => clk, reset => reset); --
    end block;
    -- CP-element group 206:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	45 
    -- CP-element group 206: marked-predecessors 
    -- CP-element group 206: 	208 
    -- CP-element group 206: 	259 
    -- CP-element group 206: 	299 
    -- CP-element group 206: 	330 
    -- CP-element group 206: 	365 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	208 
    -- CP-element group 206:  members (3) 
      -- CP-element group 206: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1123_update_start_
      -- CP-element group 206: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1123_Update/$entry
      -- CP-element group 206: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1123_Update/req
      -- 
    req_2737_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2737_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(206), ack => W_ifx_xthen_ifx_xend80_taken_1062_delayed_3_0_1121_inst_req_1); -- 
    zeropad3D_A_cp_element_group_206: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_206"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(45) & zeropad3D_A_CP_1983_elements(208) & zeropad3D_A_CP_1983_elements(259) & zeropad3D_A_CP_1983_elements(299) & zeropad3D_A_CP_1983_elements(330) & zeropad3D_A_CP_1983_elements(365);
      gj_zeropad3D_A_cp_element_group_206 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(206), clk => clk, reset => reset); --
    end block;
    -- CP-element group 207:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	205 
    -- CP-element group 207: successors 
    -- CP-element group 207: marked-successors 
    -- CP-element group 207: 	110 
    -- CP-element group 207: 	114 
    -- CP-element group 207: 	205 
    -- CP-element group 207:  members (3) 
      -- CP-element group 207: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1123_sample_completed_
      -- CP-element group 207: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1123_Sample/$exit
      -- CP-element group 207: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1123_Sample/ack
      -- 
    ack_2733_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 207_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xthen_ifx_xend80_taken_1062_delayed_3_0_1121_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(207)); -- 
    -- CP-element group 208:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	206 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	257 
    -- CP-element group 208: 	297 
    -- CP-element group 208: 	328 
    -- CP-element group 208: 	363 
    -- CP-element group 208: marked-successors 
    -- CP-element group 208: 	88 
    -- CP-element group 208: 	206 
    -- CP-element group 208:  members (3) 
      -- CP-element group 208: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1123_update_completed_
      -- CP-element group 208: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1123_Update/$exit
      -- CP-element group 208: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1123_Update/ack
      -- 
    ack_2738_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 208_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xthen_ifx_xend80_taken_1062_delayed_3_0_1121_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(208)); -- 
    -- CP-element group 209:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	93 
    -- CP-element group 209: marked-predecessors 
    -- CP-element group 209: 	211 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	211 
    -- CP-element group 209:  members (3) 
      -- CP-element group 209: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1126_sample_start_
      -- CP-element group 209: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1126_Sample/$entry
      -- CP-element group 209: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1126_Sample/rr
      -- 
    rr_2746_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2746_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(209), ack => type_cast_1126_inst_req_0); -- 
    zeropad3D_A_cp_element_group_209: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_209"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(93) & zeropad3D_A_CP_1983_elements(211);
      gj_zeropad3D_A_cp_element_group_209 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(209), clk => clk, reset => reset); --
    end block;
    -- CP-element group 210:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	45 
    -- CP-element group 210: marked-predecessors 
    -- CP-element group 210: 	212 
    -- CP-element group 210: 	259 
    -- CP-element group 210: 	299 
    -- CP-element group 210: 	330 
    -- CP-element group 210: 	365 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	212 
    -- CP-element group 210:  members (3) 
      -- CP-element group 210: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1126_update_start_
      -- CP-element group 210: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1126_Update/$entry
      -- CP-element group 210: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1126_Update/cr
      -- 
    cr_2751_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2751_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(210), ack => type_cast_1126_inst_req_1); -- 
    zeropad3D_A_cp_element_group_210: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_210"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(45) & zeropad3D_A_CP_1983_elements(212) & zeropad3D_A_CP_1983_elements(259) & zeropad3D_A_CP_1983_elements(299) & zeropad3D_A_CP_1983_elements(330) & zeropad3D_A_CP_1983_elements(365);
      gj_zeropad3D_A_cp_element_group_210 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(210), clk => clk, reset => reset); --
    end block;
    -- CP-element group 211:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	209 
    -- CP-element group 211: successors 
    -- CP-element group 211: marked-successors 
    -- CP-element group 211: 	89 
    -- CP-element group 211: 	209 
    -- CP-element group 211:  members (3) 
      -- CP-element group 211: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1126_sample_completed_
      -- CP-element group 211: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1126_Sample/$exit
      -- CP-element group 211: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1126_Sample/ra
      -- 
    ra_2747_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 211_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1126_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(211)); -- 
    -- CP-element group 212:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	210 
    -- CP-element group 212: successors 
    -- CP-element group 212: 	257 
    -- CP-element group 212: 	297 
    -- CP-element group 212: 	328 
    -- CP-element group 212: 	363 
    -- CP-element group 212: marked-successors 
    -- CP-element group 212: 	88 
    -- CP-element group 212: 	210 
    -- CP-element group 212:  members (3) 
      -- CP-element group 212: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1126_update_completed_
      -- CP-element group 212: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1126_Update/$exit
      -- CP-element group 212: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1126_Update/ca
      -- 
    ca_2752_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 212_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1126_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(212)); -- 
    -- CP-element group 213:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	128 
    -- CP-element group 213: 	156 
    -- CP-element group 213: marked-predecessors 
    -- CP-element group 213: 	215 
    -- CP-element group 213: successors 
    -- CP-element group 213: 	215 
    -- CP-element group 213:  members (3) 
      -- CP-element group 213: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1130_sample_start_
      -- CP-element group 213: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1130_Sample/$entry
      -- CP-element group 213: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1130_Sample/rr
      -- 
    rr_2760_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2760_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(213), ack => type_cast_1130_inst_req_0); -- 
    zeropad3D_A_cp_element_group_213: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_213"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(128) & zeropad3D_A_CP_1983_elements(156) & zeropad3D_A_CP_1983_elements(215);
      gj_zeropad3D_A_cp_element_group_213 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(213), clk => clk, reset => reset); --
    end block;
    -- CP-element group 214:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	45 
    -- CP-element group 214: marked-predecessors 
    -- CP-element group 214: 	216 
    -- CP-element group 214: 	259 
    -- CP-element group 214: 	299 
    -- CP-element group 214: 	330 
    -- CP-element group 214: 	365 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	216 
    -- CP-element group 214:  members (3) 
      -- CP-element group 214: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1130_update_start_
      -- CP-element group 214: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1130_Update/$entry
      -- CP-element group 214: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1130_Update/cr
      -- 
    cr_2765_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2765_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(214), ack => type_cast_1130_inst_req_1); -- 
    zeropad3D_A_cp_element_group_214: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_214"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(45) & zeropad3D_A_CP_1983_elements(216) & zeropad3D_A_CP_1983_elements(259) & zeropad3D_A_CP_1983_elements(299) & zeropad3D_A_CP_1983_elements(330) & zeropad3D_A_CP_1983_elements(365);
      gj_zeropad3D_A_cp_element_group_214 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(214), clk => clk, reset => reset); --
    end block;
    -- CP-element group 215:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	213 
    -- CP-element group 215: successors 
    -- CP-element group 215: marked-successors 
    -- CP-element group 215: 	126 
    -- CP-element group 215: 	154 
    -- CP-element group 215: 	213 
    -- CP-element group 215:  members (3) 
      -- CP-element group 215: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1130_sample_completed_
      -- CP-element group 215: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1130_Sample/$exit
      -- CP-element group 215: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1130_Sample/ra
      -- 
    ra_2761_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 215_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1130_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(215)); -- 
    -- CP-element group 216:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	214 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	257 
    -- CP-element group 216: 	297 
    -- CP-element group 216: 	328 
    -- CP-element group 216: 	363 
    -- CP-element group 216: marked-successors 
    -- CP-element group 216: 	88 
    -- CP-element group 216: 	214 
    -- CP-element group 216:  members (3) 
      -- CP-element group 216: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1130_update_completed_
      -- CP-element group 216: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1130_Update/$exit
      -- CP-element group 216: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1130_Update/ca
      -- 
    ca_2766_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1130_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(216)); -- 
    -- CP-element group 217:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	128 
    -- CP-element group 217: 	156 
    -- CP-element group 217: marked-predecessors 
    -- CP-element group 217: 	219 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	219 
    -- CP-element group 217:  members (3) 
      -- CP-element group 217: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1134_sample_start_
      -- CP-element group 217: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1134_Sample/$entry
      -- CP-element group 217: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1134_Sample/rr
      -- 
    rr_2774_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2774_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(217), ack => type_cast_1134_inst_req_0); -- 
    zeropad3D_A_cp_element_group_217: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_217"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(128) & zeropad3D_A_CP_1983_elements(156) & zeropad3D_A_CP_1983_elements(219);
      gj_zeropad3D_A_cp_element_group_217 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(217), clk => clk, reset => reset); --
    end block;
    -- CP-element group 218:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	45 
    -- CP-element group 218: marked-predecessors 
    -- CP-element group 218: 	220 
    -- CP-element group 218: 	259 
    -- CP-element group 218: 	299 
    -- CP-element group 218: 	330 
    -- CP-element group 218: 	365 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	220 
    -- CP-element group 218:  members (3) 
      -- CP-element group 218: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1134_update_start_
      -- CP-element group 218: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1134_Update/$entry
      -- CP-element group 218: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1134_Update/cr
      -- 
    cr_2779_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2779_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(218), ack => type_cast_1134_inst_req_1); -- 
    zeropad3D_A_cp_element_group_218: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_218"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(45) & zeropad3D_A_CP_1983_elements(220) & zeropad3D_A_CP_1983_elements(259) & zeropad3D_A_CP_1983_elements(299) & zeropad3D_A_CP_1983_elements(330) & zeropad3D_A_CP_1983_elements(365);
      gj_zeropad3D_A_cp_element_group_218 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(218), clk => clk, reset => reset); --
    end block;
    -- CP-element group 219:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	217 
    -- CP-element group 219: successors 
    -- CP-element group 219: marked-successors 
    -- CP-element group 219: 	126 
    -- CP-element group 219: 	154 
    -- CP-element group 219: 	217 
    -- CP-element group 219:  members (3) 
      -- CP-element group 219: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1134_sample_completed_
      -- CP-element group 219: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1134_Sample/$exit
      -- CP-element group 219: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1134_Sample/ra
      -- 
    ra_2775_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 219_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1134_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(219)); -- 
    -- CP-element group 220:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	218 
    -- CP-element group 220: successors 
    -- CP-element group 220: 	257 
    -- CP-element group 220: 	297 
    -- CP-element group 220: 	328 
    -- CP-element group 220: 	363 
    -- CP-element group 220: marked-successors 
    -- CP-element group 220: 	88 
    -- CP-element group 220: 	218 
    -- CP-element group 220:  members (3) 
      -- CP-element group 220: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1134_update_completed_
      -- CP-element group 220: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1134_Update/$exit
      -- CP-element group 220: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1134_Update/ca
      -- 
    ca_2780_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1134_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(220)); -- 
    -- CP-element group 221:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	112 
    -- CP-element group 221: 	116 
    -- CP-element group 221: marked-predecessors 
    -- CP-element group 221: 	223 
    -- CP-element group 221: successors 
    -- CP-element group 221: 	223 
    -- CP-element group 221:  members (3) 
      -- CP-element group 221: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1151_Sample/req
      -- CP-element group 221: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1151_Sample/$entry
      -- CP-element group 221: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1151_sample_start_
      -- 
    req_2788_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2788_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(221), ack => W_ifx_xthen_ifx_xend80_taken_1078_delayed_3_0_1149_inst_req_0); -- 
    zeropad3D_A_cp_element_group_221: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_221"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(112) & zeropad3D_A_CP_1983_elements(116) & zeropad3D_A_CP_1983_elements(223);
      gj_zeropad3D_A_cp_element_group_221 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(221), clk => clk, reset => reset); --
    end block;
    -- CP-element group 222:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: marked-predecessors 
    -- CP-element group 222: 	224 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	224 
    -- CP-element group 222:  members (3) 
      -- CP-element group 222: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1151_Update/$entry
      -- CP-element group 222: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1151_Update/req
      -- CP-element group 222: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1151_update_start_
      -- 
    req_2793_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2793_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(222), ack => W_ifx_xthen_ifx_xend80_taken_1078_delayed_3_0_1149_inst_req_1); -- 
    zeropad3D_A_cp_element_group_222: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_222"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= zeropad3D_A_CP_1983_elements(224);
      gj_zeropad3D_A_cp_element_group_222 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(222), clk => clk, reset => reset); --
    end block;
    -- CP-element group 223:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	221 
    -- CP-element group 223: successors 
    -- CP-element group 223: marked-successors 
    -- CP-element group 223: 	110 
    -- CP-element group 223: 	114 
    -- CP-element group 223: 	221 
    -- CP-element group 223:  members (3) 
      -- CP-element group 223: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1151_Sample/ack
      -- CP-element group 223: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1151_Sample/$exit
      -- CP-element group 223: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1151_sample_completed_
      -- 
    ack_2789_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 223_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xthen_ifx_xend80_taken_1078_delayed_3_0_1149_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(223)); -- 
    -- CP-element group 224:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	222 
    -- CP-element group 224: successors 
    -- CP-element group 224: 	43 
    -- CP-element group 224: marked-successors 
    -- CP-element group 224: 	222 
    -- CP-element group 224:  members (3) 
      -- CP-element group 224: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1151_Update/$exit
      -- CP-element group 224: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1151_Update/ack
      -- CP-element group 224: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1151_update_completed_
      -- 
    ack_2794_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xthen_ifx_xend80_taken_1078_delayed_3_0_1149_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(224)); -- 
    -- CP-element group 225:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	164 
    -- CP-element group 225: 	172 
    -- CP-element group 225: 	176 
    -- CP-element group 225: 	180 
    -- CP-element group 225: 	192 
    -- CP-element group 225: 	196 
    -- CP-element group 225: 	200 
    -- CP-element group 225: 	204 
    -- CP-element group 225: marked-predecessors 
    -- CP-element group 225: 	227 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	227 
    -- CP-element group 225:  members (3) 
      -- CP-element group 225: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1234_Sample/rr
      -- CP-element group 225: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1234_sample_start_
      -- CP-element group 225: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1234_Sample/$entry
      -- 
    rr_2802_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2802_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(225), ack => type_cast_1234_inst_req_0); -- 
    zeropad3D_A_cp_element_group_225: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 1);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_225"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(164) & zeropad3D_A_CP_1983_elements(172) & zeropad3D_A_CP_1983_elements(176) & zeropad3D_A_CP_1983_elements(180) & zeropad3D_A_CP_1983_elements(192) & zeropad3D_A_CP_1983_elements(196) & zeropad3D_A_CP_1983_elements(200) & zeropad3D_A_CP_1983_elements(204) & zeropad3D_A_CP_1983_elements(227);
      gj_zeropad3D_A_cp_element_group_225 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(225), clk => clk, reset => reset); --
    end block;
    -- CP-element group 226:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: marked-predecessors 
    -- CP-element group 226: 	228 
    -- CP-element group 226: 	263 
    -- CP-element group 226: 	267 
    -- CP-element group 226: 	271 
    -- CP-element group 226: 	275 
    -- CP-element group 226: 	283 
    -- CP-element group 226: 	287 
    -- CP-element group 226: 	291 
    -- CP-element group 226: 	295 
    -- CP-element group 226: successors 
    -- CP-element group 226: 	228 
    -- CP-element group 226:  members (3) 
      -- CP-element group 226: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1234_Update/$entry
      -- CP-element group 226: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1234_Update/cr
      -- CP-element group 226: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1234_update_start_
      -- 
    cr_2807_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2807_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(226), ack => type_cast_1234_inst_req_1); -- 
    zeropad3D_A_cp_element_group_226: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_226"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(228) & zeropad3D_A_CP_1983_elements(263) & zeropad3D_A_CP_1983_elements(267) & zeropad3D_A_CP_1983_elements(271) & zeropad3D_A_CP_1983_elements(275) & zeropad3D_A_CP_1983_elements(283) & zeropad3D_A_CP_1983_elements(287) & zeropad3D_A_CP_1983_elements(291) & zeropad3D_A_CP_1983_elements(295);
      gj_zeropad3D_A_cp_element_group_226 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(226), clk => clk, reset => reset); --
    end block;
    -- CP-element group 227:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	225 
    -- CP-element group 227: successors 
    -- CP-element group 227: marked-successors 
    -- CP-element group 227: 	162 
    -- CP-element group 227: 	170 
    -- CP-element group 227: 	174 
    -- CP-element group 227: 	178 
    -- CP-element group 227: 	190 
    -- CP-element group 227: 	194 
    -- CP-element group 227: 	198 
    -- CP-element group 227: 	202 
    -- CP-element group 227: 	225 
    -- CP-element group 227:  members (3) 
      -- CP-element group 227: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1234_Sample/ra
      -- CP-element group 227: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1234_sample_completed_
      -- CP-element group 227: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1234_Sample/$exit
      -- 
    ra_2803_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 227_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1234_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(227)); -- 
    -- CP-element group 228:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	226 
    -- CP-element group 228: successors 
    -- CP-element group 228: 	261 
    -- CP-element group 228: 	265 
    -- CP-element group 228: 	269 
    -- CP-element group 228: 	273 
    -- CP-element group 228: 	281 
    -- CP-element group 228: 	285 
    -- CP-element group 228: 	289 
    -- CP-element group 228: 	293 
    -- CP-element group 228: marked-successors 
    -- CP-element group 228: 	226 
    -- CP-element group 228:  members (3) 
      -- CP-element group 228: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1234_Update/$exit
      -- CP-element group 228: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1234_Update/ca
      -- CP-element group 228: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1234_update_completed_
      -- 
    ca_2808_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 228_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1234_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(228)); -- 
    -- CP-element group 229:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	164 
    -- CP-element group 229: 	172 
    -- CP-element group 229: 	176 
    -- CP-element group 229: 	180 
    -- CP-element group 229: marked-predecessors 
    -- CP-element group 229: 	231 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	231 
    -- CP-element group 229:  members (3) 
      -- CP-element group 229: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1238_Sample/req
      -- CP-element group 229: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1238_Sample/$entry
      -- CP-element group 229: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1238_sample_start_
      -- 
    req_2816_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2816_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(229), ack => W_ifx_xend80_exec_guard_1161_delayed_1_0_1236_inst_req_0); -- 
    zeropad3D_A_cp_element_group_229: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_229"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(164) & zeropad3D_A_CP_1983_elements(172) & zeropad3D_A_CP_1983_elements(176) & zeropad3D_A_CP_1983_elements(180) & zeropad3D_A_CP_1983_elements(231);
      gj_zeropad3D_A_cp_element_group_229 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(229), clk => clk, reset => reset); --
    end block;
    -- CP-element group 230:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: marked-predecessors 
    -- CP-element group 230: 	232 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	232 
    -- CP-element group 230:  members (3) 
      -- CP-element group 230: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1238_Update/$entry
      -- CP-element group 230: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1238_Update/req
      -- CP-element group 230: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1238_update_start_
      -- 
    req_2821_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2821_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(230), ack => W_ifx_xend80_exec_guard_1161_delayed_1_0_1236_inst_req_1); -- 
    zeropad3D_A_cp_element_group_230: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_230"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= zeropad3D_A_CP_1983_elements(232);
      gj_zeropad3D_A_cp_element_group_230 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(230), clk => clk, reset => reset); --
    end block;
    -- CP-element group 231:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	229 
    -- CP-element group 231: successors 
    -- CP-element group 231: marked-successors 
    -- CP-element group 231: 	162 
    -- CP-element group 231: 	170 
    -- CP-element group 231: 	174 
    -- CP-element group 231: 	178 
    -- CP-element group 231: 	229 
    -- CP-element group 231:  members (3) 
      -- CP-element group 231: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1238_Sample/$exit
      -- CP-element group 231: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1238_Sample/ack
      -- CP-element group 231: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1238_sample_completed_
      -- 
    ack_2817_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 231_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xend80_exec_guard_1161_delayed_1_0_1236_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(231)); -- 
    -- CP-element group 232:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	230 
    -- CP-element group 232: successors 
    -- CP-element group 232: 	404 
    -- CP-element group 232: marked-successors 
    -- CP-element group 232: 	230 
    -- CP-element group 232:  members (3) 
      -- CP-element group 232: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1238_update_completed_
      -- CP-element group 232: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1238_Update/$exit
      -- CP-element group 232: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1238_Update/ack
      -- 
    ack_2822_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 232_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xend80_exec_guard_1161_delayed_1_0_1236_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(232)); -- 
    -- CP-element group 233:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	164 
    -- CP-element group 233: 	172 
    -- CP-element group 233: 	176 
    -- CP-element group 233: 	180 
    -- CP-element group 233: marked-predecessors 
    -- CP-element group 233: 	235 
    -- CP-element group 233: successors 
    -- CP-element group 233: 	235 
    -- CP-element group 233:  members (3) 
      -- CP-element group 233: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1247_Sample/req
      -- CP-element group 233: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1247_sample_start_
      -- CP-element group 233: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1247_Sample/$entry
      -- 
    req_2830_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2830_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(233), ack => W_ifx_xend80_exec_guard_1167_delayed_1_0_1245_inst_req_0); -- 
    zeropad3D_A_cp_element_group_233: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_233"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(164) & zeropad3D_A_CP_1983_elements(172) & zeropad3D_A_CP_1983_elements(176) & zeropad3D_A_CP_1983_elements(180) & zeropad3D_A_CP_1983_elements(235);
      gj_zeropad3D_A_cp_element_group_233 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(233), clk => clk, reset => reset); --
    end block;
    -- CP-element group 234:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: marked-predecessors 
    -- CP-element group 234: 	236 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	236 
    -- CP-element group 234:  members (3) 
      -- CP-element group 234: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1247_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1247_update_start_
      -- CP-element group 234: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1247_Update/req
      -- 
    req_2835_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2835_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(234), ack => W_ifx_xend80_exec_guard_1167_delayed_1_0_1245_inst_req_1); -- 
    zeropad3D_A_cp_element_group_234: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_234"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= zeropad3D_A_CP_1983_elements(236);
      gj_zeropad3D_A_cp_element_group_234 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(234), clk => clk, reset => reset); --
    end block;
    -- CP-element group 235:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	233 
    -- CP-element group 235: successors 
    -- CP-element group 235: marked-successors 
    -- CP-element group 235: 	162 
    -- CP-element group 235: 	170 
    -- CP-element group 235: 	174 
    -- CP-element group 235: 	178 
    -- CP-element group 235: 	233 
    -- CP-element group 235:  members (3) 
      -- CP-element group 235: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1247_Sample/ack
      -- CP-element group 235: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1247_sample_completed_
      -- CP-element group 235: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1247_Sample/$exit
      -- 
    ack_2831_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 235_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xend80_exec_guard_1167_delayed_1_0_1245_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(235)); -- 
    -- CP-element group 236:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	234 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	404 
    -- CP-element group 236: marked-successors 
    -- CP-element group 236: 	234 
    -- CP-element group 236:  members (3) 
      -- CP-element group 236: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1247_Update/$exit
      -- CP-element group 236: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1247_update_completed_
      -- CP-element group 236: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1247_Update/ack
      -- 
    ack_2836_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 236_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xend80_exec_guard_1167_delayed_1_0_1245_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(236)); -- 
    -- CP-element group 237:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	164 
    -- CP-element group 237: 	172 
    -- CP-element group 237: 	176 
    -- CP-element group 237: 	180 
    -- CP-element group 237: marked-predecessors 
    -- CP-element group 237: 	239 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	239 
    -- CP-element group 237:  members (3) 
      -- CP-element group 237: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1257_Sample/req
      -- CP-element group 237: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1257_Sample/$entry
      -- CP-element group 237: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1257_sample_start_
      -- 
    req_2844_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2844_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(237), ack => W_ifx_xend80_exec_guard_1174_delayed_1_0_1255_inst_req_0); -- 
    zeropad3D_A_cp_element_group_237: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_237"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(164) & zeropad3D_A_CP_1983_elements(172) & zeropad3D_A_CP_1983_elements(176) & zeropad3D_A_CP_1983_elements(180) & zeropad3D_A_CP_1983_elements(239);
      gj_zeropad3D_A_cp_element_group_237 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(237), clk => clk, reset => reset); --
    end block;
    -- CP-element group 238:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: marked-predecessors 
    -- CP-element group 238: 	240 
    -- CP-element group 238: successors 
    -- CP-element group 238: 	240 
    -- CP-element group 238:  members (3) 
      -- CP-element group 238: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1257_Update/req
      -- CP-element group 238: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1257_Update/$entry
      -- CP-element group 238: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1257_update_start_
      -- 
    req_2849_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2849_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(238), ack => W_ifx_xend80_exec_guard_1174_delayed_1_0_1255_inst_req_1); -- 
    zeropad3D_A_cp_element_group_238: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_238"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= zeropad3D_A_CP_1983_elements(240);
      gj_zeropad3D_A_cp_element_group_238 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(238), clk => clk, reset => reset); --
    end block;
    -- CP-element group 239:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	237 
    -- CP-element group 239: successors 
    -- CP-element group 239: marked-successors 
    -- CP-element group 239: 	162 
    -- CP-element group 239: 	170 
    -- CP-element group 239: 	174 
    -- CP-element group 239: 	178 
    -- CP-element group 239: 	237 
    -- CP-element group 239:  members (3) 
      -- CP-element group 239: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1257_Sample/ack
      -- CP-element group 239: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1257_Sample/$exit
      -- CP-element group 239: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1257_sample_completed_
      -- 
    ack_2845_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 239_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xend80_exec_guard_1174_delayed_1_0_1255_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(239)); -- 
    -- CP-element group 240:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	238 
    -- CP-element group 240: successors 
    -- CP-element group 240: 	404 
    -- CP-element group 240: marked-successors 
    -- CP-element group 240: 	238 
    -- CP-element group 240:  members (3) 
      -- CP-element group 240: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1257_Update/ack
      -- CP-element group 240: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1257_Update/$exit
      -- CP-element group 240: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1257_update_completed_
      -- 
    ack_2850_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 240_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xend80_exec_guard_1174_delayed_1_0_1255_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(240)); -- 
    -- CP-element group 241:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	42 
    -- CP-element group 241: marked-predecessors 
    -- CP-element group 241: 	243 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	243 
    -- CP-element group 241:  members (3) 
      -- CP-element group 241: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1260_Sample/rr
      -- CP-element group 241: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1260_Sample/$entry
      -- CP-element group 241: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1260_sample_start_
      -- 
    rr_2858_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2858_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(241), ack => type_cast_1260_inst_req_0); -- 
    zeropad3D_A_cp_element_group_241: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_241"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(42) & zeropad3D_A_CP_1983_elements(243);
      gj_zeropad3D_A_cp_element_group_241 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(241), clk => clk, reset => reset); --
    end block;
    -- CP-element group 242:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: marked-predecessors 
    -- CP-element group 242: 	244 
    -- CP-element group 242: 	263 
    -- CP-element group 242: 	267 
    -- CP-element group 242: 	271 
    -- CP-element group 242: 	275 
    -- CP-element group 242: 	283 
    -- CP-element group 242: 	287 
    -- CP-element group 242: 	291 
    -- CP-element group 242: 	295 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	244 
    -- CP-element group 242:  members (3) 
      -- CP-element group 242: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1260_Update/cr
      -- CP-element group 242: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1260_Update/$entry
      -- CP-element group 242: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1260_update_start_
      -- 
    cr_2863_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2863_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(242), ack => type_cast_1260_inst_req_1); -- 
    zeropad3D_A_cp_element_group_242: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_242"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(244) & zeropad3D_A_CP_1983_elements(263) & zeropad3D_A_CP_1983_elements(267) & zeropad3D_A_CP_1983_elements(271) & zeropad3D_A_CP_1983_elements(275) & zeropad3D_A_CP_1983_elements(283) & zeropad3D_A_CP_1983_elements(287) & zeropad3D_A_CP_1983_elements(291) & zeropad3D_A_CP_1983_elements(295);
      gj_zeropad3D_A_cp_element_group_242 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(242), clk => clk, reset => reset); --
    end block;
    -- CP-element group 243:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	241 
    -- CP-element group 243: successors 
    -- CP-element group 243: marked-successors 
    -- CP-element group 243: 	241 
    -- CP-element group 243:  members (3) 
      -- CP-element group 243: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1260_Sample/$exit
      -- CP-element group 243: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1260_Sample/ra
      -- CP-element group 243: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1260_sample_completed_
      -- 
    ra_2859_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 243_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1260_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(243)); -- 
    -- CP-element group 244:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	242 
    -- CP-element group 244: successors 
    -- CP-element group 244: 	261 
    -- CP-element group 244: 	265 
    -- CP-element group 244: 	269 
    -- CP-element group 244: 	273 
    -- CP-element group 244: 	281 
    -- CP-element group 244: 	285 
    -- CP-element group 244: 	289 
    -- CP-element group 244: 	293 
    -- CP-element group 244: marked-successors 
    -- CP-element group 244: 	242 
    -- CP-element group 244:  members (3) 
      -- CP-element group 244: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1260_Update/$exit
      -- CP-element group 244: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1260_Update/ca
      -- CP-element group 244: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1260_update_completed_
      -- 
    ca_2864_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 244_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1260_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(244)); -- 
    -- CP-element group 245:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	164 
    -- CP-element group 245: 	172 
    -- CP-element group 245: 	176 
    -- CP-element group 245: 	180 
    -- CP-element group 245: marked-predecessors 
    -- CP-element group 245: 	247 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	247 
    -- CP-element group 245:  members (3) 
      -- CP-element group 245: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1271_sample_start_
      -- CP-element group 245: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1271_Sample/$entry
      -- CP-element group 245: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1271_Sample/req
      -- 
    req_2872_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2872_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(245), ack => W_ifx_xend80_exec_guard_1182_delayed_1_0_1269_inst_req_0); -- 
    zeropad3D_A_cp_element_group_245: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_245"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(164) & zeropad3D_A_CP_1983_elements(172) & zeropad3D_A_CP_1983_elements(176) & zeropad3D_A_CP_1983_elements(180) & zeropad3D_A_CP_1983_elements(247);
      gj_zeropad3D_A_cp_element_group_245 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(245), clk => clk, reset => reset); --
    end block;
    -- CP-element group 246:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: marked-predecessors 
    -- CP-element group 246: 	248 
    -- CP-element group 246: successors 
    -- CP-element group 246: 	248 
    -- CP-element group 246:  members (3) 
      -- CP-element group 246: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1271_update_start_
      -- CP-element group 246: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1271_Update/$entry
      -- CP-element group 246: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1271_Update/req
      -- 
    req_2877_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2877_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(246), ack => W_ifx_xend80_exec_guard_1182_delayed_1_0_1269_inst_req_1); -- 
    zeropad3D_A_cp_element_group_246: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_246"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= zeropad3D_A_CP_1983_elements(248);
      gj_zeropad3D_A_cp_element_group_246 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(246), clk => clk, reset => reset); --
    end block;
    -- CP-element group 247:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	245 
    -- CP-element group 247: successors 
    -- CP-element group 247: marked-successors 
    -- CP-element group 247: 	162 
    -- CP-element group 247: 	170 
    -- CP-element group 247: 	174 
    -- CP-element group 247: 	178 
    -- CP-element group 247: 	245 
    -- CP-element group 247:  members (3) 
      -- CP-element group 247: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1271_sample_completed_
      -- CP-element group 247: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1271_Sample/$exit
      -- CP-element group 247: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1271_Sample/ack
      -- 
    ack_2873_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 247_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xend80_exec_guard_1182_delayed_1_0_1269_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(247)); -- 
    -- CP-element group 248:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	246 
    -- CP-element group 248: successors 
    -- CP-element group 248: 	404 
    -- CP-element group 248: marked-successors 
    -- CP-element group 248: 	246 
    -- CP-element group 248:  members (3) 
      -- CP-element group 248: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1271_update_completed_
      -- CP-element group 248: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1271_Update/$exit
      -- CP-element group 248: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1271_Update/ack
      -- 
    ack_2878_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 248_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xend80_exec_guard_1182_delayed_1_0_1269_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(248)); -- 
    -- CP-element group 249:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	164 
    -- CP-element group 249: 	172 
    -- CP-element group 249: 	176 
    -- CP-element group 249: 	180 
    -- CP-element group 249: marked-predecessors 
    -- CP-element group 249: 	251 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	251 
    -- CP-element group 249:  members (3) 
      -- CP-element group 249: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1280_Sample/req
      -- CP-element group 249: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1280_Sample/$entry
      -- CP-element group 249: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1280_sample_start_
      -- 
    req_2886_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2886_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(249), ack => W_ifx_xend80_exec_guard_1189_delayed_1_0_1278_inst_req_0); -- 
    zeropad3D_A_cp_element_group_249: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_249"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(164) & zeropad3D_A_CP_1983_elements(172) & zeropad3D_A_CP_1983_elements(176) & zeropad3D_A_CP_1983_elements(180) & zeropad3D_A_CP_1983_elements(251);
      gj_zeropad3D_A_cp_element_group_249 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(249), clk => clk, reset => reset); --
    end block;
    -- CP-element group 250:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: marked-predecessors 
    -- CP-element group 250: 	252 
    -- CP-element group 250: 	263 
    -- CP-element group 250: 	267 
    -- CP-element group 250: 	271 
    -- CP-element group 250: 	275 
    -- CP-element group 250: 	283 
    -- CP-element group 250: 	287 
    -- CP-element group 250: 	291 
    -- CP-element group 250: successors 
    -- CP-element group 250: 	252 
    -- CP-element group 250:  members (3) 
      -- CP-element group 250: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1280_Update/$entry
      -- CP-element group 250: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1280_Update/req
      -- CP-element group 250: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1280_update_start_
      -- 
    req_2891_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2891_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(250), ack => W_ifx_xend80_exec_guard_1189_delayed_1_0_1278_inst_req_1); -- 
    zeropad3D_A_cp_element_group_250: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_250"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(252) & zeropad3D_A_CP_1983_elements(263) & zeropad3D_A_CP_1983_elements(267) & zeropad3D_A_CP_1983_elements(271) & zeropad3D_A_CP_1983_elements(275) & zeropad3D_A_CP_1983_elements(283) & zeropad3D_A_CP_1983_elements(287) & zeropad3D_A_CP_1983_elements(291);
      gj_zeropad3D_A_cp_element_group_250 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(250), clk => clk, reset => reset); --
    end block;
    -- CP-element group 251:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	249 
    -- CP-element group 251: successors 
    -- CP-element group 251: marked-successors 
    -- CP-element group 251: 	162 
    -- CP-element group 251: 	170 
    -- CP-element group 251: 	174 
    -- CP-element group 251: 	178 
    -- CP-element group 251: 	249 
    -- CP-element group 251:  members (3) 
      -- CP-element group 251: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1280_Sample/ack
      -- CP-element group 251: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1280_Sample/$exit
      -- CP-element group 251: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1280_sample_completed_
      -- 
    ack_2887_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 251_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xend80_exec_guard_1189_delayed_1_0_1278_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(251)); -- 
    -- CP-element group 252:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	250 
    -- CP-element group 252: successors 
    -- CP-element group 252: 	261 
    -- CP-element group 252: 	265 
    -- CP-element group 252: 	269 
    -- CP-element group 252: 	273 
    -- CP-element group 252: 	281 
    -- CP-element group 252: 	285 
    -- CP-element group 252: 	289 
    -- CP-element group 252: marked-successors 
    -- CP-element group 252: 	250 
    -- CP-element group 252:  members (3) 
      -- CP-element group 252: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1280_update_completed_
      -- CP-element group 252: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1280_Update/$exit
      -- CP-element group 252: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1280_Update/ack
      -- 
    ack_2892_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 252_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xend80_exec_guard_1189_delayed_1_0_1278_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(252)); -- 
    -- CP-element group 253:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	164 
    -- CP-element group 253: 	172 
    -- CP-element group 253: 	176 
    -- CP-element group 253: 	180 
    -- CP-element group 253: marked-predecessors 
    -- CP-element group 253: 	255 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	255 
    -- CP-element group 253:  members (3) 
      -- CP-element group 253: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1288_Sample/req
      -- CP-element group 253: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1288_Sample/$entry
      -- CP-element group 253: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1288_sample_start_
      -- 
    req_2900_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2900_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(253), ack => W_ifx_xend80_exec_guard_1194_delayed_1_0_1286_inst_req_0); -- 
    zeropad3D_A_cp_element_group_253: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_253"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(164) & zeropad3D_A_CP_1983_elements(172) & zeropad3D_A_CP_1983_elements(176) & zeropad3D_A_CP_1983_elements(180) & zeropad3D_A_CP_1983_elements(255);
      gj_zeropad3D_A_cp_element_group_253 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(253), clk => clk, reset => reset); --
    end block;
    -- CP-element group 254:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: marked-predecessors 
    -- CP-element group 254: 	256 
    -- CP-element group 254: 	295 
    -- CP-element group 254: successors 
    -- CP-element group 254: 	256 
    -- CP-element group 254:  members (3) 
      -- CP-element group 254: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1288_Update/req
      -- CP-element group 254: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1288_Update/$entry
      -- CP-element group 254: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1288_update_start_
      -- 
    req_2905_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2905_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(254), ack => W_ifx_xend80_exec_guard_1194_delayed_1_0_1286_inst_req_1); -- 
    zeropad3D_A_cp_element_group_254: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_254"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(256) & zeropad3D_A_CP_1983_elements(295);
      gj_zeropad3D_A_cp_element_group_254 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(254), clk => clk, reset => reset); --
    end block;
    -- CP-element group 255:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	253 
    -- CP-element group 255: successors 
    -- CP-element group 255: marked-successors 
    -- CP-element group 255: 	162 
    -- CP-element group 255: 	170 
    -- CP-element group 255: 	174 
    -- CP-element group 255: 	178 
    -- CP-element group 255: 	253 
    -- CP-element group 255:  members (3) 
      -- CP-element group 255: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1288_Sample/ack
      -- CP-element group 255: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1288_Sample/$exit
      -- CP-element group 255: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1288_sample_completed_
      -- 
    ack_2901_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 255_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xend80_exec_guard_1194_delayed_1_0_1286_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(255)); -- 
    -- CP-element group 256:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	254 
    -- CP-element group 256: successors 
    -- CP-element group 256: 	293 
    -- CP-element group 256: marked-successors 
    -- CP-element group 256: 	254 
    -- CP-element group 256:  members (3) 
      -- CP-element group 256: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1288_Update/ack
      -- CP-element group 256: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1288_Update/$exit
      -- CP-element group 256: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1288_update_completed_
      -- 
    ack_2906_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 256_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xend80_exec_guard_1194_delayed_1_0_1286_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(256)); -- 
    -- CP-element group 257:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	164 
    -- CP-element group 257: 	172 
    -- CP-element group 257: 	176 
    -- CP-element group 257: 	208 
    -- CP-element group 257: 	212 
    -- CP-element group 257: 	216 
    -- CP-element group 257: 	220 
    -- CP-element group 257: marked-predecessors 
    -- CP-element group 257: 	259 
    -- CP-element group 257: successors 
    -- CP-element group 257: 	259 
    -- CP-element group 257:  members (3) 
      -- CP-element group 257: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1300_Sample/req
      -- CP-element group 257: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1300_Sample/$entry
      -- CP-element group 257: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1300_sample_start_
      -- 
    req_2914_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2914_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(257), ack => W_jx_x0_1204_delayed_1_0_1298_inst_req_0); -- 
    zeropad3D_A_cp_element_group_257: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_257"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(164) & zeropad3D_A_CP_1983_elements(172) & zeropad3D_A_CP_1983_elements(176) & zeropad3D_A_CP_1983_elements(208) & zeropad3D_A_CP_1983_elements(212) & zeropad3D_A_CP_1983_elements(216) & zeropad3D_A_CP_1983_elements(220) & zeropad3D_A_CP_1983_elements(259);
      gj_zeropad3D_A_cp_element_group_257 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(257), clk => clk, reset => reset); --
    end block;
    -- CP-element group 258:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: marked-predecessors 
    -- CP-element group 258: 	260 
    -- CP-element group 258: 	263 
    -- CP-element group 258: successors 
    -- CP-element group 258: 	260 
    -- CP-element group 258:  members (3) 
      -- CP-element group 258: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1300_Update/req
      -- CP-element group 258: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1300_Update/$entry
      -- CP-element group 258: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1300_update_start_
      -- 
    req_2919_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2919_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(258), ack => W_jx_x0_1204_delayed_1_0_1298_inst_req_1); -- 
    zeropad3D_A_cp_element_group_258: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_258"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(260) & zeropad3D_A_CP_1983_elements(263);
      gj_zeropad3D_A_cp_element_group_258 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(258), clk => clk, reset => reset); --
    end block;
    -- CP-element group 259:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	257 
    -- CP-element group 259: successors 
    -- CP-element group 259: marked-successors 
    -- CP-element group 259: 	162 
    -- CP-element group 259: 	170 
    -- CP-element group 259: 	174 
    -- CP-element group 259: 	206 
    -- CP-element group 259: 	210 
    -- CP-element group 259: 	214 
    -- CP-element group 259: 	218 
    -- CP-element group 259: 	257 
    -- CP-element group 259:  members (3) 
      -- CP-element group 259: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1300_Sample/ack
      -- CP-element group 259: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1300_Sample/$exit
      -- CP-element group 259: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1300_sample_completed_
      -- 
    ack_2915_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 259_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_jx_x0_1204_delayed_1_0_1298_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(259)); -- 
    -- CP-element group 260:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	258 
    -- CP-element group 260: successors 
    -- CP-element group 260: 	261 
    -- CP-element group 260: marked-successors 
    -- CP-element group 260: 	258 
    -- CP-element group 260:  members (3) 
      -- CP-element group 260: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1300_Update/ack
      -- CP-element group 260: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1300_Update/$exit
      -- CP-element group 260: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1300_update_completed_
      -- 
    ack_2920_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 260_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_jx_x0_1204_delayed_1_0_1298_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(260)); -- 
    -- CP-element group 261:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	228 
    -- CP-element group 261: 	244 
    -- CP-element group 261: 	252 
    -- CP-element group 261: 	260 
    -- CP-element group 261: marked-predecessors 
    -- CP-element group 261: 	263 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	263 
    -- CP-element group 261:  members (3) 
      -- CP-element group 261: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1304_Sample/rr
      -- CP-element group 261: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1304_Sample/$entry
      -- CP-element group 261: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1304_sample_start_
      -- 
    rr_2928_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2928_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(261), ack => type_cast_1304_inst_req_0); -- 
    zeropad3D_A_cp_element_group_261: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_261"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(228) & zeropad3D_A_CP_1983_elements(244) & zeropad3D_A_CP_1983_elements(252) & zeropad3D_A_CP_1983_elements(260) & zeropad3D_A_CP_1983_elements(263);
      gj_zeropad3D_A_cp_element_group_261 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(261), clk => clk, reset => reset); --
    end block;
    -- CP-element group 262:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: marked-predecessors 
    -- CP-element group 262: 	392 
    -- CP-element group 262: 	264 
    -- CP-element group 262: 	303 
    -- CP-element group 262: 	307 
    -- CP-element group 262: 	311 
    -- CP-element group 262: 	334 
    -- CP-element group 262: 	338 
    -- CP-element group 262: 	342 
    -- CP-element group 262: 	357 
    -- CP-element group 262: 	369 
    -- CP-element group 262: 	373 
    -- CP-element group 262: 	377 
    -- CP-element group 262: successors 
    -- CP-element group 262: 	264 
    -- CP-element group 262:  members (3) 
      -- CP-element group 262: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1304_Update/$entry
      -- CP-element group 262: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1304_Update/cr
      -- CP-element group 262: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1304_update_start_
      -- 
    cr_2933_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2933_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(262), ack => type_cast_1304_inst_req_1); -- 
    zeropad3D_A_cp_element_group_262: block -- 
      constant place_capacities: IntegerArray(0 to 11) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1);
      constant place_markings: IntegerArray(0 to 11)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1);
      constant place_delays: IntegerArray(0 to 11) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_262"; 
      signal preds: BooleanArray(1 to 12); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(392) & zeropad3D_A_CP_1983_elements(264) & zeropad3D_A_CP_1983_elements(303) & zeropad3D_A_CP_1983_elements(307) & zeropad3D_A_CP_1983_elements(311) & zeropad3D_A_CP_1983_elements(334) & zeropad3D_A_CP_1983_elements(338) & zeropad3D_A_CP_1983_elements(342) & zeropad3D_A_CP_1983_elements(357) & zeropad3D_A_CP_1983_elements(369) & zeropad3D_A_CP_1983_elements(373) & zeropad3D_A_CP_1983_elements(377);
      gj_zeropad3D_A_cp_element_group_262 : generic_join generic map(name => joinName, number_of_predecessors => 12, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(262), clk => clk, reset => reset); --
    end block;
    -- CP-element group 263:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	261 
    -- CP-element group 263: successors 
    -- CP-element group 263: marked-successors 
    -- CP-element group 263: 	226 
    -- CP-element group 263: 	242 
    -- CP-element group 263: 	250 
    -- CP-element group 263: 	258 
    -- CP-element group 263: 	261 
    -- CP-element group 263:  members (3) 
      -- CP-element group 263: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1304_Sample/ra
      -- CP-element group 263: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1304_Sample/$exit
      -- CP-element group 263: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1304_sample_completed_
      -- 
    ra_2929_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 263_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1304_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(263)); -- 
    -- CP-element group 264:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	262 
    -- CP-element group 264: successors 
    -- CP-element group 264: 	390 
    -- CP-element group 264: 	301 
    -- CP-element group 264: 	305 
    -- CP-element group 264: 	309 
    -- CP-element group 264: 	332 
    -- CP-element group 264: 	336 
    -- CP-element group 264: 	340 
    -- CP-element group 264: 	355 
    -- CP-element group 264: 	367 
    -- CP-element group 264: 	371 
    -- CP-element group 264: 	375 
    -- CP-element group 264: marked-successors 
    -- CP-element group 264: 	262 
    -- CP-element group 264:  members (3) 
      -- CP-element group 264: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1304_Update/$exit
      -- CP-element group 264: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1304_Update/ca
      -- CP-element group 264: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1304_update_completed_
      -- 
    ca_2934_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 264_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1304_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(264)); -- 
    -- CP-element group 265:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	228 
    -- CP-element group 265: 	244 
    -- CP-element group 265: 	252 
    -- CP-element group 265: marked-predecessors 
    -- CP-element group 265: 	267 
    -- CP-element group 265: successors 
    -- CP-element group 265: 	267 
    -- CP-element group 265:  members (3) 
      -- CP-element group 265: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1308_Sample/req
      -- CP-element group 265: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1308_Sample/$entry
      -- CP-element group 265: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1308_sample_start_
      -- 
    req_2942_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2942_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(265), ack => W_lorx_xlhsx_xfalse135_exec_guard_1207_delayed_1_0_1306_inst_req_0); -- 
    zeropad3D_A_cp_element_group_265: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_265"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(228) & zeropad3D_A_CP_1983_elements(244) & zeropad3D_A_CP_1983_elements(252) & zeropad3D_A_CP_1983_elements(267);
      gj_zeropad3D_A_cp_element_group_265 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(265), clk => clk, reset => reset); --
    end block;
    -- CP-element group 266:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: marked-predecessors 
    -- CP-element group 266: 	268 
    -- CP-element group 266: successors 
    -- CP-element group 266: 	268 
    -- CP-element group 266:  members (3) 
      -- CP-element group 266: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1308_Update/req
      -- CP-element group 266: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1308_Update/$entry
      -- CP-element group 266: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1308_update_start_
      -- 
    req_2947_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2947_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(266), ack => W_lorx_xlhsx_xfalse135_exec_guard_1207_delayed_1_0_1306_inst_req_1); -- 
    zeropad3D_A_cp_element_group_266: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_266"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= zeropad3D_A_CP_1983_elements(268);
      gj_zeropad3D_A_cp_element_group_266 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(266), clk => clk, reset => reset); --
    end block;
    -- CP-element group 267:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	265 
    -- CP-element group 267: successors 
    -- CP-element group 267: marked-successors 
    -- CP-element group 267: 	226 
    -- CP-element group 267: 	242 
    -- CP-element group 267: 	250 
    -- CP-element group 267: 	265 
    -- CP-element group 267:  members (3) 
      -- CP-element group 267: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1308_Sample/ack
      -- CP-element group 267: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1308_Sample/$exit
      -- CP-element group 267: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1308_sample_completed_
      -- 
    ack_2943_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 267_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_lorx_xlhsx_xfalse135_exec_guard_1207_delayed_1_0_1306_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(267)); -- 
    -- CP-element group 268:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	266 
    -- CP-element group 268: successors 
    -- CP-element group 268: 	404 
    -- CP-element group 268: marked-successors 
    -- CP-element group 268: 	266 
    -- CP-element group 268:  members (3) 
      -- CP-element group 268: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1308_Update/ack
      -- CP-element group 268: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1308_Update/$exit
      -- CP-element group 268: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1308_update_completed_
      -- 
    ack_2948_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 268_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_lorx_xlhsx_xfalse135_exec_guard_1207_delayed_1_0_1306_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(268)); -- 
    -- CP-element group 269:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: 	228 
    -- CP-element group 269: 	244 
    -- CP-element group 269: 	252 
    -- CP-element group 269: marked-predecessors 
    -- CP-element group 269: 	271 
    -- CP-element group 269: successors 
    -- CP-element group 269: 	271 
    -- CP-element group 269:  members (3) 
      -- CP-element group 269: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1317_Sample/req
      -- CP-element group 269: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1317_Sample/$entry
      -- CP-element group 269: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1317_sample_start_
      -- 
    req_2956_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2956_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(269), ack => W_lorx_xlhsx_xfalse135_exec_guard_1213_delayed_1_0_1315_inst_req_0); -- 
    zeropad3D_A_cp_element_group_269: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_269"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(228) & zeropad3D_A_CP_1983_elements(244) & zeropad3D_A_CP_1983_elements(252) & zeropad3D_A_CP_1983_elements(271);
      gj_zeropad3D_A_cp_element_group_269 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(269), clk => clk, reset => reset); --
    end block;
    -- CP-element group 270:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: marked-predecessors 
    -- CP-element group 270: 	272 
    -- CP-element group 270: successors 
    -- CP-element group 270: 	272 
    -- CP-element group 270:  members (3) 
      -- CP-element group 270: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1317_Update/req
      -- CP-element group 270: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1317_Update/$entry
      -- CP-element group 270: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1317_update_start_
      -- 
    req_2961_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2961_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(270), ack => W_lorx_xlhsx_xfalse135_exec_guard_1213_delayed_1_0_1315_inst_req_1); -- 
    zeropad3D_A_cp_element_group_270: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_270"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= zeropad3D_A_CP_1983_elements(272);
      gj_zeropad3D_A_cp_element_group_270 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(270), clk => clk, reset => reset); --
    end block;
    -- CP-element group 271:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	269 
    -- CP-element group 271: successors 
    -- CP-element group 271: marked-successors 
    -- CP-element group 271: 	226 
    -- CP-element group 271: 	242 
    -- CP-element group 271: 	250 
    -- CP-element group 271: 	269 
    -- CP-element group 271:  members (3) 
      -- CP-element group 271: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1317_Sample/ack
      -- CP-element group 271: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1317_Sample/$exit
      -- CP-element group 271: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1317_sample_completed_
      -- 
    ack_2957_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 271_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_lorx_xlhsx_xfalse135_exec_guard_1213_delayed_1_0_1315_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(271)); -- 
    -- CP-element group 272:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	270 
    -- CP-element group 272: successors 
    -- CP-element group 272: 	404 
    -- CP-element group 272: marked-successors 
    -- CP-element group 272: 	270 
    -- CP-element group 272:  members (3) 
      -- CP-element group 272: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1317_Update/ack
      -- CP-element group 272: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1317_Update/$exit
      -- CP-element group 272: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1317_update_completed_
      -- 
    ack_2962_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 272_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_lorx_xlhsx_xfalse135_exec_guard_1213_delayed_1_0_1315_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(272)); -- 
    -- CP-element group 273:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: 	228 
    -- CP-element group 273: 	244 
    -- CP-element group 273: 	252 
    -- CP-element group 273: marked-predecessors 
    -- CP-element group 273: 	275 
    -- CP-element group 273: successors 
    -- CP-element group 273: 	275 
    -- CP-element group 273:  members (3) 
      -- CP-element group 273: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1327_Sample/req
      -- CP-element group 273: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1327_Sample/$entry
      -- CP-element group 273: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1327_sample_start_
      -- 
    req_2970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(273), ack => W_lorx_xlhsx_xfalse135_exec_guard_1220_delayed_1_0_1325_inst_req_0); -- 
    zeropad3D_A_cp_element_group_273: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_273"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(228) & zeropad3D_A_CP_1983_elements(244) & zeropad3D_A_CP_1983_elements(252) & zeropad3D_A_CP_1983_elements(275);
      gj_zeropad3D_A_cp_element_group_273 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(273), clk => clk, reset => reset); --
    end block;
    -- CP-element group 274:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: marked-predecessors 
    -- CP-element group 274: 	276 
    -- CP-element group 274: successors 
    -- CP-element group 274: 	276 
    -- CP-element group 274:  members (3) 
      -- CP-element group 274: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1327_Update/req
      -- CP-element group 274: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1327_Update/$entry
      -- CP-element group 274: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1327_update_start_
      -- 
    req_2975_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2975_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(274), ack => W_lorx_xlhsx_xfalse135_exec_guard_1220_delayed_1_0_1325_inst_req_1); -- 
    zeropad3D_A_cp_element_group_274: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_274"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= zeropad3D_A_CP_1983_elements(276);
      gj_zeropad3D_A_cp_element_group_274 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(274), clk => clk, reset => reset); --
    end block;
    -- CP-element group 275:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	273 
    -- CP-element group 275: successors 
    -- CP-element group 275: marked-successors 
    -- CP-element group 275: 	226 
    -- CP-element group 275: 	242 
    -- CP-element group 275: 	250 
    -- CP-element group 275: 	273 
    -- CP-element group 275:  members (3) 
      -- CP-element group 275: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1327_Sample/ack
      -- CP-element group 275: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1327_Sample/$exit
      -- CP-element group 275: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1327_sample_completed_
      -- 
    ack_2971_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 275_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_lorx_xlhsx_xfalse135_exec_guard_1220_delayed_1_0_1325_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(275)); -- 
    -- CP-element group 276:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	274 
    -- CP-element group 276: successors 
    -- CP-element group 276: 	404 
    -- CP-element group 276: marked-successors 
    -- CP-element group 276: 	274 
    -- CP-element group 276:  members (3) 
      -- CP-element group 276: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1327_Update/ack
      -- CP-element group 276: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1327_Update/$exit
      -- CP-element group 276: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1327_update_completed_
      -- 
    ack_2976_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 276_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_lorx_xlhsx_xfalse135_exec_guard_1220_delayed_1_0_1325_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(276)); -- 
    -- CP-element group 277:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	42 
    -- CP-element group 277: marked-predecessors 
    -- CP-element group 277: 	279 
    -- CP-element group 277: successors 
    -- CP-element group 277: 	279 
    -- CP-element group 277:  members (3) 
      -- CP-element group 277: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1330_Sample/rr
      -- CP-element group 277: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1330_Sample/$entry
      -- CP-element group 277: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1330_sample_start_
      -- 
    rr_2984_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2984_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(277), ack => type_cast_1330_inst_req_0); -- 
    zeropad3D_A_cp_element_group_277: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_277"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(42) & zeropad3D_A_CP_1983_elements(279);
      gj_zeropad3D_A_cp_element_group_277 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(277), clk => clk, reset => reset); --
    end block;
    -- CP-element group 278:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: marked-predecessors 
    -- CP-element group 278: 	392 
    -- CP-element group 278: 	280 
    -- CP-element group 278: 	303 
    -- CP-element group 278: 	307 
    -- CP-element group 278: 	311 
    -- CP-element group 278: 	334 
    -- CP-element group 278: 	338 
    -- CP-element group 278: 	342 
    -- CP-element group 278: 	357 
    -- CP-element group 278: 	369 
    -- CP-element group 278: 	373 
    -- CP-element group 278: 	377 
    -- CP-element group 278: successors 
    -- CP-element group 278: 	280 
    -- CP-element group 278:  members (3) 
      -- CP-element group 278: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1330_Update/$entry
      -- CP-element group 278: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1330_Update/cr
      -- CP-element group 278: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1330_update_start_
      -- 
    cr_2989_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2989_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(278), ack => type_cast_1330_inst_req_1); -- 
    zeropad3D_A_cp_element_group_278: block -- 
      constant place_capacities: IntegerArray(0 to 11) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1);
      constant place_markings: IntegerArray(0 to 11)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1);
      constant place_delays: IntegerArray(0 to 11) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_278"; 
      signal preds: BooleanArray(1 to 12); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(392) & zeropad3D_A_CP_1983_elements(280) & zeropad3D_A_CP_1983_elements(303) & zeropad3D_A_CP_1983_elements(307) & zeropad3D_A_CP_1983_elements(311) & zeropad3D_A_CP_1983_elements(334) & zeropad3D_A_CP_1983_elements(338) & zeropad3D_A_CP_1983_elements(342) & zeropad3D_A_CP_1983_elements(357) & zeropad3D_A_CP_1983_elements(369) & zeropad3D_A_CP_1983_elements(373) & zeropad3D_A_CP_1983_elements(377);
      gj_zeropad3D_A_cp_element_group_278 : generic_join generic map(name => joinName, number_of_predecessors => 12, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(278), clk => clk, reset => reset); --
    end block;
    -- CP-element group 279:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	277 
    -- CP-element group 279: successors 
    -- CP-element group 279: marked-successors 
    -- CP-element group 279: 	277 
    -- CP-element group 279:  members (3) 
      -- CP-element group 279: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1330_Sample/ra
      -- CP-element group 279: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1330_Sample/$exit
      -- CP-element group 279: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1330_sample_completed_
      -- 
    ra_2985_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 279_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1330_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(279)); -- 
    -- CP-element group 280:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	278 
    -- CP-element group 280: successors 
    -- CP-element group 280: 	390 
    -- CP-element group 280: 	301 
    -- CP-element group 280: 	305 
    -- CP-element group 280: 	309 
    -- CP-element group 280: 	332 
    -- CP-element group 280: 	336 
    -- CP-element group 280: 	340 
    -- CP-element group 280: 	355 
    -- CP-element group 280: 	367 
    -- CP-element group 280: 	371 
    -- CP-element group 280: 	375 
    -- CP-element group 280: marked-successors 
    -- CP-element group 280: 	278 
    -- CP-element group 280:  members (3) 
      -- CP-element group 280: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1330_Update/$exit
      -- CP-element group 280: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1330_update_completed_
      -- CP-element group 280: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1330_Update/ca
      -- 
    ca_2990_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 280_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1330_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(280)); -- 
    -- CP-element group 281:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	228 
    -- CP-element group 281: 	244 
    -- CP-element group 281: 	252 
    -- CP-element group 281: marked-predecessors 
    -- CP-element group 281: 	283 
    -- CP-element group 281: successors 
    -- CP-element group 281: 	283 
    -- CP-element group 281:  members (3) 
      -- CP-element group 281: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1341_Sample/req
      -- CP-element group 281: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1341_Sample/$entry
      -- CP-element group 281: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1341_sample_start_
      -- 
    req_2998_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2998_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(281), ack => W_lorx_xlhsx_xfalse135_exec_guard_1228_delayed_1_0_1339_inst_req_0); -- 
    zeropad3D_A_cp_element_group_281: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_281"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(228) & zeropad3D_A_CP_1983_elements(244) & zeropad3D_A_CP_1983_elements(252) & zeropad3D_A_CP_1983_elements(283);
      gj_zeropad3D_A_cp_element_group_281 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(281), clk => clk, reset => reset); --
    end block;
    -- CP-element group 282:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: marked-predecessors 
    -- CP-element group 282: 	284 
    -- CP-element group 282: successors 
    -- CP-element group 282: 	284 
    -- CP-element group 282:  members (3) 
      -- CP-element group 282: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1341_Update/req
      -- CP-element group 282: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1341_Update/$entry
      -- CP-element group 282: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1341_update_start_
      -- 
    req_3003_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3003_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(282), ack => W_lorx_xlhsx_xfalse135_exec_guard_1228_delayed_1_0_1339_inst_req_1); -- 
    zeropad3D_A_cp_element_group_282: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_282"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= zeropad3D_A_CP_1983_elements(284);
      gj_zeropad3D_A_cp_element_group_282 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(282), clk => clk, reset => reset); --
    end block;
    -- CP-element group 283:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: 	281 
    -- CP-element group 283: successors 
    -- CP-element group 283: marked-successors 
    -- CP-element group 283: 	226 
    -- CP-element group 283: 	242 
    -- CP-element group 283: 	250 
    -- CP-element group 283: 	281 
    -- CP-element group 283:  members (3) 
      -- CP-element group 283: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1341_Sample/ack
      -- CP-element group 283: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1341_Sample/$exit
      -- CP-element group 283: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1341_sample_completed_
      -- 
    ack_2999_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 283_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_lorx_xlhsx_xfalse135_exec_guard_1228_delayed_1_0_1339_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(283)); -- 
    -- CP-element group 284:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	282 
    -- CP-element group 284: successors 
    -- CP-element group 284: 	404 
    -- CP-element group 284: marked-successors 
    -- CP-element group 284: 	282 
    -- CP-element group 284:  members (3) 
      -- CP-element group 284: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1341_Update/ack
      -- CP-element group 284: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1341_Update/$exit
      -- CP-element group 284: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1341_update_completed_
      -- 
    ack_3004_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 284_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_lorx_xlhsx_xfalse135_exec_guard_1228_delayed_1_0_1339_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(284)); -- 
    -- CP-element group 285:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: 	228 
    -- CP-element group 285: 	244 
    -- CP-element group 285: 	252 
    -- CP-element group 285: marked-predecessors 
    -- CP-element group 285: 	287 
    -- CP-element group 285: successors 
    -- CP-element group 285: 	287 
    -- CP-element group 285:  members (3) 
      -- CP-element group 285: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1350_Sample/req
      -- CP-element group 285: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1350_Sample/$entry
      -- CP-element group 285: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1350_sample_start_
      -- 
    req_3012_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3012_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(285), ack => W_lorx_xlhsx_xfalse135_exec_guard_1235_delayed_1_0_1348_inst_req_0); -- 
    zeropad3D_A_cp_element_group_285: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_285"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(228) & zeropad3D_A_CP_1983_elements(244) & zeropad3D_A_CP_1983_elements(252) & zeropad3D_A_CP_1983_elements(287);
      gj_zeropad3D_A_cp_element_group_285 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(285), clk => clk, reset => reset); --
    end block;
    -- CP-element group 286:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: marked-predecessors 
    -- CP-element group 286: 	392 
    -- CP-element group 286: 	288 
    -- CP-element group 286: 	334 
    -- CP-element group 286: 	338 
    -- CP-element group 286: 	342 
    -- CP-element group 286: 	357 
    -- CP-element group 286: 	369 
    -- CP-element group 286: 	373 
    -- CP-element group 286: 	377 
    -- CP-element group 286: successors 
    -- CP-element group 286: 	288 
    -- CP-element group 286:  members (3) 
      -- CP-element group 286: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1350_Update/req
      -- CP-element group 286: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1350_Update/$entry
      -- CP-element group 286: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1350_update_start_
      -- 
    req_3017_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3017_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(286), ack => W_lorx_xlhsx_xfalse135_exec_guard_1235_delayed_1_0_1348_inst_req_1); -- 
    zeropad3D_A_cp_element_group_286: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_286"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(392) & zeropad3D_A_CP_1983_elements(288) & zeropad3D_A_CP_1983_elements(334) & zeropad3D_A_CP_1983_elements(338) & zeropad3D_A_CP_1983_elements(342) & zeropad3D_A_CP_1983_elements(357) & zeropad3D_A_CP_1983_elements(369) & zeropad3D_A_CP_1983_elements(373) & zeropad3D_A_CP_1983_elements(377);
      gj_zeropad3D_A_cp_element_group_286 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(286), clk => clk, reset => reset); --
    end block;
    -- CP-element group 287:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	285 
    -- CP-element group 287: successors 
    -- CP-element group 287: marked-successors 
    -- CP-element group 287: 	226 
    -- CP-element group 287: 	242 
    -- CP-element group 287: 	250 
    -- CP-element group 287: 	285 
    -- CP-element group 287:  members (3) 
      -- CP-element group 287: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1350_Sample/ack
      -- CP-element group 287: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1350_Sample/$exit
      -- CP-element group 287: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1350_sample_completed_
      -- 
    ack_3013_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 287_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_lorx_xlhsx_xfalse135_exec_guard_1235_delayed_1_0_1348_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(287)); -- 
    -- CP-element group 288:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	286 
    -- CP-element group 288: successors 
    -- CP-element group 288: 	390 
    -- CP-element group 288: 	332 
    -- CP-element group 288: 	336 
    -- CP-element group 288: 	340 
    -- CP-element group 288: 	355 
    -- CP-element group 288: 	367 
    -- CP-element group 288: 	371 
    -- CP-element group 288: 	375 
    -- CP-element group 288: marked-successors 
    -- CP-element group 288: 	286 
    -- CP-element group 288:  members (3) 
      -- CP-element group 288: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1350_Update/ack
      -- CP-element group 288: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1350_Update/$exit
      -- CP-element group 288: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1350_update_completed_
      -- 
    ack_3018_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 288_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_lorx_xlhsx_xfalse135_exec_guard_1235_delayed_1_0_1348_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(288)); -- 
    -- CP-element group 289:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: 	228 
    -- CP-element group 289: 	244 
    -- CP-element group 289: 	252 
    -- CP-element group 289: marked-predecessors 
    -- CP-element group 289: 	291 
    -- CP-element group 289: successors 
    -- CP-element group 289: 	291 
    -- CP-element group 289:  members (3) 
      -- CP-element group 289: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1358_sample_start_
      -- CP-element group 289: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1358_Sample/req
      -- CP-element group 289: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1358_Sample/$entry
      -- 
    req_3026_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3026_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(289), ack => W_lorx_xlhsx_xfalse135_exec_guard_1240_delayed_1_0_1356_inst_req_0); -- 
    zeropad3D_A_cp_element_group_289: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_289"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(228) & zeropad3D_A_CP_1983_elements(244) & zeropad3D_A_CP_1983_elements(252) & zeropad3D_A_CP_1983_elements(291);
      gj_zeropad3D_A_cp_element_group_289 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(289), clk => clk, reset => reset); --
    end block;
    -- CP-element group 290:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: marked-predecessors 
    -- CP-element group 290: 	292 
    -- CP-element group 290: 	303 
    -- CP-element group 290: 	307 
    -- CP-element group 290: 	311 
    -- CP-element group 290: successors 
    -- CP-element group 290: 	292 
    -- CP-element group 290:  members (3) 
      -- CP-element group 290: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1358_Update/$entry
      -- CP-element group 290: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1358_Update/req
      -- CP-element group 290: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1358_update_start_
      -- 
    req_3031_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3031_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(290), ack => W_lorx_xlhsx_xfalse135_exec_guard_1240_delayed_1_0_1356_inst_req_1); -- 
    zeropad3D_A_cp_element_group_290: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_290"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(292) & zeropad3D_A_CP_1983_elements(303) & zeropad3D_A_CP_1983_elements(307) & zeropad3D_A_CP_1983_elements(311);
      gj_zeropad3D_A_cp_element_group_290 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(290), clk => clk, reset => reset); --
    end block;
    -- CP-element group 291:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	289 
    -- CP-element group 291: successors 
    -- CP-element group 291: marked-successors 
    -- CP-element group 291: 	226 
    -- CP-element group 291: 	242 
    -- CP-element group 291: 	250 
    -- CP-element group 291: 	289 
    -- CP-element group 291:  members (3) 
      -- CP-element group 291: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1358_Sample/ack
      -- CP-element group 291: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1358_sample_completed_
      -- CP-element group 291: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1358_Sample/$exit
      -- 
    ack_3027_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 291_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_lorx_xlhsx_xfalse135_exec_guard_1240_delayed_1_0_1356_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(291)); -- 
    -- CP-element group 292:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	290 
    -- CP-element group 292: successors 
    -- CP-element group 292: 	301 
    -- CP-element group 292: 	305 
    -- CP-element group 292: 	309 
    -- CP-element group 292: marked-successors 
    -- CP-element group 292: 	290 
    -- CP-element group 292:  members (3) 
      -- CP-element group 292: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1358_Update/$exit
      -- CP-element group 292: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1358_update_completed_
      -- CP-element group 292: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1358_Update/ack
      -- 
    ack_3032_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 292_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_lorx_xlhsx_xfalse135_exec_guard_1240_delayed_1_0_1356_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(292)); -- 
    -- CP-element group 293:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: 	228 
    -- CP-element group 293: 	244 
    -- CP-element group 293: 	256 
    -- CP-element group 293: marked-predecessors 
    -- CP-element group 293: 	295 
    -- CP-element group 293: successors 
    -- CP-element group 293: 	295 
    -- CP-element group 293:  members (3) 
      -- CP-element group 293: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1367_Sample/req
      -- CP-element group 293: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1367_Sample/$entry
      -- CP-element group 293: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1367_sample_start_
      -- 
    req_3040_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3040_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(293), ack => W_ifx_xend80_ifx_xthen152_taken_1246_delayed_1_0_1365_inst_req_0); -- 
    zeropad3D_A_cp_element_group_293: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_293"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(228) & zeropad3D_A_CP_1983_elements(244) & zeropad3D_A_CP_1983_elements(256) & zeropad3D_A_CP_1983_elements(295);
      gj_zeropad3D_A_cp_element_group_293 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(293), clk => clk, reset => reset); --
    end block;
    -- CP-element group 294:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: marked-predecessors 
    -- CP-element group 294: 	296 
    -- CP-element group 294: 	303 
    -- CP-element group 294: 	307 
    -- CP-element group 294: 	311 
    -- CP-element group 294: successors 
    -- CP-element group 294: 	296 
    -- CP-element group 294:  members (3) 
      -- CP-element group 294: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1367_Update/req
      -- CP-element group 294: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1367_Update/$entry
      -- CP-element group 294: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1367_update_start_
      -- 
    req_3045_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3045_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(294), ack => W_ifx_xend80_ifx_xthen152_taken_1246_delayed_1_0_1365_inst_req_1); -- 
    zeropad3D_A_cp_element_group_294: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_294"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(296) & zeropad3D_A_CP_1983_elements(303) & zeropad3D_A_CP_1983_elements(307) & zeropad3D_A_CP_1983_elements(311);
      gj_zeropad3D_A_cp_element_group_294 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(294), clk => clk, reset => reset); --
    end block;
    -- CP-element group 295:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 295: predecessors 
    -- CP-element group 295: 	293 
    -- CP-element group 295: successors 
    -- CP-element group 295: marked-successors 
    -- CP-element group 295: 	226 
    -- CP-element group 295: 	242 
    -- CP-element group 295: 	254 
    -- CP-element group 295: 	293 
    -- CP-element group 295:  members (3) 
      -- CP-element group 295: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1367_Sample/ack
      -- CP-element group 295: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1367_Sample/$exit
      -- CP-element group 295: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1367_sample_completed_
      -- 
    ack_3041_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 295_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xend80_ifx_xthen152_taken_1246_delayed_1_0_1365_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(295)); -- 
    -- CP-element group 296:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 296: predecessors 
    -- CP-element group 296: 	294 
    -- CP-element group 296: successors 
    -- CP-element group 296: 	301 
    -- CP-element group 296: 	305 
    -- CP-element group 296: 	309 
    -- CP-element group 296: marked-successors 
    -- CP-element group 296: 	294 
    -- CP-element group 296:  members (3) 
      -- CP-element group 296: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1367_Update/ack
      -- CP-element group 296: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1367_Update/$exit
      -- CP-element group 296: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1367_update_completed_
      -- 
    ack_3046_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 296_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xend80_ifx_xthen152_taken_1246_delayed_1_0_1365_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(296)); -- 
    -- CP-element group 297:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 297: predecessors 
    -- CP-element group 297: 	164 
    -- CP-element group 297: 	172 
    -- CP-element group 297: 	176 
    -- CP-element group 297: 	184 
    -- CP-element group 297: 	188 
    -- CP-element group 297: 	192 
    -- CP-element group 297: 	196 
    -- CP-element group 297: 	200 
    -- CP-element group 297: 	204 
    -- CP-element group 297: 	208 
    -- CP-element group 297: 	212 
    -- CP-element group 297: 	216 
    -- CP-element group 297: 	220 
    -- CP-element group 297: marked-predecessors 
    -- CP-element group 297: 	299 
    -- CP-element group 297: successors 
    -- CP-element group 297: 	299 
    -- CP-element group 297:  members (3) 
      -- CP-element group 297: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1375_sample_start_
      -- CP-element group 297: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1375_Sample/req
      -- CP-element group 297: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1375_Sample/$entry
      -- 
    req_3054_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3054_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(297), ack => W_add96_1252_delayed_2_0_1373_inst_req_0); -- 
    zeropad3D_A_cp_element_group_297: block -- 
      constant place_capacities: IntegerArray(0 to 13) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1);
      constant place_markings: IntegerArray(0 to 13)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 1);
      constant place_delays: IntegerArray(0 to 13) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_297"; 
      signal preds: BooleanArray(1 to 14); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(164) & zeropad3D_A_CP_1983_elements(172) & zeropad3D_A_CP_1983_elements(176) & zeropad3D_A_CP_1983_elements(184) & zeropad3D_A_CP_1983_elements(188) & zeropad3D_A_CP_1983_elements(192) & zeropad3D_A_CP_1983_elements(196) & zeropad3D_A_CP_1983_elements(200) & zeropad3D_A_CP_1983_elements(204) & zeropad3D_A_CP_1983_elements(208) & zeropad3D_A_CP_1983_elements(212) & zeropad3D_A_CP_1983_elements(216) & zeropad3D_A_CP_1983_elements(220) & zeropad3D_A_CP_1983_elements(299);
      gj_zeropad3D_A_cp_element_group_297 : generic_join generic map(name => joinName, number_of_predecessors => 14, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(297), clk => clk, reset => reset); --
    end block;
    -- CP-element group 298:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 298: predecessors 
    -- CP-element group 298: marked-predecessors 
    -- CP-element group 298: 	300 
    -- CP-element group 298: 	303 
    -- CP-element group 298: successors 
    -- CP-element group 298: 	300 
    -- CP-element group 298:  members (3) 
      -- CP-element group 298: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1375_update_start_
      -- CP-element group 298: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1375_Update/req
      -- CP-element group 298: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1375_Update/$entry
      -- 
    req_3059_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3059_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(298), ack => W_add96_1252_delayed_2_0_1373_inst_req_1); -- 
    zeropad3D_A_cp_element_group_298: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_298"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(300) & zeropad3D_A_CP_1983_elements(303);
      gj_zeropad3D_A_cp_element_group_298 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(298), clk => clk, reset => reset); --
    end block;
    -- CP-element group 299:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 299: predecessors 
    -- CP-element group 299: 	297 
    -- CP-element group 299: successors 
    -- CP-element group 299: marked-successors 
    -- CP-element group 299: 	162 
    -- CP-element group 299: 	170 
    -- CP-element group 299: 	174 
    -- CP-element group 299: 	182 
    -- CP-element group 299: 	186 
    -- CP-element group 299: 	190 
    -- CP-element group 299: 	194 
    -- CP-element group 299: 	198 
    -- CP-element group 299: 	202 
    -- CP-element group 299: 	206 
    -- CP-element group 299: 	210 
    -- CP-element group 299: 	214 
    -- CP-element group 299: 	218 
    -- CP-element group 299: 	297 
    -- CP-element group 299:  members (3) 
      -- CP-element group 299: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1375_sample_completed_
      -- CP-element group 299: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1375_Sample/ack
      -- CP-element group 299: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1375_Sample/$exit
      -- 
    ack_3055_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 299_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_add96_1252_delayed_2_0_1373_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(299)); -- 
    -- CP-element group 300:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 300: predecessors 
    -- CP-element group 300: 	298 
    -- CP-element group 300: successors 
    -- CP-element group 300: 	301 
    -- CP-element group 300: marked-successors 
    -- CP-element group 300: 	298 
    -- CP-element group 300:  members (3) 
      -- CP-element group 300: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1375_Update/ack
      -- CP-element group 300: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1375_Update/$exit
      -- CP-element group 300: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1375_update_completed_
      -- 
    ack_3060_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 300_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_add96_1252_delayed_2_0_1373_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(300)); -- 
    -- CP-element group 301:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 301: predecessors 
    -- CP-element group 301: 	264 
    -- CP-element group 301: 	280 
    -- CP-element group 301: 	292 
    -- CP-element group 301: 	296 
    -- CP-element group 301: 	300 
    -- CP-element group 301: marked-predecessors 
    -- CP-element group 301: 	303 
    -- CP-element group 301: successors 
    -- CP-element group 301: 	303 
    -- CP-element group 301:  members (3) 
      -- CP-element group 301: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1380_sample_start_
      -- CP-element group 301: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1380_Sample/rr
      -- CP-element group 301: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1380_Sample/$entry
      -- 
    rr_3068_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3068_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(301), ack => type_cast_1380_inst_req_0); -- 
    zeropad3D_A_cp_element_group_301: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_301"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(264) & zeropad3D_A_CP_1983_elements(280) & zeropad3D_A_CP_1983_elements(292) & zeropad3D_A_CP_1983_elements(296) & zeropad3D_A_CP_1983_elements(300) & zeropad3D_A_CP_1983_elements(303);
      gj_zeropad3D_A_cp_element_group_301 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(301), clk => clk, reset => reset); --
    end block;
    -- CP-element group 302:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 302: predecessors 
    -- CP-element group 302: marked-predecessors 
    -- CP-element group 302: 	304 
    -- CP-element group 302: 	315 
    -- CP-element group 302: successors 
    -- CP-element group 302: 	304 
    -- CP-element group 302:  members (3) 
      -- CP-element group 302: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1380_update_start_
      -- CP-element group 302: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1380_Update/$entry
      -- CP-element group 302: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1380_Update/cr
      -- 
    cr_3073_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3073_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(302), ack => type_cast_1380_inst_req_1); -- 
    zeropad3D_A_cp_element_group_302: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_302"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(304) & zeropad3D_A_CP_1983_elements(315);
      gj_zeropad3D_A_cp_element_group_302 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(302), clk => clk, reset => reset); --
    end block;
    -- CP-element group 303:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 303: predecessors 
    -- CP-element group 303: 	301 
    -- CP-element group 303: successors 
    -- CP-element group 303: marked-successors 
    -- CP-element group 303: 	262 
    -- CP-element group 303: 	278 
    -- CP-element group 303: 	290 
    -- CP-element group 303: 	294 
    -- CP-element group 303: 	298 
    -- CP-element group 303: 	301 
    -- CP-element group 303:  members (3) 
      -- CP-element group 303: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1380_Sample/$exit
      -- CP-element group 303: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1380_sample_completed_
      -- CP-element group 303: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1380_Sample/ra
      -- 
    ra_3069_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 303_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1380_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(303)); -- 
    -- CP-element group 304:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 304: predecessors 
    -- CP-element group 304: 	302 
    -- CP-element group 304: successors 
    -- CP-element group 304: 	313 
    -- CP-element group 304: marked-successors 
    -- CP-element group 304: 	302 
    -- CP-element group 304:  members (3) 
      -- CP-element group 304: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1380_update_completed_
      -- CP-element group 304: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1380_Update/$exit
      -- CP-element group 304: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1380_Update/ca
      -- 
    ca_3074_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 304_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1380_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(304)); -- 
    -- CP-element group 305:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 305: predecessors 
    -- CP-element group 305: 	264 
    -- CP-element group 305: 	280 
    -- CP-element group 305: 	292 
    -- CP-element group 305: 	296 
    -- CP-element group 305: marked-predecessors 
    -- CP-element group 305: 	307 
    -- CP-element group 305: successors 
    -- CP-element group 305: 	307 
    -- CP-element group 305:  members (3) 
      -- CP-element group 305: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1384_sample_start_
      -- CP-element group 305: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1384_Sample/$entry
      -- CP-element group 305: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1384_Sample/req
      -- 
    req_3082_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3082_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(305), ack => W_ifx_xthen152_exec_guard_1256_delayed_1_0_1382_inst_req_0); -- 
    zeropad3D_A_cp_element_group_305: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_305"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(264) & zeropad3D_A_CP_1983_elements(280) & zeropad3D_A_CP_1983_elements(292) & zeropad3D_A_CP_1983_elements(296) & zeropad3D_A_CP_1983_elements(307);
      gj_zeropad3D_A_cp_element_group_305 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(305), clk => clk, reset => reset); --
    end block;
    -- CP-element group 306:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 306: predecessors 
    -- CP-element group 306: marked-predecessors 
    -- CP-element group 306: 	308 
    -- CP-element group 306: successors 
    -- CP-element group 306: 	308 
    -- CP-element group 306:  members (3) 
      -- CP-element group 306: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1384_update_start_
      -- CP-element group 306: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1384_Update/$entry
      -- CP-element group 306: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1384_Update/req
      -- 
    req_3087_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3087_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(306), ack => W_ifx_xthen152_exec_guard_1256_delayed_1_0_1382_inst_req_1); -- 
    zeropad3D_A_cp_element_group_306: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_306"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= zeropad3D_A_CP_1983_elements(308);
      gj_zeropad3D_A_cp_element_group_306 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(306), clk => clk, reset => reset); --
    end block;
    -- CP-element group 307:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 307: predecessors 
    -- CP-element group 307: 	305 
    -- CP-element group 307: successors 
    -- CP-element group 307: marked-successors 
    -- CP-element group 307: 	262 
    -- CP-element group 307: 	278 
    -- CP-element group 307: 	290 
    -- CP-element group 307: 	294 
    -- CP-element group 307: 	305 
    -- CP-element group 307:  members (3) 
      -- CP-element group 307: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1384_sample_completed_
      -- CP-element group 307: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1384_Sample/$exit
      -- CP-element group 307: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1384_Sample/ack
      -- 
    ack_3083_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 307_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xthen152_exec_guard_1256_delayed_1_0_1382_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(307)); -- 
    -- CP-element group 308:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 308: predecessors 
    -- CP-element group 308: 	306 
    -- CP-element group 308: successors 
    -- CP-element group 308: 	404 
    -- CP-element group 308: marked-successors 
    -- CP-element group 308: 	306 
    -- CP-element group 308:  members (3) 
      -- CP-element group 308: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1384_update_completed_
      -- CP-element group 308: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1384_Update/$exit
      -- CP-element group 308: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1384_Update/ack
      -- 
    ack_3088_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 308_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xthen152_exec_guard_1256_delayed_1_0_1382_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(308)); -- 
    -- CP-element group 309:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 309: predecessors 
    -- CP-element group 309: 	264 
    -- CP-element group 309: 	280 
    -- CP-element group 309: 	292 
    -- CP-element group 309: 	296 
    -- CP-element group 309: marked-predecessors 
    -- CP-element group 309: 	311 
    -- CP-element group 309: successors 
    -- CP-element group 309: 	311 
    -- CP-element group 309:  members (3) 
      -- CP-element group 309: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1397_sample_start_
      -- CP-element group 309: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1397_Sample/$entry
      -- CP-element group 309: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1397_Sample/req
      -- 
    req_3096_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3096_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(309), ack => W_ifx_xthen152_exec_guard_1266_delayed_1_0_1395_inst_req_0); -- 
    zeropad3D_A_cp_element_group_309: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_309"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(264) & zeropad3D_A_CP_1983_elements(280) & zeropad3D_A_CP_1983_elements(292) & zeropad3D_A_CP_1983_elements(296) & zeropad3D_A_CP_1983_elements(311);
      gj_zeropad3D_A_cp_element_group_309 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(309), clk => clk, reset => reset); --
    end block;
    -- CP-element group 310:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 310: predecessors 
    -- CP-element group 310: marked-predecessors 
    -- CP-element group 310: 	312 
    -- CP-element group 310: 	315 
    -- CP-element group 310: successors 
    -- CP-element group 310: 	312 
    -- CP-element group 310:  members (3) 
      -- CP-element group 310: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1397_update_start_
      -- CP-element group 310: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1397_Update/$entry
      -- CP-element group 310: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1397_Update/req
      -- 
    req_3101_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3101_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(310), ack => W_ifx_xthen152_exec_guard_1266_delayed_1_0_1395_inst_req_1); -- 
    zeropad3D_A_cp_element_group_310: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_310"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(312) & zeropad3D_A_CP_1983_elements(315);
      gj_zeropad3D_A_cp_element_group_310 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(310), clk => clk, reset => reset); --
    end block;
    -- CP-element group 311:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 311: predecessors 
    -- CP-element group 311: 	309 
    -- CP-element group 311: successors 
    -- CP-element group 311: marked-successors 
    -- CP-element group 311: 	262 
    -- CP-element group 311: 	278 
    -- CP-element group 311: 	290 
    -- CP-element group 311: 	294 
    -- CP-element group 311: 	309 
    -- CP-element group 311:  members (3) 
      -- CP-element group 311: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1397_sample_completed_
      -- CP-element group 311: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1397_Sample/$exit
      -- CP-element group 311: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1397_Sample/ack
      -- 
    ack_3097_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 311_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xthen152_exec_guard_1266_delayed_1_0_1395_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(311)); -- 
    -- CP-element group 312:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 312: predecessors 
    -- CP-element group 312: 	310 
    -- CP-element group 312: successors 
    -- CP-element group 312: 	313 
    -- CP-element group 312: marked-successors 
    -- CP-element group 312: 	310 
    -- CP-element group 312:  members (3) 
      -- CP-element group 312: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1397_update_completed_
      -- CP-element group 312: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1397_Update/$exit
      -- CP-element group 312: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1397_Update/ack
      -- 
    ack_3102_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 312_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xthen152_exec_guard_1266_delayed_1_0_1395_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(312)); -- 
    -- CP-element group 313:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 313: predecessors 
    -- CP-element group 313: 	304 
    -- CP-element group 313: 	312 
    -- CP-element group 313: marked-predecessors 
    -- CP-element group 313: 	315 
    -- CP-element group 313: successors 
    -- CP-element group 313: 	315 
    -- CP-element group 313:  members (3) 
      -- CP-element group 313: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1402_sample_start_
      -- CP-element group 313: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1402_Sample/$entry
      -- CP-element group 313: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1402_Sample/rr
      -- 
    rr_3110_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3110_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(313), ack => type_cast_1402_inst_req_0); -- 
    zeropad3D_A_cp_element_group_313: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_313"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(304) & zeropad3D_A_CP_1983_elements(312) & zeropad3D_A_CP_1983_elements(315);
      gj_zeropad3D_A_cp_element_group_313 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(313), clk => clk, reset => reset); --
    end block;
    -- CP-element group 314:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 314: predecessors 
    -- CP-element group 314: marked-predecessors 
    -- CP-element group 314: 	316 
    -- CP-element group 314: 	320 
    -- CP-element group 314: successors 
    -- CP-element group 314: 	316 
    -- CP-element group 314:  members (3) 
      -- CP-element group 314: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1402_update_start_
      -- CP-element group 314: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1402_Update/$entry
      -- CP-element group 314: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1402_Update/cr
      -- 
    cr_3115_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3115_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(314), ack => type_cast_1402_inst_req_1); -- 
    zeropad3D_A_cp_element_group_314: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_314"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(316) & zeropad3D_A_CP_1983_elements(320);
      gj_zeropad3D_A_cp_element_group_314 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(314), clk => clk, reset => reset); --
    end block;
    -- CP-element group 315:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 315: predecessors 
    -- CP-element group 315: 	313 
    -- CP-element group 315: successors 
    -- CP-element group 315: marked-successors 
    -- CP-element group 315: 	302 
    -- CP-element group 315: 	310 
    -- CP-element group 315: 	313 
    -- CP-element group 315:  members (3) 
      -- CP-element group 315: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1402_sample_completed_
      -- CP-element group 315: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1402_Sample/$exit
      -- CP-element group 315: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1402_Sample/ra
      -- 
    ra_3111_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 315_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1402_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(315)); -- 
    -- CP-element group 316:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 316: predecessors 
    -- CP-element group 316: 	314 
    -- CP-element group 316: successors 
    -- CP-element group 316: 	320 
    -- CP-element group 316: marked-successors 
    -- CP-element group 316: 	314 
    -- CP-element group 316:  members (16) 
      -- CP-element group 316: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1402_update_completed_
      -- CP-element group 316: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1402_Update/$exit
      -- CP-element group 316: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1402_Update/ca
      -- CP-element group 316: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1408_index_resized_1
      -- CP-element group 316: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1408_index_scaled_1
      -- CP-element group 316: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1408_index_computed_1
      -- CP-element group 316: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1408_index_resize_1/$entry
      -- CP-element group 316: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1408_index_resize_1/$exit
      -- CP-element group 316: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1408_index_resize_1/index_resize_req
      -- CP-element group 316: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1408_index_resize_1/index_resize_ack
      -- CP-element group 316: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1408_index_scale_1/$entry
      -- CP-element group 316: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1408_index_scale_1/$exit
      -- CP-element group 316: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1408_index_scale_1/scale_rename_req
      -- CP-element group 316: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1408_index_scale_1/scale_rename_ack
      -- CP-element group 316: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1408_final_index_sum_regn_Sample/$entry
      -- CP-element group 316: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1408_final_index_sum_regn_Sample/req
      -- 
    ca_3116_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 316_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1402_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(316)); -- 
    req_3141_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3141_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(316), ack => array_obj_ref_1408_index_offset_req_0); -- 
    -- CP-element group 317:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 317: predecessors 
    -- CP-element group 317: 	321 
    -- CP-element group 317: marked-predecessors 
    -- CP-element group 317: 	322 
    -- CP-element group 317: successors 
    -- CP-element group 317: 	322 
    -- CP-element group 317:  members (3) 
      -- CP-element group 317: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/addr_of_1409_sample_start_
      -- CP-element group 317: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/addr_of_1409_request/$entry
      -- CP-element group 317: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/addr_of_1409_request/req
      -- 
    req_3156_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3156_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(317), ack => addr_of_1409_final_reg_req_0); -- 
    zeropad3D_A_cp_element_group_317: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_317"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(321) & zeropad3D_A_CP_1983_elements(322);
      gj_zeropad3D_A_cp_element_group_317 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(317), clk => clk, reset => reset); --
    end block;
    -- CP-element group 318:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 318: predecessors 
    -- CP-element group 318: 	42 
    -- CP-element group 318: marked-predecessors 
    -- CP-element group 318: 	323 
    -- CP-element group 318: 	326 
    -- CP-element group 318: successors 
    -- CP-element group 318: 	323 
    -- CP-element group 318:  members (3) 
      -- CP-element group 318: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/addr_of_1409_update_start_
      -- CP-element group 318: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/addr_of_1409_complete/$entry
      -- CP-element group 318: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/addr_of_1409_complete/req
      -- 
    req_3161_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3161_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(318), ack => addr_of_1409_final_reg_req_1); -- 
    zeropad3D_A_cp_element_group_318: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_318"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(42) & zeropad3D_A_CP_1983_elements(323) & zeropad3D_A_CP_1983_elements(326);
      gj_zeropad3D_A_cp_element_group_318 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(318), clk => clk, reset => reset); --
    end block;
    -- CP-element group 319:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 319: predecessors 
    -- CP-element group 319: 	42 
    -- CP-element group 319: marked-predecessors 
    -- CP-element group 319: 	321 
    -- CP-element group 319: 	322 
    -- CP-element group 319: successors 
    -- CP-element group 319: 	321 
    -- CP-element group 319:  members (3) 
      -- CP-element group 319: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1408_final_index_sum_regn_update_start
      -- CP-element group 319: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1408_final_index_sum_regn_Update/$entry
      -- CP-element group 319: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1408_final_index_sum_regn_Update/req
      -- 
    req_3146_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3146_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(319), ack => array_obj_ref_1408_index_offset_req_1); -- 
    zeropad3D_A_cp_element_group_319: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_319"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(42) & zeropad3D_A_CP_1983_elements(321) & zeropad3D_A_CP_1983_elements(322);
      gj_zeropad3D_A_cp_element_group_319 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(319), clk => clk, reset => reset); --
    end block;
    -- CP-element group 320:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 320: predecessors 
    -- CP-element group 320: 	316 
    -- CP-element group 320: successors 
    -- CP-element group 320: 	404 
    -- CP-element group 320: marked-successors 
    -- CP-element group 320: 	314 
    -- CP-element group 320:  members (3) 
      -- CP-element group 320: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1408_final_index_sum_regn_sample_complete
      -- CP-element group 320: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1408_final_index_sum_regn_Sample/$exit
      -- CP-element group 320: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1408_final_index_sum_regn_Sample/ack
      -- 
    ack_3142_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 320_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1408_index_offset_ack_0, ack => zeropad3D_A_CP_1983_elements(320)); -- 
    -- CP-element group 321:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 321: predecessors 
    -- CP-element group 321: 	319 
    -- CP-element group 321: successors 
    -- CP-element group 321: 	317 
    -- CP-element group 321: marked-successors 
    -- CP-element group 321: 	319 
    -- CP-element group 321:  members (8) 
      -- CP-element group 321: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1408_root_address_calculated
      -- CP-element group 321: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1408_offset_calculated
      -- CP-element group 321: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1408_final_index_sum_regn_Update/$exit
      -- CP-element group 321: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1408_final_index_sum_regn_Update/ack
      -- CP-element group 321: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1408_base_plus_offset/$entry
      -- CP-element group 321: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1408_base_plus_offset/$exit
      -- CP-element group 321: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1408_base_plus_offset/sum_rename_req
      -- CP-element group 321: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1408_base_plus_offset/sum_rename_ack
      -- 
    ack_3147_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 321_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1408_index_offset_ack_1, ack => zeropad3D_A_CP_1983_elements(321)); -- 
    -- CP-element group 322:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 322: predecessors 
    -- CP-element group 322: 	317 
    -- CP-element group 322: successors 
    -- CP-element group 322: marked-successors 
    -- CP-element group 322: 	317 
    -- CP-element group 322: 	319 
    -- CP-element group 322:  members (3) 
      -- CP-element group 322: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/addr_of_1409_sample_completed_
      -- CP-element group 322: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/addr_of_1409_request/$exit
      -- CP-element group 322: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/addr_of_1409_request/ack
      -- 
    ack_3157_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 322_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1409_final_reg_ack_0, ack => zeropad3D_A_CP_1983_elements(322)); -- 
    -- CP-element group 323:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 323: predecessors 
    -- CP-element group 323: 	318 
    -- CP-element group 323: successors 
    -- CP-element group 323: 	324 
    -- CP-element group 323: marked-successors 
    -- CP-element group 323: 	318 
    -- CP-element group 323:  members (19) 
      -- CP-element group 323: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/addr_of_1409_update_completed_
      -- CP-element group 323: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/addr_of_1409_complete/$exit
      -- CP-element group 323: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/addr_of_1409_complete/ack
      -- CP-element group 323: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1413_base_address_calculated
      -- CP-element group 323: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1413_word_address_calculated
      -- CP-element group 323: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1413_root_address_calculated
      -- CP-element group 323: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1413_base_address_resized
      -- CP-element group 323: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1413_base_addr_resize/$entry
      -- CP-element group 323: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1413_base_addr_resize/$exit
      -- CP-element group 323: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1413_base_addr_resize/base_resize_req
      -- CP-element group 323: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1413_base_addr_resize/base_resize_ack
      -- CP-element group 323: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1413_base_plus_offset/$entry
      -- CP-element group 323: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1413_base_plus_offset/$exit
      -- CP-element group 323: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1413_base_plus_offset/sum_rename_req
      -- CP-element group 323: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1413_base_plus_offset/sum_rename_ack
      -- CP-element group 323: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1413_word_addrgen/$entry
      -- CP-element group 323: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1413_word_addrgen/$exit
      -- CP-element group 323: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1413_word_addrgen/root_register_req
      -- CP-element group 323: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1413_word_addrgen/root_register_ack
      -- 
    ack_3162_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 323_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1409_final_reg_ack_1, ack => zeropad3D_A_CP_1983_elements(323)); -- 
    -- CP-element group 324:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 324: predecessors 
    -- CP-element group 324: 	323 
    -- CP-element group 324: marked-predecessors 
    -- CP-element group 324: 	400 
    -- CP-element group 324: 	326 
    -- CP-element group 324: successors 
    -- CP-element group 324: 	326 
    -- CP-element group 324:  members (9) 
      -- CP-element group 324: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1413_sample_start_
      -- CP-element group 324: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1413_Sample/$entry
      -- CP-element group 324: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1413_Sample/ptr_deref_1413_Split/$entry
      -- CP-element group 324: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1413_Sample/ptr_deref_1413_Split/$exit
      -- CP-element group 324: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1413_Sample/ptr_deref_1413_Split/split_req
      -- CP-element group 324: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1413_Sample/ptr_deref_1413_Split/split_ack
      -- CP-element group 324: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1413_Sample/word_access_start/$entry
      -- CP-element group 324: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1413_Sample/word_access_start/word_0/$entry
      -- CP-element group 324: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1413_Sample/word_access_start/word_0/rr
      -- 
    rr_3200_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3200_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(324), ack => ptr_deref_1413_store_0_req_0); -- 
    zeropad3D_A_cp_element_group_324: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_324"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(323) & zeropad3D_A_CP_1983_elements(400) & zeropad3D_A_CP_1983_elements(326);
      gj_zeropad3D_A_cp_element_group_324 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(324), clk => clk, reset => reset); --
    end block;
    -- CP-element group 325:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 325: predecessors 
    -- CP-element group 325: marked-predecessors 
    -- CP-element group 325: 	327 
    -- CP-element group 325: successors 
    -- CP-element group 325: 	327 
    -- CP-element group 325:  members (5) 
      -- CP-element group 325: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1413_update_start_
      -- CP-element group 325: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1413_Update/$entry
      -- CP-element group 325: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1413_Update/word_access_complete/$entry
      -- CP-element group 325: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1413_Update/word_access_complete/word_0/$entry
      -- CP-element group 325: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1413_Update/word_access_complete/word_0/cr
      -- 
    cr_3211_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3211_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(325), ack => ptr_deref_1413_store_0_req_1); -- 
    zeropad3D_A_cp_element_group_325: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_325"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= zeropad3D_A_CP_1983_elements(327);
      gj_zeropad3D_A_cp_element_group_325 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(325), clk => clk, reset => reset); --
    end block;
    -- CP-element group 326:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 326: predecessors 
    -- CP-element group 326: 	324 
    -- CP-element group 326: successors 
    -- CP-element group 326: 	403 
    -- CP-element group 326: marked-successors 
    -- CP-element group 326: 	318 
    -- CP-element group 326: 	324 
    -- CP-element group 326:  members (5) 
      -- CP-element group 326: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1413_sample_completed_
      -- CP-element group 326: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1413_Sample/$exit
      -- CP-element group 326: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1413_Sample/word_access_start/$exit
      -- CP-element group 326: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1413_Sample/word_access_start/word_0/$exit
      -- CP-element group 326: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1413_Sample/word_access_start/word_0/ra
      -- 
    ra_3201_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 326_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1413_store_0_ack_0, ack => zeropad3D_A_CP_1983_elements(326)); -- 
    -- CP-element group 327:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 327: predecessors 
    -- CP-element group 327: 	325 
    -- CP-element group 327: successors 
    -- CP-element group 327: 	404 
    -- CP-element group 327: marked-successors 
    -- CP-element group 327: 	325 
    -- CP-element group 327:  members (5) 
      -- CP-element group 327: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1413_update_completed_
      -- CP-element group 327: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1413_Update/$exit
      -- CP-element group 327: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1413_Update/word_access_complete/$exit
      -- CP-element group 327: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1413_Update/word_access_complete/word_0/$exit
      -- CP-element group 327: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1413_Update/word_access_complete/word_0/ca
      -- 
    ca_3212_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 327_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1413_store_0_ack_1, ack => zeropad3D_A_CP_1983_elements(327)); -- 
    -- CP-element group 328:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 328: predecessors 
    -- CP-element group 328: 	164 
    -- CP-element group 328: 	172 
    -- CP-element group 328: 	176 
    -- CP-element group 328: 	184 
    -- CP-element group 328: 	188 
    -- CP-element group 328: 	192 
    -- CP-element group 328: 	196 
    -- CP-element group 328: 	200 
    -- CP-element group 328: 	204 
    -- CP-element group 328: 	208 
    -- CP-element group 328: 	212 
    -- CP-element group 328: 	216 
    -- CP-element group 328: 	220 
    -- CP-element group 328: marked-predecessors 
    -- CP-element group 328: 	330 
    -- CP-element group 328: successors 
    -- CP-element group 328: 	330 
    -- CP-element group 328:  members (3) 
      -- CP-element group 328: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1422_sample_start_
      -- CP-element group 328: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1422_Sample/$entry
      -- CP-element group 328: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1422_Sample/req
      -- 
    req_3220_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3220_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(328), ack => W_add118_1290_delayed_2_0_1420_inst_req_0); -- 
    zeropad3D_A_cp_element_group_328: block -- 
      constant place_capacities: IntegerArray(0 to 13) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1);
      constant place_markings: IntegerArray(0 to 13)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 1);
      constant place_delays: IntegerArray(0 to 13) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_328"; 
      signal preds: BooleanArray(1 to 14); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(164) & zeropad3D_A_CP_1983_elements(172) & zeropad3D_A_CP_1983_elements(176) & zeropad3D_A_CP_1983_elements(184) & zeropad3D_A_CP_1983_elements(188) & zeropad3D_A_CP_1983_elements(192) & zeropad3D_A_CP_1983_elements(196) & zeropad3D_A_CP_1983_elements(200) & zeropad3D_A_CP_1983_elements(204) & zeropad3D_A_CP_1983_elements(208) & zeropad3D_A_CP_1983_elements(212) & zeropad3D_A_CP_1983_elements(216) & zeropad3D_A_CP_1983_elements(220) & zeropad3D_A_CP_1983_elements(330);
      gj_zeropad3D_A_cp_element_group_328 : generic_join generic map(name => joinName, number_of_predecessors => 14, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(328), clk => clk, reset => reset); --
    end block;
    -- CP-element group 329:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 329: predecessors 
    -- CP-element group 329: marked-predecessors 
    -- CP-element group 329: 	331 
    -- CP-element group 329: 	334 
    -- CP-element group 329: successors 
    -- CP-element group 329: 	331 
    -- CP-element group 329:  members (3) 
      -- CP-element group 329: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1422_update_start_
      -- CP-element group 329: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1422_Update/$entry
      -- CP-element group 329: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1422_Update/req
      -- 
    req_3225_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3225_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(329), ack => W_add118_1290_delayed_2_0_1420_inst_req_1); -- 
    zeropad3D_A_cp_element_group_329: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_329"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(331) & zeropad3D_A_CP_1983_elements(334);
      gj_zeropad3D_A_cp_element_group_329 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(329), clk => clk, reset => reset); --
    end block;
    -- CP-element group 330:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 330: predecessors 
    -- CP-element group 330: 	328 
    -- CP-element group 330: successors 
    -- CP-element group 330: marked-successors 
    -- CP-element group 330: 	162 
    -- CP-element group 330: 	170 
    -- CP-element group 330: 	174 
    -- CP-element group 330: 	182 
    -- CP-element group 330: 	186 
    -- CP-element group 330: 	190 
    -- CP-element group 330: 	194 
    -- CP-element group 330: 	198 
    -- CP-element group 330: 	202 
    -- CP-element group 330: 	206 
    -- CP-element group 330: 	210 
    -- CP-element group 330: 	214 
    -- CP-element group 330: 	218 
    -- CP-element group 330: 	328 
    -- CP-element group 330:  members (3) 
      -- CP-element group 330: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1422_sample_completed_
      -- CP-element group 330: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1422_Sample/$exit
      -- CP-element group 330: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1422_Sample/ack
      -- 
    ack_3221_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 330_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_add118_1290_delayed_2_0_1420_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(330)); -- 
    -- CP-element group 331:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 331: predecessors 
    -- CP-element group 331: 	329 
    -- CP-element group 331: successors 
    -- CP-element group 331: 	332 
    -- CP-element group 331: marked-successors 
    -- CP-element group 331: 	329 
    -- CP-element group 331:  members (3) 
      -- CP-element group 331: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1422_update_completed_
      -- CP-element group 331: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1422_Update/$exit
      -- CP-element group 331: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1422_Update/ack
      -- 
    ack_3226_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 331_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_add118_1290_delayed_2_0_1420_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(331)); -- 
    -- CP-element group 332:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 332: predecessors 
    -- CP-element group 332: 	264 
    -- CP-element group 332: 	280 
    -- CP-element group 332: 	288 
    -- CP-element group 332: 	331 
    -- CP-element group 332: marked-predecessors 
    -- CP-element group 332: 	334 
    -- CP-element group 332: successors 
    -- CP-element group 332: 	334 
    -- CP-element group 332:  members (3) 
      -- CP-element group 332: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1427_sample_start_
      -- CP-element group 332: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1427_Sample/$entry
      -- CP-element group 332: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1427_Sample/rr
      -- 
    rr_3234_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3234_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(332), ack => type_cast_1427_inst_req_0); -- 
    zeropad3D_A_cp_element_group_332: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_332"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(264) & zeropad3D_A_CP_1983_elements(280) & zeropad3D_A_CP_1983_elements(288) & zeropad3D_A_CP_1983_elements(331) & zeropad3D_A_CP_1983_elements(334);
      gj_zeropad3D_A_cp_element_group_332 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(332), clk => clk, reset => reset); --
    end block;
    -- CP-element group 333:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 333: predecessors 
    -- CP-element group 333: marked-predecessors 
    -- CP-element group 333: 	335 
    -- CP-element group 333: 	346 
    -- CP-element group 333: successors 
    -- CP-element group 333: 	335 
    -- CP-element group 333:  members (3) 
      -- CP-element group 333: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1427_update_start_
      -- CP-element group 333: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1427_Update/$entry
      -- CP-element group 333: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1427_Update/cr
      -- 
    cr_3239_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3239_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(333), ack => type_cast_1427_inst_req_1); -- 
    zeropad3D_A_cp_element_group_333: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_333"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(335) & zeropad3D_A_CP_1983_elements(346);
      gj_zeropad3D_A_cp_element_group_333 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(333), clk => clk, reset => reset); --
    end block;
    -- CP-element group 334:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 334: predecessors 
    -- CP-element group 334: 	332 
    -- CP-element group 334: successors 
    -- CP-element group 334: marked-successors 
    -- CP-element group 334: 	262 
    -- CP-element group 334: 	278 
    -- CP-element group 334: 	286 
    -- CP-element group 334: 	329 
    -- CP-element group 334: 	332 
    -- CP-element group 334:  members (3) 
      -- CP-element group 334: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1427_sample_completed_
      -- CP-element group 334: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1427_Sample/$exit
      -- CP-element group 334: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1427_Sample/ra
      -- 
    ra_3235_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 334_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1427_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(334)); -- 
    -- CP-element group 335:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 335: predecessors 
    -- CP-element group 335: 	333 
    -- CP-element group 335: successors 
    -- CP-element group 335: 	344 
    -- CP-element group 335: marked-successors 
    -- CP-element group 335: 	333 
    -- CP-element group 335:  members (3) 
      -- CP-element group 335: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1427_update_completed_
      -- CP-element group 335: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1427_Update/$exit
      -- CP-element group 335: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1427_Update/ca
      -- 
    ca_3240_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 335_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1427_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(335)); -- 
    -- CP-element group 336:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 336: predecessors 
    -- CP-element group 336: 	264 
    -- CP-element group 336: 	280 
    -- CP-element group 336: 	288 
    -- CP-element group 336: marked-predecessors 
    -- CP-element group 336: 	338 
    -- CP-element group 336: successors 
    -- CP-element group 336: 	338 
    -- CP-element group 336:  members (3) 
      -- CP-element group 336: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1431_sample_start_
      -- CP-element group 336: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1431_Sample/$entry
      -- CP-element group 336: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1431_Sample/req
      -- 
    req_3248_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3248_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(336), ack => W_ifx_xelse155_exec_guard_1294_delayed_1_0_1429_inst_req_0); -- 
    zeropad3D_A_cp_element_group_336: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_336"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(264) & zeropad3D_A_CP_1983_elements(280) & zeropad3D_A_CP_1983_elements(288) & zeropad3D_A_CP_1983_elements(338);
      gj_zeropad3D_A_cp_element_group_336 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(336), clk => clk, reset => reset); --
    end block;
    -- CP-element group 337:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 337: predecessors 
    -- CP-element group 337: marked-predecessors 
    -- CP-element group 337: 	339 
    -- CP-element group 337: successors 
    -- CP-element group 337: 	339 
    -- CP-element group 337:  members (3) 
      -- CP-element group 337: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1431_update_start_
      -- CP-element group 337: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1431_Update/$entry
      -- CP-element group 337: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1431_Update/req
      -- 
    req_3253_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3253_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(337), ack => W_ifx_xelse155_exec_guard_1294_delayed_1_0_1429_inst_req_1); -- 
    zeropad3D_A_cp_element_group_337: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_337"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= zeropad3D_A_CP_1983_elements(339);
      gj_zeropad3D_A_cp_element_group_337 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(337), clk => clk, reset => reset); --
    end block;
    -- CP-element group 338:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 338: predecessors 
    -- CP-element group 338: 	336 
    -- CP-element group 338: successors 
    -- CP-element group 338: marked-successors 
    -- CP-element group 338: 	262 
    -- CP-element group 338: 	278 
    -- CP-element group 338: 	286 
    -- CP-element group 338: 	336 
    -- CP-element group 338:  members (3) 
      -- CP-element group 338: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1431_sample_completed_
      -- CP-element group 338: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1431_Sample/$exit
      -- CP-element group 338: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1431_Sample/ack
      -- 
    ack_3249_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 338_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xelse155_exec_guard_1294_delayed_1_0_1429_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(338)); -- 
    -- CP-element group 339:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 339: predecessors 
    -- CP-element group 339: 	337 
    -- CP-element group 339: successors 
    -- CP-element group 339: 	404 
    -- CP-element group 339: marked-successors 
    -- CP-element group 339: 	337 
    -- CP-element group 339:  members (3) 
      -- CP-element group 339: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1431_update_completed_
      -- CP-element group 339: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1431_Update/$exit
      -- CP-element group 339: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1431_Update/ack
      -- 
    ack_3254_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 339_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xelse155_exec_guard_1294_delayed_1_0_1429_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(339)); -- 
    -- CP-element group 340:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 340: predecessors 
    -- CP-element group 340: 	264 
    -- CP-element group 340: 	280 
    -- CP-element group 340: 	288 
    -- CP-element group 340: marked-predecessors 
    -- CP-element group 340: 	342 
    -- CP-element group 340: successors 
    -- CP-element group 340: 	342 
    -- CP-element group 340:  members (3) 
      -- CP-element group 340: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1444_sample_start_
      -- CP-element group 340: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1444_Sample/$entry
      -- CP-element group 340: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1444_Sample/req
      -- 
    req_3262_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3262_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(340), ack => W_ifx_xelse155_exec_guard_1304_delayed_1_0_1442_inst_req_0); -- 
    zeropad3D_A_cp_element_group_340: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_340"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(264) & zeropad3D_A_CP_1983_elements(280) & zeropad3D_A_CP_1983_elements(288) & zeropad3D_A_CP_1983_elements(342);
      gj_zeropad3D_A_cp_element_group_340 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(340), clk => clk, reset => reset); --
    end block;
    -- CP-element group 341:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 341: predecessors 
    -- CP-element group 341: marked-predecessors 
    -- CP-element group 341: 	343 
    -- CP-element group 341: 	346 
    -- CP-element group 341: successors 
    -- CP-element group 341: 	343 
    -- CP-element group 341:  members (3) 
      -- CP-element group 341: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1444_update_start_
      -- CP-element group 341: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1444_Update/$entry
      -- CP-element group 341: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1444_Update/req
      -- 
    req_3267_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3267_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(341), ack => W_ifx_xelse155_exec_guard_1304_delayed_1_0_1442_inst_req_1); -- 
    zeropad3D_A_cp_element_group_341: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_341"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(343) & zeropad3D_A_CP_1983_elements(346);
      gj_zeropad3D_A_cp_element_group_341 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(341), clk => clk, reset => reset); --
    end block;
    -- CP-element group 342:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 342: predecessors 
    -- CP-element group 342: 	340 
    -- CP-element group 342: successors 
    -- CP-element group 342: marked-successors 
    -- CP-element group 342: 	262 
    -- CP-element group 342: 	278 
    -- CP-element group 342: 	286 
    -- CP-element group 342: 	340 
    -- CP-element group 342:  members (3) 
      -- CP-element group 342: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1444_sample_completed_
      -- CP-element group 342: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1444_Sample/$exit
      -- CP-element group 342: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1444_Sample/ack
      -- 
    ack_3263_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 342_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xelse155_exec_guard_1304_delayed_1_0_1442_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(342)); -- 
    -- CP-element group 343:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 343: predecessors 
    -- CP-element group 343: 	341 
    -- CP-element group 343: successors 
    -- CP-element group 343: 	344 
    -- CP-element group 343: marked-successors 
    -- CP-element group 343: 	341 
    -- CP-element group 343:  members (3) 
      -- CP-element group 343: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1444_update_completed_
      -- CP-element group 343: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1444_Update/$exit
      -- CP-element group 343: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1444_Update/ack
      -- 
    ack_3268_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 343_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xelse155_exec_guard_1304_delayed_1_0_1442_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(343)); -- 
    -- CP-element group 344:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 344: predecessors 
    -- CP-element group 344: 	335 
    -- CP-element group 344: 	343 
    -- CP-element group 344: marked-predecessors 
    -- CP-element group 344: 	346 
    -- CP-element group 344: successors 
    -- CP-element group 344: 	346 
    -- CP-element group 344:  members (3) 
      -- CP-element group 344: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1449_sample_start_
      -- CP-element group 344: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1449_Sample/$entry
      -- CP-element group 344: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1449_Sample/rr
      -- 
    rr_3276_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3276_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(344), ack => type_cast_1449_inst_req_0); -- 
    zeropad3D_A_cp_element_group_344: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_344"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(335) & zeropad3D_A_CP_1983_elements(343) & zeropad3D_A_CP_1983_elements(346);
      gj_zeropad3D_A_cp_element_group_344 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(344), clk => clk, reset => reset); --
    end block;
    -- CP-element group 345:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 345: predecessors 
    -- CP-element group 345: marked-predecessors 
    -- CP-element group 345: 	347 
    -- CP-element group 345: 	351 
    -- CP-element group 345: successors 
    -- CP-element group 345: 	347 
    -- CP-element group 345:  members (3) 
      -- CP-element group 345: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1449_update_start_
      -- CP-element group 345: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1449_Update/$entry
      -- CP-element group 345: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1449_Update/cr
      -- 
    cr_3281_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3281_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(345), ack => type_cast_1449_inst_req_1); -- 
    zeropad3D_A_cp_element_group_345: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_345"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(347) & zeropad3D_A_CP_1983_elements(351);
      gj_zeropad3D_A_cp_element_group_345 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(345), clk => clk, reset => reset); --
    end block;
    -- CP-element group 346:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 346: predecessors 
    -- CP-element group 346: 	344 
    -- CP-element group 346: successors 
    -- CP-element group 346: marked-successors 
    -- CP-element group 346: 	333 
    -- CP-element group 346: 	341 
    -- CP-element group 346: 	344 
    -- CP-element group 346:  members (3) 
      -- CP-element group 346: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1449_sample_completed_
      -- CP-element group 346: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1449_Sample/$exit
      -- CP-element group 346: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1449_Sample/ra
      -- 
    ra_3277_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 346_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1449_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(346)); -- 
    -- CP-element group 347:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 347: predecessors 
    -- CP-element group 347: 	345 
    -- CP-element group 347: successors 
    -- CP-element group 347: 	351 
    -- CP-element group 347: marked-successors 
    -- CP-element group 347: 	345 
    -- CP-element group 347:  members (16) 
      -- CP-element group 347: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1449_update_completed_
      -- CP-element group 347: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1449_Update/$exit
      -- CP-element group 347: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1449_Update/ca
      -- CP-element group 347: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1455_index_resized_1
      -- CP-element group 347: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1455_index_scaled_1
      -- CP-element group 347: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1455_index_computed_1
      -- CP-element group 347: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1455_index_resize_1/$entry
      -- CP-element group 347: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1455_index_resize_1/$exit
      -- CP-element group 347: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1455_index_resize_1/index_resize_req
      -- CP-element group 347: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1455_index_resize_1/index_resize_ack
      -- CP-element group 347: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1455_index_scale_1/$entry
      -- CP-element group 347: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1455_index_scale_1/$exit
      -- CP-element group 347: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1455_index_scale_1/scale_rename_req
      -- CP-element group 347: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1455_index_scale_1/scale_rename_ack
      -- CP-element group 347: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1455_final_index_sum_regn_Sample/$entry
      -- CP-element group 347: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1455_final_index_sum_regn_Sample/req
      -- 
    ca_3282_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 347_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1449_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(347)); -- 
    req_3307_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3307_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(347), ack => array_obj_ref_1455_index_offset_req_0); -- 
    -- CP-element group 348:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 348: predecessors 
    -- CP-element group 348: 	352 
    -- CP-element group 348: marked-predecessors 
    -- CP-element group 348: 	353 
    -- CP-element group 348: successors 
    -- CP-element group 348: 	353 
    -- CP-element group 348:  members (3) 
      -- CP-element group 348: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/addr_of_1456_sample_start_
      -- CP-element group 348: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/addr_of_1456_request/$entry
      -- CP-element group 348: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/addr_of_1456_request/req
      -- 
    req_3322_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3322_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(348), ack => addr_of_1456_final_reg_req_0); -- 
    zeropad3D_A_cp_element_group_348: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_348"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(352) & zeropad3D_A_CP_1983_elements(353);
      gj_zeropad3D_A_cp_element_group_348 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(348), clk => clk, reset => reset); --
    end block;
    -- CP-element group 349:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 349: predecessors 
    -- CP-element group 349: 	42 
    -- CP-element group 349: marked-predecessors 
    -- CP-element group 349: 	354 
    -- CP-element group 349: 	361 
    -- CP-element group 349: successors 
    -- CP-element group 349: 	354 
    -- CP-element group 349:  members (3) 
      -- CP-element group 349: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/addr_of_1456_update_start_
      -- CP-element group 349: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/addr_of_1456_complete/$entry
      -- CP-element group 349: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/addr_of_1456_complete/req
      -- 
    req_3327_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3327_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(349), ack => addr_of_1456_final_reg_req_1); -- 
    zeropad3D_A_cp_element_group_349: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_349"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(42) & zeropad3D_A_CP_1983_elements(354) & zeropad3D_A_CP_1983_elements(361);
      gj_zeropad3D_A_cp_element_group_349 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(349), clk => clk, reset => reset); --
    end block;
    -- CP-element group 350:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 350: predecessors 
    -- CP-element group 350: 	42 
    -- CP-element group 350: marked-predecessors 
    -- CP-element group 350: 	352 
    -- CP-element group 350: 	353 
    -- CP-element group 350: successors 
    -- CP-element group 350: 	352 
    -- CP-element group 350:  members (3) 
      -- CP-element group 350: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1455_final_index_sum_regn_update_start
      -- CP-element group 350: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1455_final_index_sum_regn_Update/$entry
      -- CP-element group 350: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1455_final_index_sum_regn_Update/req
      -- 
    req_3312_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3312_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(350), ack => array_obj_ref_1455_index_offset_req_1); -- 
    zeropad3D_A_cp_element_group_350: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_350"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(42) & zeropad3D_A_CP_1983_elements(352) & zeropad3D_A_CP_1983_elements(353);
      gj_zeropad3D_A_cp_element_group_350 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(350), clk => clk, reset => reset); --
    end block;
    -- CP-element group 351:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 351: predecessors 
    -- CP-element group 351: 	347 
    -- CP-element group 351: successors 
    -- CP-element group 351: 	404 
    -- CP-element group 351: marked-successors 
    -- CP-element group 351: 	345 
    -- CP-element group 351:  members (3) 
      -- CP-element group 351: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1455_final_index_sum_regn_sample_complete
      -- CP-element group 351: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1455_final_index_sum_regn_Sample/$exit
      -- CP-element group 351: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1455_final_index_sum_regn_Sample/ack
      -- 
    ack_3308_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 351_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1455_index_offset_ack_0, ack => zeropad3D_A_CP_1983_elements(351)); -- 
    -- CP-element group 352:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 352: predecessors 
    -- CP-element group 352: 	350 
    -- CP-element group 352: successors 
    -- CP-element group 352: 	348 
    -- CP-element group 352: marked-successors 
    -- CP-element group 352: 	350 
    -- CP-element group 352:  members (8) 
      -- CP-element group 352: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1455_root_address_calculated
      -- CP-element group 352: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1455_offset_calculated
      -- CP-element group 352: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1455_final_index_sum_regn_Update/$exit
      -- CP-element group 352: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1455_final_index_sum_regn_Update/ack
      -- CP-element group 352: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1455_base_plus_offset/$entry
      -- CP-element group 352: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1455_base_plus_offset/$exit
      -- CP-element group 352: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1455_base_plus_offset/sum_rename_req
      -- CP-element group 352: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1455_base_plus_offset/sum_rename_ack
      -- 
    ack_3313_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 352_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1455_index_offset_ack_1, ack => zeropad3D_A_CP_1983_elements(352)); -- 
    -- CP-element group 353:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 353: predecessors 
    -- CP-element group 353: 	348 
    -- CP-element group 353: successors 
    -- CP-element group 353: marked-successors 
    -- CP-element group 353: 	348 
    -- CP-element group 353: 	350 
    -- CP-element group 353:  members (3) 
      -- CP-element group 353: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/addr_of_1456_sample_completed_
      -- CP-element group 353: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/addr_of_1456_request/$exit
      -- CP-element group 353: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/addr_of_1456_request/ack
      -- 
    ack_3323_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 353_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1456_final_reg_ack_0, ack => zeropad3D_A_CP_1983_elements(353)); -- 
    -- CP-element group 354:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 354: predecessors 
    -- CP-element group 354: 	349 
    -- CP-element group 354: successors 
    -- CP-element group 354: 	359 
    -- CP-element group 354: marked-successors 
    -- CP-element group 354: 	349 
    -- CP-element group 354:  members (19) 
      -- CP-element group 354: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1464_base_addr_resize/$exit
      -- CP-element group 354: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1464_base_addr_resize/$entry
      -- CP-element group 354: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1464_word_addrgen/root_register_req
      -- CP-element group 354: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1464_base_addr_resize/base_resize_req
      -- CP-element group 354: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1464_base_addr_resize/base_resize_ack
      -- CP-element group 354: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1464_word_addrgen/root_register_ack
      -- CP-element group 354: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1464_base_plus_offset/$entry
      -- CP-element group 354: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1464_base_address_resized
      -- CP-element group 354: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1464_word_addrgen/$exit
      -- CP-element group 354: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1464_word_addrgen/$entry
      -- CP-element group 354: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1464_base_plus_offset/sum_rename_ack
      -- CP-element group 354: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1464_base_plus_offset/sum_rename_req
      -- CP-element group 354: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1464_base_plus_offset/$exit
      -- CP-element group 354: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1464_root_address_calculated
      -- CP-element group 354: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/addr_of_1456_update_completed_
      -- CP-element group 354: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1464_word_address_calculated
      -- CP-element group 354: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1464_base_address_calculated
      -- CP-element group 354: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/addr_of_1456_complete/$exit
      -- CP-element group 354: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/addr_of_1456_complete/ack
      -- 
    ack_3328_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 354_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1456_final_reg_ack_1, ack => zeropad3D_A_CP_1983_elements(354)); -- 
    -- CP-element group 355:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 355: predecessors 
    -- CP-element group 355: 	264 
    -- CP-element group 355: 	280 
    -- CP-element group 355: 	288 
    -- CP-element group 355: marked-predecessors 
    -- CP-element group 355: 	357 
    -- CP-element group 355: successors 
    -- CP-element group 355: 	357 
    -- CP-element group 355:  members (3) 
      -- CP-element group 355: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1460_sample_start_
      -- CP-element group 355: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1460_Sample/$entry
      -- CP-element group 355: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1460_Sample/req
      -- 
    req_3336_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3336_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(355), ack => W_ifx_xelse155_exec_guard_1317_delayed_9_0_1458_inst_req_0); -- 
    zeropad3D_A_cp_element_group_355: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_355"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(264) & zeropad3D_A_CP_1983_elements(280) & zeropad3D_A_CP_1983_elements(288) & zeropad3D_A_CP_1983_elements(357);
      gj_zeropad3D_A_cp_element_group_355 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(355), clk => clk, reset => reset); --
    end block;
    -- CP-element group 356:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 356: predecessors 
    -- CP-element group 356: marked-predecessors 
    -- CP-element group 356: 	358 
    -- CP-element group 356: 	361 
    -- CP-element group 356: successors 
    -- CP-element group 356: 	358 
    -- CP-element group 356:  members (3) 
      -- CP-element group 356: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1460_update_start_
      -- CP-element group 356: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1460_Update/$entry
      -- CP-element group 356: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1460_Update/req
      -- 
    req_3341_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3341_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(356), ack => W_ifx_xelse155_exec_guard_1317_delayed_9_0_1458_inst_req_1); -- 
    zeropad3D_A_cp_element_group_356: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_356"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(358) & zeropad3D_A_CP_1983_elements(361);
      gj_zeropad3D_A_cp_element_group_356 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(356), clk => clk, reset => reset); --
    end block;
    -- CP-element group 357:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 357: predecessors 
    -- CP-element group 357: 	355 
    -- CP-element group 357: successors 
    -- CP-element group 357: marked-successors 
    -- CP-element group 357: 	262 
    -- CP-element group 357: 	278 
    -- CP-element group 357: 	286 
    -- CP-element group 357: 	355 
    -- CP-element group 357:  members (3) 
      -- CP-element group 357: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1460_sample_completed_
      -- CP-element group 357: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1460_Sample/$exit
      -- CP-element group 357: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1460_Sample/ack
      -- 
    ack_3337_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 357_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xelse155_exec_guard_1317_delayed_9_0_1458_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(357)); -- 
    -- CP-element group 358:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 358: predecessors 
    -- CP-element group 358: 	356 
    -- CP-element group 358: successors 
    -- CP-element group 358: 	359 
    -- CP-element group 358: marked-successors 
    -- CP-element group 358: 	356 
    -- CP-element group 358:  members (3) 
      -- CP-element group 358: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1460_update_completed_
      -- CP-element group 358: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1460_Update/$exit
      -- CP-element group 358: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1460_Update/ack
      -- 
    ack_3342_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 358_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xelse155_exec_guard_1317_delayed_9_0_1458_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(358)); -- 
    -- CP-element group 359:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 359: predecessors 
    -- CP-element group 359: 	354 
    -- CP-element group 359: 	358 
    -- CP-element group 359: marked-predecessors 
    -- CP-element group 359: 	361 
    -- CP-element group 359: successors 
    -- CP-element group 359: 	361 
    -- CP-element group 359:  members (5) 
      -- CP-element group 359: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1464_Sample/word_access_start/word_0/$entry
      -- CP-element group 359: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1464_Sample/word_access_start/$entry
      -- CP-element group 359: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1464_Sample/$entry
      -- CP-element group 359: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1464_Sample/word_access_start/word_0/rr
      -- CP-element group 359: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1464_sample_start_
      -- 
    rr_3375_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3375_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(359), ack => ptr_deref_1464_load_0_req_0); -- 
    zeropad3D_A_cp_element_group_359: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_359"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(354) & zeropad3D_A_CP_1983_elements(358) & zeropad3D_A_CP_1983_elements(361);
      gj_zeropad3D_A_cp_element_group_359 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(359), clk => clk, reset => reset); --
    end block;
    -- CP-element group 360:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 360: predecessors 
    -- CP-element group 360: marked-predecessors 
    -- CP-element group 360: 	400 
    -- CP-element group 360: 	362 
    -- CP-element group 360: successors 
    -- CP-element group 360: 	362 
    -- CP-element group 360:  members (5) 
      -- CP-element group 360: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1464_Update/word_access_complete/word_0/$entry
      -- CP-element group 360: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1464_Update/word_access_complete/word_0/cr
      -- CP-element group 360: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1464_Update/word_access_complete/$entry
      -- CP-element group 360: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1464_Update/$entry
      -- CP-element group 360: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1464_update_start_
      -- 
    cr_3386_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3386_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(360), ack => ptr_deref_1464_load_0_req_1); -- 
    zeropad3D_A_cp_element_group_360: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_360"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(400) & zeropad3D_A_CP_1983_elements(362);
      gj_zeropad3D_A_cp_element_group_360 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(360), clk => clk, reset => reset); --
    end block;
    -- CP-element group 361:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 361: predecessors 
    -- CP-element group 361: 	359 
    -- CP-element group 361: successors 
    -- CP-element group 361: marked-successors 
    -- CP-element group 361: 	349 
    -- CP-element group 361: 	356 
    -- CP-element group 361: 	359 
    -- CP-element group 361:  members (5) 
      -- CP-element group 361: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1464_Sample/word_access_start/$exit
      -- CP-element group 361: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1464_Sample/$exit
      -- CP-element group 361: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1464_Sample/word_access_start/word_0/ra
      -- CP-element group 361: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1464_Sample/word_access_start/word_0/$exit
      -- CP-element group 361: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1464_sample_completed_
      -- 
    ra_3376_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 361_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1464_load_0_ack_0, ack => zeropad3D_A_CP_1983_elements(361)); -- 
    -- CP-element group 362:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 362: predecessors 
    -- CP-element group 362: 	360 
    -- CP-element group 362: successors 
    -- CP-element group 362: 	398 
    -- CP-element group 362: marked-successors 
    -- CP-element group 362: 	360 
    -- CP-element group 362:  members (9) 
      -- CP-element group 362: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1464_Update/word_access_complete/word_0/$exit
      -- CP-element group 362: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1464_Update/word_access_complete/word_0/ca
      -- CP-element group 362: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1464_Update/ptr_deref_1464_Merge/merge_ack
      -- CP-element group 362: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1464_Update/word_access_complete/$exit
      -- CP-element group 362: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1464_Update/$exit
      -- CP-element group 362: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1464_Update/ptr_deref_1464_Merge/merge_req
      -- CP-element group 362: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1464_Update/ptr_deref_1464_Merge/$exit
      -- CP-element group 362: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1464_Update/ptr_deref_1464_Merge/$entry
      -- CP-element group 362: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1464_update_completed_
      -- 
    ca_3387_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 362_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1464_load_0_ack_1, ack => zeropad3D_A_CP_1983_elements(362)); -- 
    -- CP-element group 363:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 363: predecessors 
    -- CP-element group 363: 	164 
    -- CP-element group 363: 	172 
    -- CP-element group 363: 	176 
    -- CP-element group 363: 	184 
    -- CP-element group 363: 	188 
    -- CP-element group 363: 	192 
    -- CP-element group 363: 	196 
    -- CP-element group 363: 	200 
    -- CP-element group 363: 	204 
    -- CP-element group 363: 	208 
    -- CP-element group 363: 	212 
    -- CP-element group 363: 	216 
    -- CP-element group 363: 	220 
    -- CP-element group 363: marked-predecessors 
    -- CP-element group 363: 	365 
    -- CP-element group 363: successors 
    -- CP-element group 363: 	365 
    -- CP-element group 363:  members (3) 
      -- CP-element group 363: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1468_sample_start_
      -- CP-element group 363: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1468_Sample/req
      -- CP-element group 363: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1468_Sample/$entry
      -- 
    req_3400_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3400_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(363), ack => W_add96_1324_delayed_2_0_1466_inst_req_0); -- 
    zeropad3D_A_cp_element_group_363: block -- 
      constant place_capacities: IntegerArray(0 to 13) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1);
      constant place_markings: IntegerArray(0 to 13)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 1);
      constant place_delays: IntegerArray(0 to 13) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_363"; 
      signal preds: BooleanArray(1 to 14); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(164) & zeropad3D_A_CP_1983_elements(172) & zeropad3D_A_CP_1983_elements(176) & zeropad3D_A_CP_1983_elements(184) & zeropad3D_A_CP_1983_elements(188) & zeropad3D_A_CP_1983_elements(192) & zeropad3D_A_CP_1983_elements(196) & zeropad3D_A_CP_1983_elements(200) & zeropad3D_A_CP_1983_elements(204) & zeropad3D_A_CP_1983_elements(208) & zeropad3D_A_CP_1983_elements(212) & zeropad3D_A_CP_1983_elements(216) & zeropad3D_A_CP_1983_elements(220) & zeropad3D_A_CP_1983_elements(365);
      gj_zeropad3D_A_cp_element_group_363 : generic_join generic map(name => joinName, number_of_predecessors => 14, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(363), clk => clk, reset => reset); --
    end block;
    -- CP-element group 364:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 364: predecessors 
    -- CP-element group 364: marked-predecessors 
    -- CP-element group 364: 	366 
    -- CP-element group 364: 	369 
    -- CP-element group 364: successors 
    -- CP-element group 364: 	366 
    -- CP-element group 364:  members (3) 
      -- CP-element group 364: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1468_update_start_
      -- CP-element group 364: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1468_Update/req
      -- CP-element group 364: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1468_Update/$entry
      -- 
    req_3405_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3405_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(364), ack => W_add96_1324_delayed_2_0_1466_inst_req_1); -- 
    zeropad3D_A_cp_element_group_364: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_364"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(366) & zeropad3D_A_CP_1983_elements(369);
      gj_zeropad3D_A_cp_element_group_364 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(364), clk => clk, reset => reset); --
    end block;
    -- CP-element group 365:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 365: predecessors 
    -- CP-element group 365: 	363 
    -- CP-element group 365: successors 
    -- CP-element group 365: marked-successors 
    -- CP-element group 365: 	162 
    -- CP-element group 365: 	170 
    -- CP-element group 365: 	174 
    -- CP-element group 365: 	182 
    -- CP-element group 365: 	186 
    -- CP-element group 365: 	190 
    -- CP-element group 365: 	194 
    -- CP-element group 365: 	198 
    -- CP-element group 365: 	202 
    -- CP-element group 365: 	206 
    -- CP-element group 365: 	210 
    -- CP-element group 365: 	214 
    -- CP-element group 365: 	218 
    -- CP-element group 365: 	363 
    -- CP-element group 365:  members (3) 
      -- CP-element group 365: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1468_sample_completed_
      -- CP-element group 365: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1468_Sample/$exit
      -- CP-element group 365: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1468_Sample/ack
      -- 
    ack_3401_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 365_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_add96_1324_delayed_2_0_1466_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(365)); -- 
    -- CP-element group 366:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 366: predecessors 
    -- CP-element group 366: 	364 
    -- CP-element group 366: successors 
    -- CP-element group 366: 	367 
    -- CP-element group 366: marked-successors 
    -- CP-element group 366: 	364 
    -- CP-element group 366:  members (3) 
      -- CP-element group 366: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1468_update_completed_
      -- CP-element group 366: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1468_Update/ack
      -- CP-element group 366: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1468_Update/$exit
      -- 
    ack_3406_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 366_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_add96_1324_delayed_2_0_1466_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(366)); -- 
    -- CP-element group 367:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 367: predecessors 
    -- CP-element group 367: 	264 
    -- CP-element group 367: 	280 
    -- CP-element group 367: 	288 
    -- CP-element group 367: 	366 
    -- CP-element group 367: marked-predecessors 
    -- CP-element group 367: 	369 
    -- CP-element group 367: successors 
    -- CP-element group 367: 	369 
    -- CP-element group 367:  members (3) 
      -- CP-element group 367: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1473_Sample/rr
      -- CP-element group 367: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1473_Sample/$entry
      -- CP-element group 367: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1473_sample_start_
      -- 
    rr_3414_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3414_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(367), ack => type_cast_1473_inst_req_0); -- 
    zeropad3D_A_cp_element_group_367: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_367"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(264) & zeropad3D_A_CP_1983_elements(280) & zeropad3D_A_CP_1983_elements(288) & zeropad3D_A_CP_1983_elements(366) & zeropad3D_A_CP_1983_elements(369);
      gj_zeropad3D_A_cp_element_group_367 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(367), clk => clk, reset => reset); --
    end block;
    -- CP-element group 368:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 368: predecessors 
    -- CP-element group 368: marked-predecessors 
    -- CP-element group 368: 	381 
    -- CP-element group 368: 	370 
    -- CP-element group 368: successors 
    -- CP-element group 368: 	370 
    -- CP-element group 368:  members (3) 
      -- CP-element group 368: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1473_Update/cr
      -- CP-element group 368: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1473_Update/$entry
      -- CP-element group 368: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1473_update_start_
      -- 
    cr_3419_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3419_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(368), ack => type_cast_1473_inst_req_1); -- 
    zeropad3D_A_cp_element_group_368: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_368"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(381) & zeropad3D_A_CP_1983_elements(370);
      gj_zeropad3D_A_cp_element_group_368 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(368), clk => clk, reset => reset); --
    end block;
    -- CP-element group 369:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 369: predecessors 
    -- CP-element group 369: 	367 
    -- CP-element group 369: successors 
    -- CP-element group 369: marked-successors 
    -- CP-element group 369: 	262 
    -- CP-element group 369: 	278 
    -- CP-element group 369: 	286 
    -- CP-element group 369: 	364 
    -- CP-element group 369: 	367 
    -- CP-element group 369:  members (3) 
      -- CP-element group 369: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1473_Sample/ra
      -- CP-element group 369: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1473_Sample/$exit
      -- CP-element group 369: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1473_sample_completed_
      -- 
    ra_3415_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 369_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1473_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(369)); -- 
    -- CP-element group 370:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 370: predecessors 
    -- CP-element group 370: 	368 
    -- CP-element group 370: successors 
    -- CP-element group 370: 	379 
    -- CP-element group 370: marked-successors 
    -- CP-element group 370: 	368 
    -- CP-element group 370:  members (3) 
      -- CP-element group 370: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1473_Update/ca
      -- CP-element group 370: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1473_Update/$exit
      -- CP-element group 370: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1473_update_completed_
      -- 
    ca_3420_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 370_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1473_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(370)); -- 
    -- CP-element group 371:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 371: predecessors 
    -- CP-element group 371: 	264 
    -- CP-element group 371: 	280 
    -- CP-element group 371: 	288 
    -- CP-element group 371: marked-predecessors 
    -- CP-element group 371: 	373 
    -- CP-element group 371: successors 
    -- CP-element group 371: 	373 
    -- CP-element group 371:  members (3) 
      -- CP-element group 371: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1477_Sample/req
      -- CP-element group 371: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1477_Sample/$entry
      -- CP-element group 371: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1477_sample_start_
      -- 
    req_3428_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3428_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(371), ack => W_ifx_xelse155_exec_guard_1328_delayed_1_0_1475_inst_req_0); -- 
    zeropad3D_A_cp_element_group_371: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_371"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(264) & zeropad3D_A_CP_1983_elements(280) & zeropad3D_A_CP_1983_elements(288) & zeropad3D_A_CP_1983_elements(373);
      gj_zeropad3D_A_cp_element_group_371 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(371), clk => clk, reset => reset); --
    end block;
    -- CP-element group 372:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 372: predecessors 
    -- CP-element group 372: marked-predecessors 
    -- CP-element group 372: 	374 
    -- CP-element group 372: successors 
    -- CP-element group 372: 	374 
    -- CP-element group 372:  members (3) 
      -- CP-element group 372: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1477_Update/req
      -- CP-element group 372: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1477_Update/$entry
      -- CP-element group 372: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1477_update_start_
      -- 
    req_3433_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3433_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(372), ack => W_ifx_xelse155_exec_guard_1328_delayed_1_0_1475_inst_req_1); -- 
    zeropad3D_A_cp_element_group_372: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_372"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= zeropad3D_A_CP_1983_elements(374);
      gj_zeropad3D_A_cp_element_group_372 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(372), clk => clk, reset => reset); --
    end block;
    -- CP-element group 373:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 373: predecessors 
    -- CP-element group 373: 	371 
    -- CP-element group 373: successors 
    -- CP-element group 373: marked-successors 
    -- CP-element group 373: 	262 
    -- CP-element group 373: 	278 
    -- CP-element group 373: 	286 
    -- CP-element group 373: 	371 
    -- CP-element group 373:  members (3) 
      -- CP-element group 373: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1477_Sample/ack
      -- CP-element group 373: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1477_Sample/$exit
      -- CP-element group 373: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1477_sample_completed_
      -- 
    ack_3429_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 373_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xelse155_exec_guard_1328_delayed_1_0_1475_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(373)); -- 
    -- CP-element group 374:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 374: predecessors 
    -- CP-element group 374: 	372 
    -- CP-element group 374: successors 
    -- CP-element group 374: 	404 
    -- CP-element group 374: marked-successors 
    -- CP-element group 374: 	372 
    -- CP-element group 374:  members (3) 
      -- CP-element group 374: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1477_Update/ack
      -- CP-element group 374: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1477_Update/$exit
      -- CP-element group 374: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1477_update_completed_
      -- 
    ack_3434_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 374_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xelse155_exec_guard_1328_delayed_1_0_1475_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(374)); -- 
    -- CP-element group 375:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 375: predecessors 
    -- CP-element group 375: 	264 
    -- CP-element group 375: 	280 
    -- CP-element group 375: 	288 
    -- CP-element group 375: marked-predecessors 
    -- CP-element group 375: 	377 
    -- CP-element group 375: successors 
    -- CP-element group 375: 	377 
    -- CP-element group 375:  members (3) 
      -- CP-element group 375: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1490_sample_start_
      -- CP-element group 375: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1490_Sample/$entry
      -- CP-element group 375: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1490_Sample/req
      -- 
    req_3442_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3442_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(375), ack => W_ifx_xelse155_exec_guard_1338_delayed_1_0_1488_inst_req_0); -- 
    zeropad3D_A_cp_element_group_375: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_375"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(264) & zeropad3D_A_CP_1983_elements(280) & zeropad3D_A_CP_1983_elements(288) & zeropad3D_A_CP_1983_elements(377);
      gj_zeropad3D_A_cp_element_group_375 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(375), clk => clk, reset => reset); --
    end block;
    -- CP-element group 376:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 376: predecessors 
    -- CP-element group 376: marked-predecessors 
    -- CP-element group 376: 	381 
    -- CP-element group 376: 	378 
    -- CP-element group 376: successors 
    -- CP-element group 376: 	378 
    -- CP-element group 376:  members (3) 
      -- CP-element group 376: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1490_update_start_
      -- CP-element group 376: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1490_Update/req
      -- CP-element group 376: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1490_Update/$entry
      -- 
    req_3447_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3447_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(376), ack => W_ifx_xelse155_exec_guard_1338_delayed_1_0_1488_inst_req_1); -- 
    zeropad3D_A_cp_element_group_376: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_376"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(381) & zeropad3D_A_CP_1983_elements(378);
      gj_zeropad3D_A_cp_element_group_376 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(376), clk => clk, reset => reset); --
    end block;
    -- CP-element group 377:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 377: predecessors 
    -- CP-element group 377: 	375 
    -- CP-element group 377: successors 
    -- CP-element group 377: marked-successors 
    -- CP-element group 377: 	262 
    -- CP-element group 377: 	278 
    -- CP-element group 377: 	286 
    -- CP-element group 377: 	375 
    -- CP-element group 377:  members (3) 
      -- CP-element group 377: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1490_sample_completed_
      -- CP-element group 377: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1490_Sample/$exit
      -- CP-element group 377: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1490_Sample/ack
      -- 
    ack_3443_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 377_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xelse155_exec_guard_1338_delayed_1_0_1488_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(377)); -- 
    -- CP-element group 378:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 378: predecessors 
    -- CP-element group 378: 	376 
    -- CP-element group 378: successors 
    -- CP-element group 378: 	379 
    -- CP-element group 378: marked-successors 
    -- CP-element group 378: 	376 
    -- CP-element group 378:  members (3) 
      -- CP-element group 378: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1490_update_completed_
      -- CP-element group 378: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1490_Update/ack
      -- CP-element group 378: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1490_Update/$exit
      -- 
    ack_3448_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 378_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xelse155_exec_guard_1338_delayed_1_0_1488_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(378)); -- 
    -- CP-element group 379:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 379: predecessors 
    -- CP-element group 379: 	370 
    -- CP-element group 379: 	378 
    -- CP-element group 379: marked-predecessors 
    -- CP-element group 379: 	381 
    -- CP-element group 379: successors 
    -- CP-element group 379: 	381 
    -- CP-element group 379:  members (3) 
      -- CP-element group 379: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1495_Sample/$entry
      -- CP-element group 379: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1495_Sample/rr
      -- CP-element group 379: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1495_sample_start_
      -- 
    rr_3456_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3456_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(379), ack => type_cast_1495_inst_req_0); -- 
    zeropad3D_A_cp_element_group_379: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_379"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(370) & zeropad3D_A_CP_1983_elements(378) & zeropad3D_A_CP_1983_elements(381);
      gj_zeropad3D_A_cp_element_group_379 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(379), clk => clk, reset => reset); --
    end block;
    -- CP-element group 380:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 380: predecessors 
    -- CP-element group 380: marked-predecessors 
    -- CP-element group 380: 	382 
    -- CP-element group 380: 	386 
    -- CP-element group 380: successors 
    -- CP-element group 380: 	382 
    -- CP-element group 380:  members (3) 
      -- CP-element group 380: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1495_Update/$entry
      -- CP-element group 380: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1495_update_start_
      -- CP-element group 380: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1495_Update/cr
      -- 
    cr_3461_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3461_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(380), ack => type_cast_1495_inst_req_1); -- 
    zeropad3D_A_cp_element_group_380: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_380"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(382) & zeropad3D_A_CP_1983_elements(386);
      gj_zeropad3D_A_cp_element_group_380 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(380), clk => clk, reset => reset); --
    end block;
    -- CP-element group 381:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 381: predecessors 
    -- CP-element group 381: 	379 
    -- CP-element group 381: successors 
    -- CP-element group 381: marked-successors 
    -- CP-element group 381: 	368 
    -- CP-element group 381: 	376 
    -- CP-element group 381: 	379 
    -- CP-element group 381:  members (3) 
      -- CP-element group 381: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1495_Sample/ra
      -- CP-element group 381: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1495_Sample/$exit
      -- CP-element group 381: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1495_sample_completed_
      -- 
    ra_3457_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 381_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1495_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(381)); -- 
    -- CP-element group 382:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 382: predecessors 
    -- CP-element group 382: 	380 
    -- CP-element group 382: successors 
    -- CP-element group 382: 	386 
    -- CP-element group 382: marked-successors 
    -- CP-element group 382: 	380 
    -- CP-element group 382:  members (16) 
      -- CP-element group 382: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1495_update_completed_
      -- CP-element group 382: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1501_final_index_sum_regn_Sample/req
      -- CP-element group 382: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1501_final_index_sum_regn_Sample/$entry
      -- CP-element group 382: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1501_index_scale_1/scale_rename_ack
      -- CP-element group 382: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1501_index_scale_1/scale_rename_req
      -- CP-element group 382: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1501_index_scale_1/$exit
      -- CP-element group 382: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1501_index_scale_1/$entry
      -- CP-element group 382: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1501_index_resize_1/index_resize_ack
      -- CP-element group 382: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1501_index_resize_1/index_resize_req
      -- CP-element group 382: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1501_index_resize_1/$exit
      -- CP-element group 382: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1501_index_resize_1/$entry
      -- CP-element group 382: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1501_index_computed_1
      -- CP-element group 382: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1501_index_scaled_1
      -- CP-element group 382: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1501_index_resized_1
      -- CP-element group 382: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1495_Update/ca
      -- CP-element group 382: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/type_cast_1495_Update/$exit
      -- 
    ca_3462_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 382_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1495_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(382)); -- 
    req_3487_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3487_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(382), ack => array_obj_ref_1501_index_offset_req_0); -- 
    -- CP-element group 383:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 383: predecessors 
    -- CP-element group 383: 	387 
    -- CP-element group 383: marked-predecessors 
    -- CP-element group 383: 	388 
    -- CP-element group 383: successors 
    -- CP-element group 383: 	388 
    -- CP-element group 383:  members (3) 
      -- CP-element group 383: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/addr_of_1502_request/req
      -- CP-element group 383: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/addr_of_1502_request/$entry
      -- CP-element group 383: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/addr_of_1502_sample_start_
      -- 
    req_3502_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3502_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(383), ack => addr_of_1502_final_reg_req_0); -- 
    zeropad3D_A_cp_element_group_383: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_383"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(387) & zeropad3D_A_CP_1983_elements(388);
      gj_zeropad3D_A_cp_element_group_383 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(383), clk => clk, reset => reset); --
    end block;
    -- CP-element group 384:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 384: predecessors 
    -- CP-element group 384: 	42 
    -- CP-element group 384: marked-predecessors 
    -- CP-element group 384: 	389 
    -- CP-element group 384: 	396 
    -- CP-element group 384: successors 
    -- CP-element group 384: 	389 
    -- CP-element group 384:  members (3) 
      -- CP-element group 384: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/addr_of_1502_complete/$entry
      -- CP-element group 384: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/addr_of_1502_complete/req
      -- CP-element group 384: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/addr_of_1502_update_start_
      -- 
    req_3507_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3507_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(384), ack => addr_of_1502_final_reg_req_1); -- 
    zeropad3D_A_cp_element_group_384: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_384"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(42) & zeropad3D_A_CP_1983_elements(389) & zeropad3D_A_CP_1983_elements(396);
      gj_zeropad3D_A_cp_element_group_384 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(384), clk => clk, reset => reset); --
    end block;
    -- CP-element group 385:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 385: predecessors 
    -- CP-element group 385: 	42 
    -- CP-element group 385: marked-predecessors 
    -- CP-element group 385: 	387 
    -- CP-element group 385: 	388 
    -- CP-element group 385: successors 
    -- CP-element group 385: 	387 
    -- CP-element group 385:  members (3) 
      -- CP-element group 385: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1501_final_index_sum_regn_Update/req
      -- CP-element group 385: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1501_final_index_sum_regn_Update/$entry
      -- CP-element group 385: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1501_final_index_sum_regn_update_start
      -- 
    req_3492_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3492_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(385), ack => array_obj_ref_1501_index_offset_req_1); -- 
    zeropad3D_A_cp_element_group_385: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_385"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(42) & zeropad3D_A_CP_1983_elements(387) & zeropad3D_A_CP_1983_elements(388);
      gj_zeropad3D_A_cp_element_group_385 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(385), clk => clk, reset => reset); --
    end block;
    -- CP-element group 386:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 386: predecessors 
    -- CP-element group 386: 	382 
    -- CP-element group 386: successors 
    -- CP-element group 386: 	404 
    -- CP-element group 386: marked-successors 
    -- CP-element group 386: 	380 
    -- CP-element group 386:  members (3) 
      -- CP-element group 386: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1501_final_index_sum_regn_Sample/ack
      -- CP-element group 386: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1501_final_index_sum_regn_Sample/$exit
      -- CP-element group 386: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1501_final_index_sum_regn_sample_complete
      -- 
    ack_3488_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 386_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1501_index_offset_ack_0, ack => zeropad3D_A_CP_1983_elements(386)); -- 
    -- CP-element group 387:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 387: predecessors 
    -- CP-element group 387: 	385 
    -- CP-element group 387: successors 
    -- CP-element group 387: 	383 
    -- CP-element group 387: marked-successors 
    -- CP-element group 387: 	385 
    -- CP-element group 387:  members (8) 
      -- CP-element group 387: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1501_base_plus_offset/sum_rename_ack
      -- CP-element group 387: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1501_base_plus_offset/sum_rename_req
      -- CP-element group 387: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1501_base_plus_offset/$exit
      -- CP-element group 387: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1501_base_plus_offset/$entry
      -- CP-element group 387: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1501_final_index_sum_regn_Update/ack
      -- CP-element group 387: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1501_final_index_sum_regn_Update/$exit
      -- CP-element group 387: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1501_offset_calculated
      -- CP-element group 387: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/array_obj_ref_1501_root_address_calculated
      -- 
    ack_3493_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 387_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1501_index_offset_ack_1, ack => zeropad3D_A_CP_1983_elements(387)); -- 
    -- CP-element group 388:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 388: predecessors 
    -- CP-element group 388: 	383 
    -- CP-element group 388: successors 
    -- CP-element group 388: marked-successors 
    -- CP-element group 388: 	383 
    -- CP-element group 388: 	385 
    -- CP-element group 388:  members (3) 
      -- CP-element group 388: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/addr_of_1502_request/ack
      -- CP-element group 388: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/addr_of_1502_request/$exit
      -- CP-element group 388: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/addr_of_1502_sample_completed_
      -- 
    ack_3503_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 388_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1502_final_reg_ack_0, ack => zeropad3D_A_CP_1983_elements(388)); -- 
    -- CP-element group 389:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 389: predecessors 
    -- CP-element group 389: 	384 
    -- CP-element group 389: successors 
    -- CP-element group 389: 	394 
    -- CP-element group 389: marked-successors 
    -- CP-element group 389: 	384 
    -- CP-element group 389:  members (3) 
      -- CP-element group 389: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/addr_of_1502_complete/$exit
      -- CP-element group 389: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/addr_of_1502_complete/ack
      -- CP-element group 389: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/addr_of_1502_update_completed_
      -- 
    ack_3508_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 389_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1502_final_reg_ack_1, ack => zeropad3D_A_CP_1983_elements(389)); -- 
    -- CP-element group 390:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 390: predecessors 
    -- CP-element group 390: 	264 
    -- CP-element group 390: 	280 
    -- CP-element group 390: 	288 
    -- CP-element group 390: marked-predecessors 
    -- CP-element group 390: 	392 
    -- CP-element group 390: successors 
    -- CP-element group 390: 	392 
    -- CP-element group 390:  members (3) 
      -- CP-element group 390: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1506_sample_start_
      -- CP-element group 390: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1506_Sample/$entry
      -- CP-element group 390: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1506_Sample/req
      -- 
    req_3516_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3516_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(390), ack => W_ifx_xelse155_exec_guard_1351_delayed_15_0_1504_inst_req_0); -- 
    zeropad3D_A_cp_element_group_390: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_390"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(264) & zeropad3D_A_CP_1983_elements(280) & zeropad3D_A_CP_1983_elements(288) & zeropad3D_A_CP_1983_elements(392);
      gj_zeropad3D_A_cp_element_group_390 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(390), clk => clk, reset => reset); --
    end block;
    -- CP-element group 391:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 391: predecessors 
    -- CP-element group 391: marked-predecessors 
    -- CP-element group 391: 	393 
    -- CP-element group 391: successors 
    -- CP-element group 391: 	393 
    -- CP-element group 391:  members (3) 
      -- CP-element group 391: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1506_update_start_
      -- CP-element group 391: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1506_Update/req
      -- CP-element group 391: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1506_Update/$entry
      -- 
    req_3521_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3521_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(391), ack => W_ifx_xelse155_exec_guard_1351_delayed_15_0_1504_inst_req_1); -- 
    zeropad3D_A_cp_element_group_391: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_391"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= zeropad3D_A_CP_1983_elements(393);
      gj_zeropad3D_A_cp_element_group_391 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(391), clk => clk, reset => reset); --
    end block;
    -- CP-element group 392:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 392: predecessors 
    -- CP-element group 392: 	390 
    -- CP-element group 392: successors 
    -- CP-element group 392: marked-successors 
    -- CP-element group 392: 	390 
    -- CP-element group 392: 	262 
    -- CP-element group 392: 	278 
    -- CP-element group 392: 	286 
    -- CP-element group 392:  members (3) 
      -- CP-element group 392: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1506_sample_completed_
      -- CP-element group 392: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1506_Sample/ack
      -- CP-element group 392: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1506_Sample/$exit
      -- 
    ack_3517_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 392_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xelse155_exec_guard_1351_delayed_15_0_1504_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(392)); -- 
    -- CP-element group 393:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 393: predecessors 
    -- CP-element group 393: 	391 
    -- CP-element group 393: successors 
    -- CP-element group 393: 	404 
    -- CP-element group 393: marked-successors 
    -- CP-element group 393: 	391 
    -- CP-element group 393:  members (3) 
      -- CP-element group 393: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1506_update_completed_
      -- CP-element group 393: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1506_Update/ack
      -- CP-element group 393: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1506_Update/$exit
      -- 
    ack_3522_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 393_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_ifx_xelse155_exec_guard_1351_delayed_15_0_1504_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(393)); -- 
    -- CP-element group 394:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 394: predecessors 
    -- CP-element group 394: 	389 
    -- CP-element group 394: marked-predecessors 
    -- CP-element group 394: 	396 
    -- CP-element group 394: successors 
    -- CP-element group 394: 	396 
    -- CP-element group 394:  members (3) 
      -- CP-element group 394: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1509_Sample/req
      -- CP-element group 394: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1509_Sample/$entry
      -- CP-element group 394: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1509_sample_start_
      -- 
    req_3530_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3530_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(394), ack => W_arrayidx166_1352_delayed_6_0_1507_inst_req_0); -- 
    zeropad3D_A_cp_element_group_394: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_394"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(389) & zeropad3D_A_CP_1983_elements(396);
      gj_zeropad3D_A_cp_element_group_394 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(394), clk => clk, reset => reset); --
    end block;
    -- CP-element group 395:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 395: predecessors 
    -- CP-element group 395: marked-predecessors 
    -- CP-element group 395: 	400 
    -- CP-element group 395: 	397 
    -- CP-element group 395: successors 
    -- CP-element group 395: 	397 
    -- CP-element group 395:  members (3) 
      -- CP-element group 395: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1509_Update/req
      -- CP-element group 395: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1509_Update/$entry
      -- CP-element group 395: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1509_update_start_
      -- 
    req_3535_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3535_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(395), ack => W_arrayidx166_1352_delayed_6_0_1507_inst_req_1); -- 
    zeropad3D_A_cp_element_group_395: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_395"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(400) & zeropad3D_A_CP_1983_elements(397);
      gj_zeropad3D_A_cp_element_group_395 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(395), clk => clk, reset => reset); --
    end block;
    -- CP-element group 396:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 396: predecessors 
    -- CP-element group 396: 	394 
    -- CP-element group 396: successors 
    -- CP-element group 396: marked-successors 
    -- CP-element group 396: 	384 
    -- CP-element group 396: 	394 
    -- CP-element group 396:  members (3) 
      -- CP-element group 396: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1509_Sample/ack
      -- CP-element group 396: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1509_Sample/$exit
      -- CP-element group 396: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1509_sample_completed_
      -- 
    ack_3531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 396_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_arrayidx166_1352_delayed_6_0_1507_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(396)); -- 
    -- CP-element group 397:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 397: predecessors 
    -- CP-element group 397: 	395 
    -- CP-element group 397: successors 
    -- CP-element group 397: 	398 
    -- CP-element group 397: marked-successors 
    -- CP-element group 397: 	395 
    -- CP-element group 397:  members (19) 
      -- CP-element group 397: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1512_word_addrgen/$entry
      -- CP-element group 397: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1512_word_addrgen/root_register_req
      -- CP-element group 397: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1512_word_addrgen/$exit
      -- CP-element group 397: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1512_base_plus_offset/sum_rename_req
      -- CP-element group 397: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1512_base_plus_offset/$entry
      -- CP-element group 397: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1512_word_addrgen/root_register_ack
      -- CP-element group 397: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1512_base_plus_offset/sum_rename_ack
      -- CP-element group 397: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1512_base_plus_offset/$exit
      -- CP-element group 397: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1512_base_addr_resize/base_resize_ack
      -- CP-element group 397: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1512_base_addr_resize/base_resize_req
      -- CP-element group 397: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1512_base_addr_resize/$exit
      -- CP-element group 397: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1512_base_addr_resize/$entry
      -- CP-element group 397: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1512_base_address_resized
      -- CP-element group 397: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1512_root_address_calculated
      -- CP-element group 397: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1512_word_address_calculated
      -- CP-element group 397: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1512_base_address_calculated
      -- CP-element group 397: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1509_Update/ack
      -- CP-element group 397: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1509_Update/$exit
      -- CP-element group 397: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/assign_stmt_1509_update_completed_
      -- 
    ack_3536_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 397_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_arrayidx166_1352_delayed_6_0_1507_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(397)); -- 
    -- CP-element group 398:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 398: predecessors 
    -- CP-element group 398: 	403 
    -- CP-element group 398: 	397 
    -- CP-element group 398: 	362 
    -- CP-element group 398: marked-predecessors 
    -- CP-element group 398: 	400 
    -- CP-element group 398: successors 
    -- CP-element group 398: 	400 
    -- CP-element group 398:  members (9) 
      -- CP-element group 398: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1512_Sample/ptr_deref_1512_Split/split_ack
      -- CP-element group 398: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1512_Sample/$entry
      -- CP-element group 398: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1512_Sample/word_access_start/$entry
      -- CP-element group 398: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1512_Sample/ptr_deref_1512_Split/$entry
      -- CP-element group 398: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1512_Sample/ptr_deref_1512_Split/$exit
      -- CP-element group 398: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1512_Sample/ptr_deref_1512_Split/split_req
      -- CP-element group 398: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1512_Sample/word_access_start/word_0/$entry
      -- CP-element group 398: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1512_sample_start_
      -- CP-element group 398: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1512_Sample/word_access_start/word_0/rr
      -- 
    rr_3574_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3574_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(398), ack => ptr_deref_1512_store_0_req_0); -- 
    zeropad3D_A_cp_element_group_398: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_398"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(403) & zeropad3D_A_CP_1983_elements(397) & zeropad3D_A_CP_1983_elements(362) & zeropad3D_A_CP_1983_elements(400);
      gj_zeropad3D_A_cp_element_group_398 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(398), clk => clk, reset => reset); --
    end block;
    -- CP-element group 399:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 399: predecessors 
    -- CP-element group 399: marked-predecessors 
    -- CP-element group 399: 	401 
    -- CP-element group 399: successors 
    -- CP-element group 399: 	401 
    -- CP-element group 399:  members (5) 
      -- CP-element group 399: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1512_Update/word_access_complete/word_0/$entry
      -- CP-element group 399: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1512_Update/word_access_complete/word_0/cr
      -- CP-element group 399: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1512_Update/word_access_complete/$entry
      -- CP-element group 399: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1512_Update/$entry
      -- CP-element group 399: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1512_update_start_
      -- 
    cr_3585_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3585_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(399), ack => ptr_deref_1512_store_0_req_1); -- 
    zeropad3D_A_cp_element_group_399: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_399"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= zeropad3D_A_CP_1983_elements(401);
      gj_zeropad3D_A_cp_element_group_399 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(399), clk => clk, reset => reset); --
    end block;
    -- CP-element group 400:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 400: predecessors 
    -- CP-element group 400: 	398 
    -- CP-element group 400: successors 
    -- CP-element group 400: 	404 
    -- CP-element group 400: marked-successors 
    -- CP-element group 400: 	395 
    -- CP-element group 400: 	398 
    -- CP-element group 400: 	324 
    -- CP-element group 400: 	360 
    -- CP-element group 400:  members (6) 
      -- CP-element group 400: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1512_Sample/word_access_start/word_0/ra
      -- CP-element group 400: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1512_Sample/$exit
      -- CP-element group 400: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1512_Sample/word_access_start/$exit
      -- CP-element group 400: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1512_sample_completed_
      -- CP-element group 400: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ring_reenable_memory_space_0
      -- CP-element group 400: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1512_Sample/word_access_start/word_0/$exit
      -- 
    ra_3575_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 400_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1512_store_0_ack_0, ack => zeropad3D_A_CP_1983_elements(400)); -- 
    -- CP-element group 401:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 401: predecessors 
    -- CP-element group 401: 	399 
    -- CP-element group 401: successors 
    -- CP-element group 401: 	404 
    -- CP-element group 401: marked-successors 
    -- CP-element group 401: 	399 
    -- CP-element group 401:  members (5) 
      -- CP-element group 401: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1512_Update/word_access_complete/word_0/$exit
      -- CP-element group 401: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1512_Update/$exit
      -- CP-element group 401: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1512_Update/word_access_complete/$exit
      -- CP-element group 401: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1512_Update/word_access_complete/word_0/ca
      -- CP-element group 401: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1512_update_completed_
      -- 
    ca_3586_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 401_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1512_store_0_ack_1, ack => zeropad3D_A_CP_1983_elements(401)); -- 
    -- CP-element group 402:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 402: predecessors 
    -- CP-element group 402: 	42 
    -- CP-element group 402: successors 
    -- CP-element group 402: 	43 
    -- CP-element group 402:  members (1) 
      -- CP-element group 402: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group zeropad3D_A_CP_1983_elements(402) is a control-delay.
    cp_element_402_delay: control_delay_element  generic map(name => " 402_delay", delay_value => 1)  port map(req => zeropad3D_A_CP_1983_elements(42), ack => zeropad3D_A_CP_1983_elements(402), clk => clk, reset =>reset);
    -- CP-element group 403:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 403: predecessors 
    -- CP-element group 403: 	326 
    -- CP-element group 403: successors 
    -- CP-element group 403: 	398 
    -- CP-element group 403:  members (1) 
      -- CP-element group 403: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/ptr_deref_1413_ptr_deref_1512_delay
      -- 
    -- Element group zeropad3D_A_CP_1983_elements(403) is a control-delay.
    cp_element_403_delay: control_delay_element  generic map(name => " 403_delay", delay_value => 1)  port map(req => zeropad3D_A_CP_1983_elements(326), ack => zeropad3D_A_CP_1983_elements(403), clk => clk, reset =>reset);
    -- CP-element group 404:  join  transition  bypass  pipeline-parent 
    -- CP-element group 404: predecessors 
    -- CP-element group 404: 	400 
    -- CP-element group 404: 	401 
    -- CP-element group 404: 	386 
    -- CP-element group 404: 	393 
    -- CP-element group 404: 	132 
    -- CP-element group 404: 	144 
    -- CP-element group 404: 	152 
    -- CP-element group 404: 	168 
    -- CP-element group 404: 	232 
    -- CP-element group 404: 	236 
    -- CP-element group 404: 	240 
    -- CP-element group 404: 	248 
    -- CP-element group 404: 	268 
    -- CP-element group 404: 	272 
    -- CP-element group 404: 	276 
    -- CP-element group 404: 	284 
    -- CP-element group 404: 	308 
    -- CP-element group 404: 	320 
    -- CP-element group 404: 	327 
    -- CP-element group 404: 	339 
    -- CP-element group 404: 	351 
    -- CP-element group 404: 	374 
    -- CP-element group 404: successors 
    -- CP-element group 404: 	39 
    -- CP-element group 404:  members (1) 
      -- CP-element group 404: 	 branch_block_stmt_783/do_while_stmt_903/do_while_stmt_903_loop_body/$exit
      -- 
    zeropad3D_A_cp_element_group_404: block -- 
      constant place_capacities: IntegerArray(0 to 21) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 15,8 => 15,9 => 15,10 => 15,11 => 15,12 => 15,13 => 15,14 => 15,15 => 15,16 => 15,17 => 15,18 => 15,19 => 15,20 => 15,21 => 15);
      constant place_markings: IntegerArray(0 to 21)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0,21 => 0);
      constant place_delays: IntegerArray(0 to 21) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0,21 => 0);
      constant joinName: string(1 to 32) := "zeropad3D_A_cp_element_group_404"; 
      signal preds: BooleanArray(1 to 22); -- 
    begin -- 
      preds <= zeropad3D_A_CP_1983_elements(400) & zeropad3D_A_CP_1983_elements(401) & zeropad3D_A_CP_1983_elements(386) & zeropad3D_A_CP_1983_elements(393) & zeropad3D_A_CP_1983_elements(132) & zeropad3D_A_CP_1983_elements(144) & zeropad3D_A_CP_1983_elements(152) & zeropad3D_A_CP_1983_elements(168) & zeropad3D_A_CP_1983_elements(232) & zeropad3D_A_CP_1983_elements(236) & zeropad3D_A_CP_1983_elements(240) & zeropad3D_A_CP_1983_elements(248) & zeropad3D_A_CP_1983_elements(268) & zeropad3D_A_CP_1983_elements(272) & zeropad3D_A_CP_1983_elements(276) & zeropad3D_A_CP_1983_elements(284) & zeropad3D_A_CP_1983_elements(308) & zeropad3D_A_CP_1983_elements(320) & zeropad3D_A_CP_1983_elements(327) & zeropad3D_A_CP_1983_elements(339) & zeropad3D_A_CP_1983_elements(351) & zeropad3D_A_CP_1983_elements(374);
      gj_zeropad3D_A_cp_element_group_404 : generic_join generic map(name => joinName, number_of_predecessors => 22, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(404), clk => clk, reset => reset); --
    end block;
    -- CP-element group 405:  transition  input  bypass  pipeline-parent 
    -- CP-element group 405: predecessors 
    -- CP-element group 405: 	38 
    -- CP-element group 405: successors 
    -- CP-element group 405:  members (2) 
      -- CP-element group 405: 	 branch_block_stmt_783/do_while_stmt_903/loop_exit/ack
      -- CP-element group 405: 	 branch_block_stmt_783/do_while_stmt_903/loop_exit/$exit
      -- 
    ack_3593_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 405_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_903_branch_ack_0, ack => zeropad3D_A_CP_1983_elements(405)); -- 
    -- CP-element group 406:  transition  input  bypass  pipeline-parent 
    -- CP-element group 406: predecessors 
    -- CP-element group 406: 	38 
    -- CP-element group 406: successors 
    -- CP-element group 406:  members (2) 
      -- CP-element group 406: 	 branch_block_stmt_783/do_while_stmt_903/loop_taken/ack
      -- CP-element group 406: 	 branch_block_stmt_783/do_while_stmt_903/loop_taken/$exit
      -- 
    ack_3597_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 406_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_903_branch_ack_1, ack => zeropad3D_A_CP_1983_elements(406)); -- 
    -- CP-element group 407:  transition  bypass  pipeline-parent 
    -- CP-element group 407: predecessors 
    -- CP-element group 407: 	36 
    -- CP-element group 407: successors 
    -- CP-element group 407: 	1 
    -- CP-element group 407:  members (1) 
      -- CP-element group 407: 	 branch_block_stmt_783/do_while_stmt_903/$exit
      -- 
    zeropad3D_A_CP_1983_elements(407) <= zeropad3D_A_CP_1983_elements(36);
    -- CP-element group 408:  merge  transition  place  input  output  bypass 
    -- CP-element group 408: predecessors 
    -- CP-element group 408: 	1 
    -- CP-element group 408: successors 
    -- CP-element group 408: 	410 
    -- CP-element group 408:  members (15) 
      -- CP-element group 408: 	 branch_block_stmt_783/merge_stmt_1531_PhiReqMerge
      -- CP-element group 408: 	 branch_block_stmt_783/merge_stmt_1531__exit__
      -- CP-element group 408: 	 branch_block_stmt_783/assign_stmt_1536__entry__
      -- CP-element group 408: 	 branch_block_stmt_783/assign_stmt_1536/$entry
      -- CP-element group 408: 	 branch_block_stmt_783/if_stmt_1527_if_link/if_choice_transition
      -- CP-element group 408: 	 branch_block_stmt_783/if_stmt_1527_if_link/$exit
      -- CP-element group 408: 	 branch_block_stmt_783/assign_stmt_1536/WPIPE_Block0_complete_1533_sample_start_
      -- CP-element group 408: 	 branch_block_stmt_783/merge_stmt_1531_PhiAck/dummy
      -- CP-element group 408: 	 branch_block_stmt_783/merge_stmt_1531_PhiAck/$exit
      -- CP-element group 408: 	 branch_block_stmt_783/merge_stmt_1531_PhiAck/$entry
      -- CP-element group 408: 	 branch_block_stmt_783/ifx_xend167_whilex_xend_PhiReq/$exit
      -- CP-element group 408: 	 branch_block_stmt_783/ifx_xend167_whilex_xend_PhiReq/$entry
      -- CP-element group 408: 	 branch_block_stmt_783/ifx_xend167_whilex_xend
      -- CP-element group 408: 	 branch_block_stmt_783/assign_stmt_1536/WPIPE_Block0_complete_1533_Sample/req
      -- CP-element group 408: 	 branch_block_stmt_783/assign_stmt_1536/WPIPE_Block0_complete_1533_Sample/$entry
      -- 
    if_choice_transition_3611_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 408_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1527_branch_ack_1, ack => zeropad3D_A_CP_1983_elements(408)); -- 
    req_3627_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3627_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(408), ack => WPIPE_Block0_complete_1533_inst_req_0); -- 
    -- CP-element group 409:  merge  transition  place  input  bypass 
    -- CP-element group 409: predecessors 
    -- CP-element group 409: 	1 
    -- CP-element group 409: successors 
    -- CP-element group 409:  members (5) 
      -- CP-element group 409: 	 branch_block_stmt_783/if_stmt_1527_else_link/else_choice_transition
      -- CP-element group 409: 	 branch_block_stmt_783/if_stmt_1527_else_link/$exit
      -- CP-element group 409: 	 branch_block_stmt_783/if_stmt_1527__exit__
      -- CP-element group 409: 	 branch_block_stmt_783/merge_stmt_1531__entry__
      -- CP-element group 409: 	 branch_block_stmt_783/merge_stmt_1531_dead_link/$entry
      -- 
    else_choice_transition_3615_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 409_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1527_branch_ack_0, ack => zeropad3D_A_CP_1983_elements(409)); -- 
    -- CP-element group 410:  transition  input  output  bypass 
    -- CP-element group 410: predecessors 
    -- CP-element group 410: 	408 
    -- CP-element group 410: successors 
    -- CP-element group 410: 	411 
    -- CP-element group 410:  members (6) 
      -- CP-element group 410: 	 branch_block_stmt_783/assign_stmt_1536/WPIPE_Block0_complete_1533_sample_completed_
      -- CP-element group 410: 	 branch_block_stmt_783/assign_stmt_1536/WPIPE_Block0_complete_1533_update_start_
      -- CP-element group 410: 	 branch_block_stmt_783/assign_stmt_1536/WPIPE_Block0_complete_1533_Update/req
      -- CP-element group 410: 	 branch_block_stmt_783/assign_stmt_1536/WPIPE_Block0_complete_1533_Update/$entry
      -- CP-element group 410: 	 branch_block_stmt_783/assign_stmt_1536/WPIPE_Block0_complete_1533_Sample/ack
      -- CP-element group 410: 	 branch_block_stmt_783/assign_stmt_1536/WPIPE_Block0_complete_1533_Sample/$exit
      -- 
    ack_3628_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 410_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_complete_1533_inst_ack_0, ack => zeropad3D_A_CP_1983_elements(410)); -- 
    req_3632_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3632_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => zeropad3D_A_CP_1983_elements(410), ack => WPIPE_Block0_complete_1533_inst_req_1); -- 
    -- CP-element group 411:  transition  place  input  bypass 
    -- CP-element group 411: predecessors 
    -- CP-element group 411: 	410 
    -- CP-element group 411: successors 
    -- CP-element group 411:  members (16) 
      -- CP-element group 411: 	 $exit
      -- CP-element group 411: 	 branch_block_stmt_783/$exit
      -- CP-element group 411: 	 branch_block_stmt_783/branch_block_stmt_783__exit__
      -- CP-element group 411: 	 branch_block_stmt_783/assign_stmt_1536__exit__
      -- CP-element group 411: 	 branch_block_stmt_783/return__
      -- CP-element group 411: 	 branch_block_stmt_783/merge_stmt_1538__exit__
      -- CP-element group 411: 	 branch_block_stmt_783/merge_stmt_1538_PhiReqMerge
      -- CP-element group 411: 	 branch_block_stmt_783/assign_stmt_1536/$exit
      -- CP-element group 411: 	 branch_block_stmt_783/assign_stmt_1536/WPIPE_Block0_complete_1533_update_completed_
      -- CP-element group 411: 	 branch_block_stmt_783/merge_stmt_1538_PhiAck/dummy
      -- CP-element group 411: 	 branch_block_stmt_783/merge_stmt_1538_PhiAck/$exit
      -- CP-element group 411: 	 branch_block_stmt_783/merge_stmt_1538_PhiAck/$entry
      -- CP-element group 411: 	 branch_block_stmt_783/return___PhiReq/$exit
      -- CP-element group 411: 	 branch_block_stmt_783/return___PhiReq/$entry
      -- CP-element group 411: 	 branch_block_stmt_783/assign_stmt_1536/WPIPE_Block0_complete_1533_Update/ack
      -- CP-element group 411: 	 branch_block_stmt_783/assign_stmt_1536/WPIPE_Block0_complete_1533_Update/$exit
      -- 
    ack_3633_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 411_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_complete_1533_inst_ack_1, ack => zeropad3D_A_CP_1983_elements(411)); -- 
    zeropad3D_A_do_while_stmt_903_terminator_3598: loop_terminator -- 
      generic map (name => " zeropad3D_A_do_while_stmt_903_terminator_3598", max_iterations_in_flight =>15) 
      port map(loop_body_exit => zeropad3D_A_CP_1983_elements(39),loop_continue => zeropad3D_A_CP_1983_elements(406),loop_terminate => zeropad3D_A_CP_1983_elements(405),loop_back => zeropad3D_A_CP_1983_elements(37),loop_exit => zeropad3D_A_CP_1983_elements(36),clk => clk, reset => reset); -- 
    phi_stmt_905_phi_seq_2300_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= zeropad3D_A_CP_1983_elements(52);
      zeropad3D_A_CP_1983_elements(57)<= src_sample_reqs(0);
      src_sample_acks(0)  <= zeropad3D_A_CP_1983_elements(61);
      zeropad3D_A_CP_1983_elements(58)<= src_update_reqs(0);
      src_update_acks(0)  <= zeropad3D_A_CP_1983_elements(62);
      zeropad3D_A_CP_1983_elements(53) <= phi_mux_reqs(0);
      triggers(1)  <= zeropad3D_A_CP_1983_elements(54);
      zeropad3D_A_CP_1983_elements(63)<= src_sample_reqs(1);
      src_sample_acks(1)  <= zeropad3D_A_CP_1983_elements(63);
      zeropad3D_A_CP_1983_elements(64)<= src_update_reqs(1);
      src_update_acks(1)  <= zeropad3D_A_CP_1983_elements(65);
      zeropad3D_A_CP_1983_elements(55) <= phi_mux_reqs(1);
      phi_stmt_905_phi_seq_2300 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_905_phi_seq_2300") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => zeropad3D_A_CP_1983_elements(44), 
          phi_sample_ack => zeropad3D_A_CP_1983_elements(50), 
          phi_update_req => zeropad3D_A_CP_1983_elements(46), 
          phi_update_ack => zeropad3D_A_CP_1983_elements(51), 
          phi_mux_ack => zeropad3D_A_CP_1983_elements(56), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_910_phi_seq_2344_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= zeropad3D_A_CP_1983_elements(73);
      zeropad3D_A_CP_1983_elements(78)<= src_sample_reqs(0);
      src_sample_acks(0)  <= zeropad3D_A_CP_1983_elements(82);
      zeropad3D_A_CP_1983_elements(79)<= src_update_reqs(0);
      src_update_acks(0)  <= zeropad3D_A_CP_1983_elements(83);
      zeropad3D_A_CP_1983_elements(74) <= phi_mux_reqs(0);
      triggers(1)  <= zeropad3D_A_CP_1983_elements(75);
      zeropad3D_A_CP_1983_elements(84)<= src_sample_reqs(1);
      src_sample_acks(1)  <= zeropad3D_A_CP_1983_elements(84);
      zeropad3D_A_CP_1983_elements(85)<= src_update_reqs(1);
      src_update_acks(1)  <= zeropad3D_A_CP_1983_elements(86);
      zeropad3D_A_CP_1983_elements(76) <= phi_mux_reqs(1);
      phi_stmt_910_phi_seq_2344 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_910_phi_seq_2344") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => zeropad3D_A_CP_1983_elements(69), 
          phi_sample_ack => zeropad3D_A_CP_1983_elements(70), 
          phi_update_req => zeropad3D_A_CP_1983_elements(71), 
          phi_update_ack => zeropad3D_A_CP_1983_elements(72), 
          phi_mux_ack => zeropad3D_A_CP_1983_elements(77), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_915_phi_seq_2388_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= zeropad3D_A_CP_1983_elements(94);
      zeropad3D_A_CP_1983_elements(99)<= src_sample_reqs(0);
      src_sample_acks(0)  <= zeropad3D_A_CP_1983_elements(103);
      zeropad3D_A_CP_1983_elements(100)<= src_update_reqs(0);
      src_update_acks(0)  <= zeropad3D_A_CP_1983_elements(104);
      zeropad3D_A_CP_1983_elements(95) <= phi_mux_reqs(0);
      triggers(1)  <= zeropad3D_A_CP_1983_elements(96);
      zeropad3D_A_CP_1983_elements(105)<= src_sample_reqs(1);
      src_sample_acks(1)  <= zeropad3D_A_CP_1983_elements(105);
      zeropad3D_A_CP_1983_elements(106)<= src_update_reqs(1);
      src_update_acks(1)  <= zeropad3D_A_CP_1983_elements(107);
      zeropad3D_A_CP_1983_elements(97) <= phi_mux_reqs(1);
      phi_stmt_915_phi_seq_2388 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_915_phi_seq_2388") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => zeropad3D_A_CP_1983_elements(90), 
          phi_sample_ack => zeropad3D_A_CP_1983_elements(91), 
          phi_update_req => zeropad3D_A_CP_1983_elements(92), 
          phi_update_ack => zeropad3D_A_CP_1983_elements(93), 
          phi_mux_ack => zeropad3D_A_CP_1983_elements(98), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_2252_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= zeropad3D_A_CP_1983_elements(40);
        preds(1)  <= zeropad3D_A_CP_1983_elements(41);
        entry_tmerge_2252 : transition_merge -- 
          generic map(name => " entry_tmerge_2252")
          port map (preds => preds, symbol_out => zeropad3D_A_CP_1983_elements(42));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i32_i32_1392_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1439_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1485_wire : std_logic_vector(31 downto 0);
    signal MUX_1089_wire : std_logic_vector(15 downto 0);
    signal MUX_1090_wire : std_logic_vector(15 downto 0);
    signal MUX_1117_wire : std_logic_vector(15 downto 0);
    signal MUX_1118_wire : std_logic_vector(15 downto 0);
    signal MUX_1145_wire : std_logic_vector(15 downto 0);
    signal MUX_1146_wire : std_logic_vector(15 downto 0);
    signal MUX_1167_wire : std_logic_vector(15 downto 0);
    signal MUX_1168_wire : std_logic_vector(15 downto 0);
    signal NOT_u1_u1_1050_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1292_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1362_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1066_wire : std_logic_vector(0 downto 0);
    signal R_idxprom159_1454_resized : std_logic_vector(13 downto 0);
    signal R_idxprom159_1454_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom165_1500_resized : std_logic_vector(13 downto 0);
    signal R_idxprom165_1500_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_1407_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_1407_scaled : std_logic_vector(13 downto 0);
    signal add109_1224 : std_logic_vector(15 downto 0);
    signal add118_1230 : std_logic_vector(15 downto 0);
    signal add118_1290_delayed_2_0_1422 : std_logic_vector(15 downto 0);
    signal add132_879 : std_logic_vector(31 downto 0);
    signal add149_884 : std_logic_vector(31 downto 0);
    signal add61_851 : std_logic_vector(31 downto 0);
    signal add75_860 : std_logic_vector(31 downto 0);
    signal add90_1188 : std_logic_vector(15 downto 0);
    signal add96_1194 : std_logic_vector(15 downto 0);
    signal add96_1252_delayed_2_0_1375 : std_logic_vector(15 downto 0);
    signal add96_1324_delayed_2_0_1468 : std_logic_vector(15 downto 0);
    signal add_954 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1408_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1408_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1408_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1408_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1408_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1408_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1455_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1455_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1455_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1455_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1455_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1455_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1501_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1501_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1501_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1501_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1501_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1501_root_address : std_logic_vector(13 downto 0);
    signal arrayidx160_1457 : std_logic_vector(31 downto 0);
    signal arrayidx166_1352_delayed_6_0_1509 : std_logic_vector(31 downto 0);
    signal arrayidx166_1503 : std_logic_vector(31 downto 0);
    signal arrayidx_1410 : std_logic_vector(31 downto 0);
    signal call1_789 : std_logic_vector(7 downto 0);
    signal call2_792 : std_logic_vector(7 downto 0);
    signal call3_795 : std_logic_vector(7 downto 0);
    signal call4_798 : std_logic_vector(7 downto 0);
    signal call5_801 : std_logic_vector(7 downto 0);
    signal call6_804 : std_logic_vector(7 downto 0);
    signal call_786 : std_logic_vector(7 downto 0);
    signal cmp124_1244 : std_logic_vector(0 downto 0);
    signal cmp124x_xnot_1254 : std_logic_vector(0 downto 0);
    signal cmp133_1268 : std_logic_vector(0 downto 0);
    signal cmp140_1314 : std_logic_vector(0 downto 0);
    signal cmp140x_xnot_1324 : std_logic_vector(0 downto 0);
    signal cmp150_1338 : std_logic_vector(0 downto 0);
    signal cmp62_984 : std_logic_vector(0 downto 0);
    signal cmp76_1035 : std_logic_vector(0 downto 0);
    signal cmp_934 : std_logic_vector(0 downto 0);
    signal conv106_869 : std_logic_vector(15 downto 0);
    signal conv121_1235 : std_logic_vector(31 downto 0);
    signal conv137_1305 : std_logic_vector(31 downto 0);
    signal conv154_1381 : std_logic_vector(31 downto 0);
    signal conv157_1428 : std_logic_vector(31 downto 0);
    signal conv163_1474 : std_logic_vector(31 downto 0);
    signal conv27_810 : std_logic_vector(15 downto 0);
    signal conv29_814 : std_logic_vector(15 downto 0);
    signal conv33_818 : std_logic_vector(15 downto 0);
    signal conv35_822 : std_logic_vector(15 downto 0);
    signal conv44_826 : std_logic_vector(31 downto 0);
    signal conv47_924 : std_logic_vector(31 downto 0);
    signal conv56_975 : std_logic_vector(31 downto 0);
    signal conv58_836 : std_logic_vector(31 downto 0);
    signal conv60_840 : std_logic_vector(31 downto 0);
    signal conv69_1026 : std_logic_vector(31 downto 0);
    signal conv71_855 : std_logic_vector(31 downto 0);
    signal flagx_x0_1170 : std_logic_vector(15 downto 0);
    signal idxprom159_1450 : std_logic_vector(63 downto 0);
    signal idxprom165_1496 : std_logic_vector(63 downto 0);
    signal idxprom_1403 : std_logic_vector(63 downto 0);
    signal ifx_xelse155_exec_guard_1294_delayed_1_0_1431 : std_logic_vector(0 downto 0);
    signal ifx_xelse155_exec_guard_1304_delayed_1_0_1444 : std_logic_vector(0 downto 0);
    signal ifx_xelse155_exec_guard_1317_delayed_9_0_1460 : std_logic_vector(0 downto 0);
    signal ifx_xelse155_exec_guard_1328_delayed_1_0_1477 : std_logic_vector(0 downto 0);
    signal ifx_xelse155_exec_guard_1338_delayed_1_0_1490 : std_logic_vector(0 downto 0);
    signal ifx_xelse155_exec_guard_1351_delayed_15_0_1506 : std_logic_vector(0 downto 0);
    signal ifx_xelse155_exec_guard_1419 : std_logic_vector(0 downto 0);
    signal ifx_xelse_exec_guard_1004_delayed_3_0_1038 : std_logic_vector(0 downto 0);
    signal ifx_xelse_exec_guard_1009_delayed_3_0_1046 : std_logic_vector(0 downto 0);
    signal ifx_xelse_exec_guard_960 : std_logic_vector(0 downto 0);
    signal ifx_xelse_exec_guard_967_delayed_1_0_978 : std_logic_vector(0 downto 0);
    signal ifx_xelse_exec_guard_973_delayed_1_0_987 : std_logic_vector(0 downto 0);
    signal ifx_xelse_exec_guard_978_delayed_2_0_995 : std_logic_vector(0 downto 0);
    signal ifx_xelse_exec_guard_984_delayed_1_0_1007 : std_logic_vector(0 downto 0);
    signal ifx_xelse_exec_guard_992_delayed_2_0_1021 : std_logic_vector(0 downto 0);
    signal ifx_xelse_exec_guard_997_delayed_3_0_1029 : std_logic_vector(0 downto 0);
    signal ifx_xelse_ifx_xend80_taken_1052 : std_logic_vector(0 downto 0);
    signal ifx_xelse_ifx_xthen78_taken_1043 : std_logic_vector(0 downto 0);
    signal ifx_xend167_whilex_xend_taken_1524 : std_logic_vector(0 downto 0);
    signal ifx_xend80_exec_guard_1068 : std_logic_vector(0 downto 0);
    signal ifx_xend80_exec_guard_1161_delayed_1_0_1238 : std_logic_vector(0 downto 0);
    signal ifx_xend80_exec_guard_1167_delayed_1_0_1247 : std_logic_vector(0 downto 0);
    signal ifx_xend80_exec_guard_1174_delayed_1_0_1257 : std_logic_vector(0 downto 0);
    signal ifx_xend80_exec_guard_1182_delayed_1_0_1271 : std_logic_vector(0 downto 0);
    signal ifx_xend80_exec_guard_1189_delayed_1_0_1280 : std_logic_vector(0 downto 0);
    signal ifx_xend80_exec_guard_1194_delayed_1_0_1288 : std_logic_vector(0 downto 0);
    signal ifx_xend80_ifx_xthen152_taken_1246_delayed_1_0_1367 : std_logic_vector(0 downto 0);
    signal ifx_xend80_ifx_xthen152_taken_1294 : std_logic_vector(0 downto 0);
    signal ifx_xend80_lorx_xlhsx_xfalse135_taken_1285 : std_logic_vector(0 downto 0);
    signal ifx_xthen152_exec_guard_1256_delayed_1_0_1384 : std_logic_vector(0 downto 0);
    signal ifx_xthen152_exec_guard_1266_delayed_1_0_1397 : std_logic_vector(0 downto 0);
    signal ifx_xthen152_exec_guard_1372 : std_logic_vector(0 downto 0);
    signal ifx_xthen78_exec_guard_1055 : std_logic_vector(0 downto 0);
    signal ifx_xthen78_ifx_xend80_taken_1058 : std_logic_vector(0 downto 0);
    signal ifx_xthen_exec_guard_944 : std_logic_vector(0 downto 0);
    signal ifx_xthen_ifx_xend80_taken_1022_delayed_3_0_1061 : std_logic_vector(0 downto 0);
    signal ifx_xthen_ifx_xend80_taken_1028_delayed_3_0_1071 : std_logic_vector(0 downto 0);
    signal ifx_xthen_ifx_xend80_taken_1046_delayed_3_0_1095 : std_logic_vector(0 downto 0);
    signal ifx_xthen_ifx_xend80_taken_1062_delayed_3_0_1123 : std_logic_vector(0 downto 0);
    signal ifx_xthen_ifx_xend80_taken_1078_delayed_3_0_1151 : std_logic_vector(0 downto 0);
    signal ifx_xthen_ifx_xend80_taken_957 : std_logic_vector(0 downto 0);
    signal inc67_992 : std_logic_vector(15 downto 0);
    signal inc67x_xix_x2_1004 : std_logic_vector(15 downto 0);
    signal inc_970 : std_logic_vector(15 downto 0);
    signal inc_989_delayed_1_0_1010 : std_logic_vector(15 downto 0);
    signal ix_x1_1120 : std_logic_vector(15 downto 0);
    signal ix_x2_910 : std_logic_vector(15 downto 0);
    signal ix_x2_981_delayed_3_0_998 : std_logic_vector(15 downto 0);
    signal ix_x2_at_entry_892 : std_logic_vector(15 downto 0);
    signal jx_x0_1148 : std_logic_vector(15 downto 0);
    signal jx_x0_1204_delayed_1_0_1300 : std_logic_vector(15 downto 0);
    signal jx_x1_915 : std_logic_vector(15 downto 0);
    signal jx_x1_957_delayed_1_0_963 : std_logic_vector(15 downto 0);
    signal jx_x1_at_entry_897 : std_logic_vector(15 downto 0);
    signal jx_x2_1018 : std_logic_vector(15 downto 0);
    signal kx_x0_1092 : std_logic_vector(15 downto 0);
    signal kx_x1_905 : std_logic_vector(15 downto 0);
    signal kx_x1_944_delayed_1_0_947 : std_logic_vector(15 downto 0);
    signal kx_x1_at_entry_887 : std_logic_vector(15 downto 0);
    signal lorx_xlhsx_xfalse135_exec_guard_1207_delayed_1_0_1308 : std_logic_vector(0 downto 0);
    signal lorx_xlhsx_xfalse135_exec_guard_1213_delayed_1_0_1317 : std_logic_vector(0 downto 0);
    signal lorx_xlhsx_xfalse135_exec_guard_1220_delayed_1_0_1327 : std_logic_vector(0 downto 0);
    signal lorx_xlhsx_xfalse135_exec_guard_1228_delayed_1_0_1341 : std_logic_vector(0 downto 0);
    signal lorx_xlhsx_xfalse135_exec_guard_1235_delayed_1_0_1350 : std_logic_vector(0 downto 0);
    signal lorx_xlhsx_xfalse135_exec_guard_1240_delayed_1_0_1358 : std_logic_vector(0 downto 0);
    signal lorx_xlhsx_xfalse135_exec_guard_1297 : std_logic_vector(0 downto 0);
    signal lorx_xlhsx_xfalse135_ifx_xelse155_taken_1355 : std_logic_vector(0 downto 0);
    signal lorx_xlhsx_xfalse135_ifx_xthen152_taken_1364 : std_logic_vector(0 downto 0);
    signal mul108_1206 : std_logic_vector(15 downto 0);
    signal mul117_1218 : std_logic_vector(15 downto 0);
    signal mul36_865 : std_logic_vector(15 downto 0);
    signal mul89_1176 : std_logic_vector(15 downto 0);
    signal mul95_1182 : std_logic_vector(15 downto 0);
    signal mul_874 : std_logic_vector(15 downto 0);
    signal orx_xcond171_1347 : std_logic_vector(0 downto 0);
    signal orx_xcond_1277 : std_logic_vector(0 downto 0);
    signal ptr_deref_1413_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1413_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1413_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1413_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1413_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1413_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1464_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1464_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1464_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1464_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1464_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1512_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1512_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1512_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1512_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1512_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1512_word_offset_0 : std_logic_vector(13 downto 0);
    signal shl_846 : std_logic_vector(31 downto 0);
    signal shr158_1441 : std_logic_vector(31 downto 0);
    signal shr164_1487 : std_logic_vector(31 downto 0);
    signal shr_1394 : std_logic_vector(31 downto 0);
    signal sub107_1200 : std_logic_vector(15 downto 0);
    signal sub116_1212 : std_logic_vector(15 downto 0);
    signal sub_832 : std_logic_vector(31 downto 0);
    signal tmp161_1465 : std_logic_vector(63 downto 0);
    signal tobool_1520 : std_logic_vector(0 downto 0);
    signal type_cast_1015_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1030_1030_delayed_3_0_1075 : std_logic_vector(15 downto 0);
    signal type_cast_1048_1048_delayed_4_0_1099 : std_logic_vector(15 downto 0);
    signal type_cast_1051_1051_delayed_1_0_1103 : std_logic_vector(15 downto 0);
    signal type_cast_1054_1054_delayed_1_0_1107 : std_logic_vector(15 downto 0);
    signal type_cast_1064_1064_delayed_4_0_1127 : std_logic_vector(15 downto 0);
    signal type_cast_1067_1067_delayed_2_0_1131 : std_logic_vector(15 downto 0);
    signal type_cast_1070_1070_delayed_2_0_1135 : std_logic_vector(15 downto 0);
    signal type_cast_1082_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1086_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1088_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1116_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1144_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1156_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1160_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1164_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1166_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1179_1179_delayed_1_0_1261 : std_logic_vector(31 downto 0);
    signal type_cast_1225_1225_delayed_1_0_1331 : std_logic_vector(31 downto 0);
    signal type_cast_1252_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1265_wire : std_logic_vector(31 downto 0);
    signal type_cast_1322_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1335_wire : std_logic_vector(31 downto 0);
    signal type_cast_1379_wire : std_logic_vector(31 downto 0);
    signal type_cast_1388_wire : std_logic_vector(31 downto 0);
    signal type_cast_1391_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1401_wire : std_logic_vector(63 downto 0);
    signal type_cast_1415_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1426_wire : std_logic_vector(31 downto 0);
    signal type_cast_1435_wire : std_logic_vector(31 downto 0);
    signal type_cast_1438_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1448_wire : std_logic_vector(63 downto 0);
    signal type_cast_1472_wire : std_logic_vector(31 downto 0);
    signal type_cast_1481_wire : std_logic_vector(31 downto 0);
    signal type_cast_1484_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1494_wire : std_logic_vector(63 downto 0);
    signal type_cast_1518_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1535_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_830_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_844_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_908_wire : std_logic_vector(15 downto 0);
    signal type_cast_913_wire : std_logic_vector(15 downto 0);
    signal type_cast_918_wire : std_logic_vector(15 downto 0);
    signal type_cast_929_929_delayed_2_0_928 : std_logic_vector(31 downto 0);
    signal type_cast_931_wire : std_logic_vector(31 downto 0);
    signal type_cast_952_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_968_wire_constant : std_logic_vector(15 downto 0);
    signal whilex_xbody_ifx_xelse_taken_937 : std_logic_vector(0 downto 0);
    signal whilex_xbody_ifx_xthen_taken_941 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    array_obj_ref_1408_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1408_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1408_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1408_resized_base_address <= "00000000000000";
    array_obj_ref_1455_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1455_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1455_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1455_resized_base_address <= "00000000000000";
    array_obj_ref_1501_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1501_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1501_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1501_resized_base_address <= "00000000000000";
    ix_x2_at_entry_892 <= "0000000000000000";
    jx_x1_at_entry_897 <= "0000000000000000";
    kx_x1_at_entry_887 <= "0000000000000000";
    ptr_deref_1413_word_offset_0 <= "00000000000000";
    ptr_deref_1464_word_offset_0 <= "00000000000000";
    ptr_deref_1512_word_offset_0 <= "00000000000000";
    type_cast_1015_wire_constant <= "0000000000000000";
    type_cast_1082_wire_constant <= "0000000000000000";
    type_cast_1086_wire_constant <= "0000000000000000";
    type_cast_1088_wire_constant <= "0000000000000000";
    type_cast_1116_wire_constant <= "0000000000000000";
    type_cast_1144_wire_constant <= "0000000000000000";
    type_cast_1156_wire_constant <= "0000000000000000";
    type_cast_1160_wire_constant <= "0000000000000001";
    type_cast_1164_wire_constant <= "0000000000000000";
    type_cast_1166_wire_constant <= "0000000000000000";
    type_cast_1252_wire_constant <= "1";
    type_cast_1322_wire_constant <= "1";
    type_cast_1391_wire_constant <= "00000000000000000000000000000011";
    type_cast_1415_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1438_wire_constant <= "00000000000000000000000000000011";
    type_cast_1484_wire_constant <= "00000000000000000000000000000011";
    type_cast_1518_wire_constant <= "0000000000000000";
    type_cast_1535_wire_constant <= "00000001";
    type_cast_830_wire_constant <= "11111111111111111111111111111000";
    type_cast_844_wire_constant <= "00000000000000000000000000000001";
    type_cast_952_wire_constant <= "0000000000001000";
    type_cast_968_wire_constant <= "0000000000000001";
    phi_stmt_905: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_908_wire & kx_x1_at_entry_887;
      req <= phi_stmt_905_req_0 & phi_stmt_905_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_905",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_905_ack_0,
          idata => idata,
          odata => kx_x1_905,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_905
    phi_stmt_910: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_913_wire & ix_x2_at_entry_892;
      req <= phi_stmt_910_req_0 & phi_stmt_910_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_910",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_910_ack_0,
          idata => idata,
          odata => ix_x2_910,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_910
    phi_stmt_915: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_918_wire & jx_x1_at_entry_897;
      req <= phi_stmt_915_req_0 & phi_stmt_915_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_915",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_915_ack_0,
          idata => idata,
          odata => jx_x1_915,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_915
    -- flow-through select operator MUX_1017_inst
    jx_x2_1018 <= type_cast_1015_wire_constant when (cmp62_984(0) /=  '0') else inc_989_delayed_1_0_1010;
    -- flow-through select operator MUX_1089_inst
    MUX_1089_wire <= type_cast_1086_wire_constant when (ifx_xelse_ifx_xend80_taken_1052(0) /=  '0') else type_cast_1088_wire_constant;
    -- flow-through select operator MUX_1090_inst
    MUX_1090_wire <= type_cast_1082_wire_constant when (ifx_xthen78_ifx_xend80_taken_1058(0) /=  '0') else MUX_1089_wire;
    -- flow-through select operator MUX_1091_inst
    kx_x0_1092 <= type_cast_1030_1030_delayed_3_0_1075 when (ifx_xthen_ifx_xend80_taken_1028_delayed_3_0_1071(0) /=  '0') else MUX_1090_wire;
    -- flow-through select operator MUX_1117_inst
    MUX_1117_wire <= type_cast_1054_1054_delayed_1_0_1107 when (ifx_xelse_ifx_xend80_taken_1052(0) /=  '0') else type_cast_1116_wire_constant;
    -- flow-through select operator MUX_1118_inst
    MUX_1118_wire <= type_cast_1051_1051_delayed_1_0_1103 when (ifx_xthen78_ifx_xend80_taken_1058(0) /=  '0') else MUX_1117_wire;
    -- flow-through select operator MUX_1119_inst
    ix_x1_1120 <= type_cast_1048_1048_delayed_4_0_1099 when (ifx_xthen_ifx_xend80_taken_1046_delayed_3_0_1095(0) /=  '0') else MUX_1118_wire;
    -- flow-through select operator MUX_1145_inst
    MUX_1145_wire <= type_cast_1070_1070_delayed_2_0_1135 when (ifx_xelse_ifx_xend80_taken_1052(0) /=  '0') else type_cast_1144_wire_constant;
    -- flow-through select operator MUX_1146_inst
    MUX_1146_wire <= type_cast_1067_1067_delayed_2_0_1131 when (ifx_xthen78_ifx_xend80_taken_1058(0) /=  '0') else MUX_1145_wire;
    -- flow-through select operator MUX_1147_inst
    jx_x0_1148 <= type_cast_1064_1064_delayed_4_0_1127 when (ifx_xthen_ifx_xend80_taken_1062_delayed_3_0_1123(0) /=  '0') else MUX_1146_wire;
    -- flow-through select operator MUX_1167_inst
    MUX_1167_wire <= type_cast_1164_wire_constant when (ifx_xelse_ifx_xend80_taken_1052(0) /=  '0') else type_cast_1166_wire_constant;
    -- flow-through select operator MUX_1168_inst
    MUX_1168_wire <= type_cast_1160_wire_constant when (ifx_xthen78_ifx_xend80_taken_1058(0) /=  '0') else MUX_1167_wire;
    -- flow-through select operator MUX_1169_inst
    flagx_x0_1170 <= type_cast_1156_wire_constant when (ifx_xthen_ifx_xend80_taken_1078_delayed_3_0_1151(0) /=  '0') else MUX_1168_wire;
    W_add118_1290_delayed_2_0_1420_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_add118_1290_delayed_2_0_1420_inst_req_0;
      W_add118_1290_delayed_2_0_1420_inst_ack_0<= wack(0);
      rreq(0) <= W_add118_1290_delayed_2_0_1420_inst_req_1;
      W_add118_1290_delayed_2_0_1420_inst_ack_1<= rack(0);
      W_add118_1290_delayed_2_0_1420_inst : InterlockBuffer generic map ( -- 
        name => "W_add118_1290_delayed_2_0_1420_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add118_1230,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => add118_1290_delayed_2_0_1422,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_add96_1252_delayed_2_0_1373_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_add96_1252_delayed_2_0_1373_inst_req_0;
      W_add96_1252_delayed_2_0_1373_inst_ack_0<= wack(0);
      rreq(0) <= W_add96_1252_delayed_2_0_1373_inst_req_1;
      W_add96_1252_delayed_2_0_1373_inst_ack_1<= rack(0);
      W_add96_1252_delayed_2_0_1373_inst : InterlockBuffer generic map ( -- 
        name => "W_add96_1252_delayed_2_0_1373_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add96_1194,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => add96_1252_delayed_2_0_1375,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_add96_1324_delayed_2_0_1466_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_add96_1324_delayed_2_0_1466_inst_req_0;
      W_add96_1324_delayed_2_0_1466_inst_ack_0<= wack(0);
      rreq(0) <= W_add96_1324_delayed_2_0_1466_inst_req_1;
      W_add96_1324_delayed_2_0_1466_inst_ack_1<= rack(0);
      W_add96_1324_delayed_2_0_1466_inst : InterlockBuffer generic map ( -- 
        name => "W_add96_1324_delayed_2_0_1466_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add96_1194,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => add96_1324_delayed_2_0_1468,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_arrayidx166_1352_delayed_6_0_1507_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_arrayidx166_1352_delayed_6_0_1507_inst_req_0;
      W_arrayidx166_1352_delayed_6_0_1507_inst_ack_0<= wack(0);
      rreq(0) <= W_arrayidx166_1352_delayed_6_0_1507_inst_req_1;
      W_arrayidx166_1352_delayed_6_0_1507_inst_ack_1<= rack(0);
      W_arrayidx166_1352_delayed_6_0_1507_inst : InterlockBuffer generic map ( -- 
        name => "W_arrayidx166_1352_delayed_6_0_1507_inst",
        buffer_size => 6,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => arrayidx166_1503,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx166_1352_delayed_6_0_1509,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xelse155_exec_guard_1294_delayed_1_0_1429_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xelse155_exec_guard_1294_delayed_1_0_1429_inst_req_0;
      W_ifx_xelse155_exec_guard_1294_delayed_1_0_1429_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xelse155_exec_guard_1294_delayed_1_0_1429_inst_req_1;
      W_ifx_xelse155_exec_guard_1294_delayed_1_0_1429_inst_ack_1<= rack(0);
      W_ifx_xelse155_exec_guard_1294_delayed_1_0_1429_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xelse155_exec_guard_1294_delayed_1_0_1429_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xelse155_exec_guard_1419,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xelse155_exec_guard_1294_delayed_1_0_1431,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xelse155_exec_guard_1304_delayed_1_0_1442_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xelse155_exec_guard_1304_delayed_1_0_1442_inst_req_0;
      W_ifx_xelse155_exec_guard_1304_delayed_1_0_1442_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xelse155_exec_guard_1304_delayed_1_0_1442_inst_req_1;
      W_ifx_xelse155_exec_guard_1304_delayed_1_0_1442_inst_ack_1<= rack(0);
      W_ifx_xelse155_exec_guard_1304_delayed_1_0_1442_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xelse155_exec_guard_1304_delayed_1_0_1442_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xelse155_exec_guard_1419,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xelse155_exec_guard_1304_delayed_1_0_1444,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xelse155_exec_guard_1317_delayed_9_0_1458_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xelse155_exec_guard_1317_delayed_9_0_1458_inst_req_0;
      W_ifx_xelse155_exec_guard_1317_delayed_9_0_1458_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xelse155_exec_guard_1317_delayed_9_0_1458_inst_req_1;
      W_ifx_xelse155_exec_guard_1317_delayed_9_0_1458_inst_ack_1<= rack(0);
      W_ifx_xelse155_exec_guard_1317_delayed_9_0_1458_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xelse155_exec_guard_1317_delayed_9_0_1458_inst",
        buffer_size => 9,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xelse155_exec_guard_1419,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xelse155_exec_guard_1317_delayed_9_0_1460,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xelse155_exec_guard_1328_delayed_1_0_1475_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xelse155_exec_guard_1328_delayed_1_0_1475_inst_req_0;
      W_ifx_xelse155_exec_guard_1328_delayed_1_0_1475_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xelse155_exec_guard_1328_delayed_1_0_1475_inst_req_1;
      W_ifx_xelse155_exec_guard_1328_delayed_1_0_1475_inst_ack_1<= rack(0);
      W_ifx_xelse155_exec_guard_1328_delayed_1_0_1475_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xelse155_exec_guard_1328_delayed_1_0_1475_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xelse155_exec_guard_1419,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xelse155_exec_guard_1328_delayed_1_0_1477,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xelse155_exec_guard_1338_delayed_1_0_1488_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xelse155_exec_guard_1338_delayed_1_0_1488_inst_req_0;
      W_ifx_xelse155_exec_guard_1338_delayed_1_0_1488_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xelse155_exec_guard_1338_delayed_1_0_1488_inst_req_1;
      W_ifx_xelse155_exec_guard_1338_delayed_1_0_1488_inst_ack_1<= rack(0);
      W_ifx_xelse155_exec_guard_1338_delayed_1_0_1488_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xelse155_exec_guard_1338_delayed_1_0_1488_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xelse155_exec_guard_1419,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xelse155_exec_guard_1338_delayed_1_0_1490,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xelse155_exec_guard_1351_delayed_15_0_1504_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xelse155_exec_guard_1351_delayed_15_0_1504_inst_req_0;
      W_ifx_xelse155_exec_guard_1351_delayed_15_0_1504_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xelse155_exec_guard_1351_delayed_15_0_1504_inst_req_1;
      W_ifx_xelse155_exec_guard_1351_delayed_15_0_1504_inst_ack_1<= rack(0);
      W_ifx_xelse155_exec_guard_1351_delayed_15_0_1504_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xelse155_exec_guard_1351_delayed_15_0_1504_inst",
        buffer_size => 15,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xelse155_exec_guard_1419,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xelse155_exec_guard_1351_delayed_15_0_1506,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock W_ifx_xelse155_exec_guard_1417_inst
    process(lorx_xlhsx_xfalse135_ifx_xelse155_taken_1355) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := lorx_xlhsx_xfalse135_ifx_xelse155_taken_1355(0 downto 0);
      ifx_xelse155_exec_guard_1419 <= tmp_var; -- 
    end process;
    W_ifx_xelse_exec_guard_1004_delayed_3_0_1036_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xelse_exec_guard_1004_delayed_3_0_1036_inst_req_0;
      W_ifx_xelse_exec_guard_1004_delayed_3_0_1036_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xelse_exec_guard_1004_delayed_3_0_1036_inst_req_1;
      W_ifx_xelse_exec_guard_1004_delayed_3_0_1036_inst_ack_1<= rack(0);
      W_ifx_xelse_exec_guard_1004_delayed_3_0_1036_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xelse_exec_guard_1004_delayed_3_0_1036_inst",
        buffer_size => 3,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xelse_exec_guard_960,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xelse_exec_guard_1004_delayed_3_0_1038,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xelse_exec_guard_1009_delayed_3_0_1044_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xelse_exec_guard_1009_delayed_3_0_1044_inst_req_0;
      W_ifx_xelse_exec_guard_1009_delayed_3_0_1044_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xelse_exec_guard_1009_delayed_3_0_1044_inst_req_1;
      W_ifx_xelse_exec_guard_1009_delayed_3_0_1044_inst_ack_1<= rack(0);
      W_ifx_xelse_exec_guard_1009_delayed_3_0_1044_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xelse_exec_guard_1009_delayed_3_0_1044_inst",
        buffer_size => 3,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xelse_exec_guard_960,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xelse_exec_guard_1009_delayed_3_0_1046,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock W_ifx_xelse_exec_guard_958_inst
    process(whilex_xbody_ifx_xelse_taken_937) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := whilex_xbody_ifx_xelse_taken_937(0 downto 0);
      ifx_xelse_exec_guard_960 <= tmp_var; -- 
    end process;
    W_ifx_xelse_exec_guard_967_delayed_1_0_976_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xelse_exec_guard_967_delayed_1_0_976_inst_req_0;
      W_ifx_xelse_exec_guard_967_delayed_1_0_976_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xelse_exec_guard_967_delayed_1_0_976_inst_req_1;
      W_ifx_xelse_exec_guard_967_delayed_1_0_976_inst_ack_1<= rack(0);
      W_ifx_xelse_exec_guard_967_delayed_1_0_976_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xelse_exec_guard_967_delayed_1_0_976_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xelse_exec_guard_960,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xelse_exec_guard_967_delayed_1_0_978,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xelse_exec_guard_973_delayed_1_0_985_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xelse_exec_guard_973_delayed_1_0_985_inst_req_0;
      W_ifx_xelse_exec_guard_973_delayed_1_0_985_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xelse_exec_guard_973_delayed_1_0_985_inst_req_1;
      W_ifx_xelse_exec_guard_973_delayed_1_0_985_inst_ack_1<= rack(0);
      W_ifx_xelse_exec_guard_973_delayed_1_0_985_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xelse_exec_guard_973_delayed_1_0_985_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xelse_exec_guard_960,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xelse_exec_guard_973_delayed_1_0_987,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xelse_exec_guard_978_delayed_2_0_993_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xelse_exec_guard_978_delayed_2_0_993_inst_req_0;
      W_ifx_xelse_exec_guard_978_delayed_2_0_993_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xelse_exec_guard_978_delayed_2_0_993_inst_req_1;
      W_ifx_xelse_exec_guard_978_delayed_2_0_993_inst_ack_1<= rack(0);
      W_ifx_xelse_exec_guard_978_delayed_2_0_993_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xelse_exec_guard_978_delayed_2_0_993_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xelse_exec_guard_960,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xelse_exec_guard_978_delayed_2_0_995,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xelse_exec_guard_984_delayed_1_0_1005_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xelse_exec_guard_984_delayed_1_0_1005_inst_req_0;
      W_ifx_xelse_exec_guard_984_delayed_1_0_1005_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xelse_exec_guard_984_delayed_1_0_1005_inst_req_1;
      W_ifx_xelse_exec_guard_984_delayed_1_0_1005_inst_ack_1<= rack(0);
      W_ifx_xelse_exec_guard_984_delayed_1_0_1005_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xelse_exec_guard_984_delayed_1_0_1005_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xelse_exec_guard_960,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xelse_exec_guard_984_delayed_1_0_1007,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xelse_exec_guard_992_delayed_2_0_1019_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xelse_exec_guard_992_delayed_2_0_1019_inst_req_0;
      W_ifx_xelse_exec_guard_992_delayed_2_0_1019_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xelse_exec_guard_992_delayed_2_0_1019_inst_req_1;
      W_ifx_xelse_exec_guard_992_delayed_2_0_1019_inst_ack_1<= rack(0);
      W_ifx_xelse_exec_guard_992_delayed_2_0_1019_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xelse_exec_guard_992_delayed_2_0_1019_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xelse_exec_guard_960,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xelse_exec_guard_992_delayed_2_0_1021,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xelse_exec_guard_997_delayed_3_0_1027_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xelse_exec_guard_997_delayed_3_0_1027_inst_req_0;
      W_ifx_xelse_exec_guard_997_delayed_3_0_1027_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xelse_exec_guard_997_delayed_3_0_1027_inst_req_1;
      W_ifx_xelse_exec_guard_997_delayed_3_0_1027_inst_ack_1<= rack(0);
      W_ifx_xelse_exec_guard_997_delayed_3_0_1027_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xelse_exec_guard_997_delayed_3_0_1027_inst",
        buffer_size => 3,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xelse_exec_guard_960,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xelse_exec_guard_997_delayed_3_0_1029,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xend80_exec_guard_1161_delayed_1_0_1236_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xend80_exec_guard_1161_delayed_1_0_1236_inst_req_0;
      W_ifx_xend80_exec_guard_1161_delayed_1_0_1236_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xend80_exec_guard_1161_delayed_1_0_1236_inst_req_1;
      W_ifx_xend80_exec_guard_1161_delayed_1_0_1236_inst_ack_1<= rack(0);
      W_ifx_xend80_exec_guard_1161_delayed_1_0_1236_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xend80_exec_guard_1161_delayed_1_0_1236_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xend80_exec_guard_1068,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xend80_exec_guard_1161_delayed_1_0_1238,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xend80_exec_guard_1167_delayed_1_0_1245_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xend80_exec_guard_1167_delayed_1_0_1245_inst_req_0;
      W_ifx_xend80_exec_guard_1167_delayed_1_0_1245_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xend80_exec_guard_1167_delayed_1_0_1245_inst_req_1;
      W_ifx_xend80_exec_guard_1167_delayed_1_0_1245_inst_ack_1<= rack(0);
      W_ifx_xend80_exec_guard_1167_delayed_1_0_1245_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xend80_exec_guard_1167_delayed_1_0_1245_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xend80_exec_guard_1068,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xend80_exec_guard_1167_delayed_1_0_1247,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xend80_exec_guard_1174_delayed_1_0_1255_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xend80_exec_guard_1174_delayed_1_0_1255_inst_req_0;
      W_ifx_xend80_exec_guard_1174_delayed_1_0_1255_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xend80_exec_guard_1174_delayed_1_0_1255_inst_req_1;
      W_ifx_xend80_exec_guard_1174_delayed_1_0_1255_inst_ack_1<= rack(0);
      W_ifx_xend80_exec_guard_1174_delayed_1_0_1255_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xend80_exec_guard_1174_delayed_1_0_1255_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xend80_exec_guard_1068,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xend80_exec_guard_1174_delayed_1_0_1257,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xend80_exec_guard_1182_delayed_1_0_1269_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xend80_exec_guard_1182_delayed_1_0_1269_inst_req_0;
      W_ifx_xend80_exec_guard_1182_delayed_1_0_1269_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xend80_exec_guard_1182_delayed_1_0_1269_inst_req_1;
      W_ifx_xend80_exec_guard_1182_delayed_1_0_1269_inst_ack_1<= rack(0);
      W_ifx_xend80_exec_guard_1182_delayed_1_0_1269_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xend80_exec_guard_1182_delayed_1_0_1269_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xend80_exec_guard_1068,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xend80_exec_guard_1182_delayed_1_0_1271,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xend80_exec_guard_1189_delayed_1_0_1278_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xend80_exec_guard_1189_delayed_1_0_1278_inst_req_0;
      W_ifx_xend80_exec_guard_1189_delayed_1_0_1278_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xend80_exec_guard_1189_delayed_1_0_1278_inst_req_1;
      W_ifx_xend80_exec_guard_1189_delayed_1_0_1278_inst_ack_1<= rack(0);
      W_ifx_xend80_exec_guard_1189_delayed_1_0_1278_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xend80_exec_guard_1189_delayed_1_0_1278_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xend80_exec_guard_1068,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xend80_exec_guard_1189_delayed_1_0_1280,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xend80_exec_guard_1194_delayed_1_0_1286_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xend80_exec_guard_1194_delayed_1_0_1286_inst_req_0;
      W_ifx_xend80_exec_guard_1194_delayed_1_0_1286_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xend80_exec_guard_1194_delayed_1_0_1286_inst_req_1;
      W_ifx_xend80_exec_guard_1194_delayed_1_0_1286_inst_ack_1<= rack(0);
      W_ifx_xend80_exec_guard_1194_delayed_1_0_1286_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xend80_exec_guard_1194_delayed_1_0_1286_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xend80_exec_guard_1068,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xend80_exec_guard_1194_delayed_1_0_1288,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xend80_ifx_xthen152_taken_1246_delayed_1_0_1365_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xend80_ifx_xthen152_taken_1246_delayed_1_0_1365_inst_req_0;
      W_ifx_xend80_ifx_xthen152_taken_1246_delayed_1_0_1365_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xend80_ifx_xthen152_taken_1246_delayed_1_0_1365_inst_req_1;
      W_ifx_xend80_ifx_xthen152_taken_1246_delayed_1_0_1365_inst_ack_1<= rack(0);
      W_ifx_xend80_ifx_xthen152_taken_1246_delayed_1_0_1365_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xend80_ifx_xthen152_taken_1246_delayed_1_0_1365_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xend80_ifx_xthen152_taken_1294,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xend80_ifx_xthen152_taken_1246_delayed_1_0_1367,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xthen152_exec_guard_1256_delayed_1_0_1382_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xthen152_exec_guard_1256_delayed_1_0_1382_inst_req_0;
      W_ifx_xthen152_exec_guard_1256_delayed_1_0_1382_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xthen152_exec_guard_1256_delayed_1_0_1382_inst_req_1;
      W_ifx_xthen152_exec_guard_1256_delayed_1_0_1382_inst_ack_1<= rack(0);
      W_ifx_xthen152_exec_guard_1256_delayed_1_0_1382_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xthen152_exec_guard_1256_delayed_1_0_1382_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xthen152_exec_guard_1372,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xthen152_exec_guard_1256_delayed_1_0_1384,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xthen152_exec_guard_1266_delayed_1_0_1395_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xthen152_exec_guard_1266_delayed_1_0_1395_inst_req_0;
      W_ifx_xthen152_exec_guard_1266_delayed_1_0_1395_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xthen152_exec_guard_1266_delayed_1_0_1395_inst_req_1;
      W_ifx_xthen152_exec_guard_1266_delayed_1_0_1395_inst_ack_1<= rack(0);
      W_ifx_xthen152_exec_guard_1266_delayed_1_0_1395_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xthen152_exec_guard_1266_delayed_1_0_1395_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xthen152_exec_guard_1372,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xthen152_exec_guard_1266_delayed_1_0_1397,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock W_ifx_xthen78_exec_guard_1053_inst
    process(ifx_xelse_ifx_xthen78_taken_1043) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := ifx_xelse_ifx_xthen78_taken_1043(0 downto 0);
      ifx_xthen78_exec_guard_1055 <= tmp_var; -- 
    end process;
    -- interlock W_ifx_xthen78_ifx_xend80_taken_1056_inst
    process(ifx_xthen78_exec_guard_1055) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := ifx_xthen78_exec_guard_1055(0 downto 0);
      ifx_xthen78_ifx_xend80_taken_1058 <= tmp_var; -- 
    end process;
    -- interlock W_ifx_xthen_exec_guard_942_inst
    process(whilex_xbody_ifx_xthen_taken_941) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := whilex_xbody_ifx_xthen_taken_941(0 downto 0);
      ifx_xthen_exec_guard_944 <= tmp_var; -- 
    end process;
    W_ifx_xthen_ifx_xend80_taken_1022_delayed_3_0_1059_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xthen_ifx_xend80_taken_1022_delayed_3_0_1059_inst_req_0;
      W_ifx_xthen_ifx_xend80_taken_1022_delayed_3_0_1059_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xthen_ifx_xend80_taken_1022_delayed_3_0_1059_inst_req_1;
      W_ifx_xthen_ifx_xend80_taken_1022_delayed_3_0_1059_inst_ack_1<= rack(0);
      W_ifx_xthen_ifx_xend80_taken_1022_delayed_3_0_1059_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xthen_ifx_xend80_taken_1022_delayed_3_0_1059_inst",
        buffer_size => 3,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xthen_ifx_xend80_taken_957,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xthen_ifx_xend80_taken_1022_delayed_3_0_1061,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xthen_ifx_xend80_taken_1028_delayed_3_0_1069_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xthen_ifx_xend80_taken_1028_delayed_3_0_1069_inst_req_0;
      W_ifx_xthen_ifx_xend80_taken_1028_delayed_3_0_1069_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xthen_ifx_xend80_taken_1028_delayed_3_0_1069_inst_req_1;
      W_ifx_xthen_ifx_xend80_taken_1028_delayed_3_0_1069_inst_ack_1<= rack(0);
      W_ifx_xthen_ifx_xend80_taken_1028_delayed_3_0_1069_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xthen_ifx_xend80_taken_1028_delayed_3_0_1069_inst",
        buffer_size => 3,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xthen_ifx_xend80_taken_957,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xthen_ifx_xend80_taken_1028_delayed_3_0_1071,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xthen_ifx_xend80_taken_1046_delayed_3_0_1093_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xthen_ifx_xend80_taken_1046_delayed_3_0_1093_inst_req_0;
      W_ifx_xthen_ifx_xend80_taken_1046_delayed_3_0_1093_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xthen_ifx_xend80_taken_1046_delayed_3_0_1093_inst_req_1;
      W_ifx_xthen_ifx_xend80_taken_1046_delayed_3_0_1093_inst_ack_1<= rack(0);
      W_ifx_xthen_ifx_xend80_taken_1046_delayed_3_0_1093_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xthen_ifx_xend80_taken_1046_delayed_3_0_1093_inst",
        buffer_size => 3,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xthen_ifx_xend80_taken_957,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xthen_ifx_xend80_taken_1046_delayed_3_0_1095,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xthen_ifx_xend80_taken_1062_delayed_3_0_1121_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xthen_ifx_xend80_taken_1062_delayed_3_0_1121_inst_req_0;
      W_ifx_xthen_ifx_xend80_taken_1062_delayed_3_0_1121_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xthen_ifx_xend80_taken_1062_delayed_3_0_1121_inst_req_1;
      W_ifx_xthen_ifx_xend80_taken_1062_delayed_3_0_1121_inst_ack_1<= rack(0);
      W_ifx_xthen_ifx_xend80_taken_1062_delayed_3_0_1121_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xthen_ifx_xend80_taken_1062_delayed_3_0_1121_inst",
        buffer_size => 3,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xthen_ifx_xend80_taken_957,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xthen_ifx_xend80_taken_1062_delayed_3_0_1123,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ifx_xthen_ifx_xend80_taken_1078_delayed_3_0_1149_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ifx_xthen_ifx_xend80_taken_1078_delayed_3_0_1149_inst_req_0;
      W_ifx_xthen_ifx_xend80_taken_1078_delayed_3_0_1149_inst_ack_0<= wack(0);
      rreq(0) <= W_ifx_xthen_ifx_xend80_taken_1078_delayed_3_0_1149_inst_req_1;
      W_ifx_xthen_ifx_xend80_taken_1078_delayed_3_0_1149_inst_ack_1<= rack(0);
      W_ifx_xthen_ifx_xend80_taken_1078_delayed_3_0_1149_inst : InterlockBuffer generic map ( -- 
        name => "W_ifx_xthen_ifx_xend80_taken_1078_delayed_3_0_1149_inst",
        buffer_size => 3,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ifx_xthen_ifx_xend80_taken_957,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ifx_xthen_ifx_xend80_taken_1078_delayed_3_0_1151,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock W_ifx_xthen_ifx_xend80_taken_955_inst
    process(ifx_xthen_exec_guard_944) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := ifx_xthen_exec_guard_944(0 downto 0);
      ifx_xthen_ifx_xend80_taken_957 <= tmp_var; -- 
    end process;
    W_inc_989_delayed_1_0_1008_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_inc_989_delayed_1_0_1008_inst_req_0;
      W_inc_989_delayed_1_0_1008_inst_ack_0<= wack(0);
      rreq(0) <= W_inc_989_delayed_1_0_1008_inst_req_1;
      W_inc_989_delayed_1_0_1008_inst_ack_1<= rack(0);
      W_inc_989_delayed_1_0_1008_inst : InterlockBuffer generic map ( -- 
        name => "W_inc_989_delayed_1_0_1008_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc_970,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc_989_delayed_1_0_1010,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_ix_x2_981_delayed_3_0_996_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_ix_x2_981_delayed_3_0_996_inst_req_0;
      W_ix_x2_981_delayed_3_0_996_inst_ack_0<= wack(0);
      rreq(0) <= W_ix_x2_981_delayed_3_0_996_inst_req_1;
      W_ix_x2_981_delayed_3_0_996_inst_ack_1<= rack(0);
      W_ix_x2_981_delayed_3_0_996_inst : InterlockBuffer generic map ( -- 
        name => "W_ix_x2_981_delayed_3_0_996_inst",
        buffer_size => 3,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ix_x2_910,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ix_x2_981_delayed_3_0_998,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_jx_x0_1204_delayed_1_0_1298_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_jx_x0_1204_delayed_1_0_1298_inst_req_0;
      W_jx_x0_1204_delayed_1_0_1298_inst_ack_0<= wack(0);
      rreq(0) <= W_jx_x0_1204_delayed_1_0_1298_inst_req_1;
      W_jx_x0_1204_delayed_1_0_1298_inst_ack_1<= rack(0);
      W_jx_x0_1204_delayed_1_0_1298_inst : InterlockBuffer generic map ( -- 
        name => "W_jx_x0_1204_delayed_1_0_1298_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x0_1148,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => jx_x0_1204_delayed_1_0_1300,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_jx_x1_957_delayed_1_0_961_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_jx_x1_957_delayed_1_0_961_inst_req_0;
      W_jx_x1_957_delayed_1_0_961_inst_ack_0<= wack(0);
      rreq(0) <= W_jx_x1_957_delayed_1_0_961_inst_req_1;
      W_jx_x1_957_delayed_1_0_961_inst_ack_1<= rack(0);
      W_jx_x1_957_delayed_1_0_961_inst : InterlockBuffer generic map ( -- 
        name => "W_jx_x1_957_delayed_1_0_961_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x1_915,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => jx_x1_957_delayed_1_0_963,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_kx_x1_944_delayed_1_0_945_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_kx_x1_944_delayed_1_0_945_inst_req_0;
      W_kx_x1_944_delayed_1_0_945_inst_ack_0<= wack(0);
      rreq(0) <= W_kx_x1_944_delayed_1_0_945_inst_req_1;
      W_kx_x1_944_delayed_1_0_945_inst_ack_1<= rack(0);
      W_kx_x1_944_delayed_1_0_945_inst : InterlockBuffer generic map ( -- 
        name => "W_kx_x1_944_delayed_1_0_945_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => kx_x1_905,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => kx_x1_944_delayed_1_0_947,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_lorx_xlhsx_xfalse135_exec_guard_1207_delayed_1_0_1306_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_lorx_xlhsx_xfalse135_exec_guard_1207_delayed_1_0_1306_inst_req_0;
      W_lorx_xlhsx_xfalse135_exec_guard_1207_delayed_1_0_1306_inst_ack_0<= wack(0);
      rreq(0) <= W_lorx_xlhsx_xfalse135_exec_guard_1207_delayed_1_0_1306_inst_req_1;
      W_lorx_xlhsx_xfalse135_exec_guard_1207_delayed_1_0_1306_inst_ack_1<= rack(0);
      W_lorx_xlhsx_xfalse135_exec_guard_1207_delayed_1_0_1306_inst : InterlockBuffer generic map ( -- 
        name => "W_lorx_xlhsx_xfalse135_exec_guard_1207_delayed_1_0_1306_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => lorx_xlhsx_xfalse135_exec_guard_1297,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => lorx_xlhsx_xfalse135_exec_guard_1207_delayed_1_0_1308,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_lorx_xlhsx_xfalse135_exec_guard_1213_delayed_1_0_1315_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_lorx_xlhsx_xfalse135_exec_guard_1213_delayed_1_0_1315_inst_req_0;
      W_lorx_xlhsx_xfalse135_exec_guard_1213_delayed_1_0_1315_inst_ack_0<= wack(0);
      rreq(0) <= W_lorx_xlhsx_xfalse135_exec_guard_1213_delayed_1_0_1315_inst_req_1;
      W_lorx_xlhsx_xfalse135_exec_guard_1213_delayed_1_0_1315_inst_ack_1<= rack(0);
      W_lorx_xlhsx_xfalse135_exec_guard_1213_delayed_1_0_1315_inst : InterlockBuffer generic map ( -- 
        name => "W_lorx_xlhsx_xfalse135_exec_guard_1213_delayed_1_0_1315_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => lorx_xlhsx_xfalse135_exec_guard_1297,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => lorx_xlhsx_xfalse135_exec_guard_1213_delayed_1_0_1317,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_lorx_xlhsx_xfalse135_exec_guard_1220_delayed_1_0_1325_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_lorx_xlhsx_xfalse135_exec_guard_1220_delayed_1_0_1325_inst_req_0;
      W_lorx_xlhsx_xfalse135_exec_guard_1220_delayed_1_0_1325_inst_ack_0<= wack(0);
      rreq(0) <= W_lorx_xlhsx_xfalse135_exec_guard_1220_delayed_1_0_1325_inst_req_1;
      W_lorx_xlhsx_xfalse135_exec_guard_1220_delayed_1_0_1325_inst_ack_1<= rack(0);
      W_lorx_xlhsx_xfalse135_exec_guard_1220_delayed_1_0_1325_inst : InterlockBuffer generic map ( -- 
        name => "W_lorx_xlhsx_xfalse135_exec_guard_1220_delayed_1_0_1325_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => lorx_xlhsx_xfalse135_exec_guard_1297,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => lorx_xlhsx_xfalse135_exec_guard_1220_delayed_1_0_1327,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_lorx_xlhsx_xfalse135_exec_guard_1228_delayed_1_0_1339_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_lorx_xlhsx_xfalse135_exec_guard_1228_delayed_1_0_1339_inst_req_0;
      W_lorx_xlhsx_xfalse135_exec_guard_1228_delayed_1_0_1339_inst_ack_0<= wack(0);
      rreq(0) <= W_lorx_xlhsx_xfalse135_exec_guard_1228_delayed_1_0_1339_inst_req_1;
      W_lorx_xlhsx_xfalse135_exec_guard_1228_delayed_1_0_1339_inst_ack_1<= rack(0);
      W_lorx_xlhsx_xfalse135_exec_guard_1228_delayed_1_0_1339_inst : InterlockBuffer generic map ( -- 
        name => "W_lorx_xlhsx_xfalse135_exec_guard_1228_delayed_1_0_1339_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => lorx_xlhsx_xfalse135_exec_guard_1297,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => lorx_xlhsx_xfalse135_exec_guard_1228_delayed_1_0_1341,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_lorx_xlhsx_xfalse135_exec_guard_1235_delayed_1_0_1348_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_lorx_xlhsx_xfalse135_exec_guard_1235_delayed_1_0_1348_inst_req_0;
      W_lorx_xlhsx_xfalse135_exec_guard_1235_delayed_1_0_1348_inst_ack_0<= wack(0);
      rreq(0) <= W_lorx_xlhsx_xfalse135_exec_guard_1235_delayed_1_0_1348_inst_req_1;
      W_lorx_xlhsx_xfalse135_exec_guard_1235_delayed_1_0_1348_inst_ack_1<= rack(0);
      W_lorx_xlhsx_xfalse135_exec_guard_1235_delayed_1_0_1348_inst : InterlockBuffer generic map ( -- 
        name => "W_lorx_xlhsx_xfalse135_exec_guard_1235_delayed_1_0_1348_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => lorx_xlhsx_xfalse135_exec_guard_1297,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => lorx_xlhsx_xfalse135_exec_guard_1235_delayed_1_0_1350,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_lorx_xlhsx_xfalse135_exec_guard_1240_delayed_1_0_1356_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_lorx_xlhsx_xfalse135_exec_guard_1240_delayed_1_0_1356_inst_req_0;
      W_lorx_xlhsx_xfalse135_exec_guard_1240_delayed_1_0_1356_inst_ack_0<= wack(0);
      rreq(0) <= W_lorx_xlhsx_xfalse135_exec_guard_1240_delayed_1_0_1356_inst_req_1;
      W_lorx_xlhsx_xfalse135_exec_guard_1240_delayed_1_0_1356_inst_ack_1<= rack(0);
      W_lorx_xlhsx_xfalse135_exec_guard_1240_delayed_1_0_1356_inst : InterlockBuffer generic map ( -- 
        name => "W_lorx_xlhsx_xfalse135_exec_guard_1240_delayed_1_0_1356_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => lorx_xlhsx_xfalse135_exec_guard_1297,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => lorx_xlhsx_xfalse135_exec_guard_1240_delayed_1_0_1358,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock W_lorx_xlhsx_xfalse135_exec_guard_1295_inst
    process(ifx_xend80_lorx_xlhsx_xfalse135_taken_1285) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := ifx_xend80_lorx_xlhsx_xfalse135_taken_1285(0 downto 0);
      lorx_xlhsx_xfalse135_exec_guard_1297 <= tmp_var; -- 
    end process;
    -- interlock W_whilex_xbody_ifx_xelse_taken_935_inst
    process(cmp_934) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := cmp_934(0 downto 0);
      whilex_xbody_ifx_xelse_taken_937 <= tmp_var; -- 
    end process;
    addr_of_1409_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1409_final_reg_req_0;
      addr_of_1409_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1409_final_reg_req_1;
      addr_of_1409_final_reg_ack_1<= rack(0);
      addr_of_1409_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1409_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1408_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_1410,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1456_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1456_final_reg_req_0;
      addr_of_1456_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1456_final_reg_req_1;
      addr_of_1456_final_reg_ack_1<= rack(0);
      addr_of_1456_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1456_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1455_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx160_1457,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1502_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1502_final_reg_req_0;
      addr_of_1502_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1502_final_reg_req_1;
      addr_of_1502_final_reg_ack_1<= rack(0);
      addr_of_1502_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1502_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1501_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx166_1503,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1025_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_1025_inst_req_0;
      type_cast_1025_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_1025_inst_req_1;
      type_cast_1025_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  ifx_xelse_exec_guard_992_delayed_2_0_1021(0);
      type_cast_1025_inst_gI: SplitGuardInterface generic map(name => "type_cast_1025_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_1025_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1025_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc67x_xix_x2_1004,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv69_1026,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1074_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1074_inst_req_0;
      type_cast_1074_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1074_inst_req_1;
      type_cast_1074_inst_ack_1<= rack(0);
      type_cast_1074_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1074_inst",
        buffer_size => 3,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_954,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1030_1030_delayed_3_0_1075,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1098_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1098_inst_req_0;
      type_cast_1098_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1098_inst_req_1;
      type_cast_1098_inst_ack_1<= rack(0);
      type_cast_1098_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1098_inst",
        buffer_size => 4,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ix_x2_910,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1048_1048_delayed_4_0_1099,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1102_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1102_inst_req_0;
      type_cast_1102_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1102_inst_req_1;
      type_cast_1102_inst_ack_1<= rack(0);
      type_cast_1102_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1102_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc67x_xix_x2_1004,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1051_1051_delayed_1_0_1103,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1106_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1106_inst_req_0;
      type_cast_1106_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1106_inst_req_1;
      type_cast_1106_inst_ack_1<= rack(0);
      type_cast_1106_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1106_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc67x_xix_x2_1004,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1054_1054_delayed_1_0_1107,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1126_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1126_inst_req_0;
      type_cast_1126_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1126_inst_req_1;
      type_cast_1126_inst_ack_1<= rack(0);
      type_cast_1126_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1126_inst",
        buffer_size => 4,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x1_915,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1064_1064_delayed_4_0_1127,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1130_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1130_inst_req_0;
      type_cast_1130_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1130_inst_req_1;
      type_cast_1130_inst_ack_1<= rack(0);
      type_cast_1130_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1130_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x2_1018,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1067_1067_delayed_2_0_1131,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1134_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1134_inst_req_0;
      type_cast_1134_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1134_inst_req_1;
      type_cast_1134_inst_ack_1<= rack(0);
      type_cast_1134_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1134_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x2_1018,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1070_1070_delayed_2_0_1135,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1234_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_1234_inst_req_0;
      type_cast_1234_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_1234_inst_req_1;
      type_cast_1234_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  ifx_xend80_exec_guard_1068(0);
      type_cast_1234_inst_gI: SplitGuardInterface generic map(name => "type_cast_1234_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_1234_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1234_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ix_x1_1120,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv121_1235,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1260_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1260_inst_req_0;
      type_cast_1260_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1260_inst_req_1;
      type_cast_1260_inst_ack_1<= rack(0);
      type_cast_1260_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1260_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add132_879,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1179_1179_delayed_1_0_1261,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1265_inst
    process(conv121_1235) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv121_1235(31 downto 0);
      type_cast_1265_wire <= tmp_var; -- 
    end process;
    type_cast_1304_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_1304_inst_req_0;
      type_cast_1304_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_1304_inst_req_1;
      type_cast_1304_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  lorx_xlhsx_xfalse135_exec_guard_1297(0);
      type_cast_1304_inst_gI: SplitGuardInterface generic map(name => "type_cast_1304_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_1304_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1304_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x0_1204_delayed_1_0_1300,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv137_1305,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1330_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1330_inst_req_0;
      type_cast_1330_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1330_inst_req_1;
      type_cast_1330_inst_ack_1<= rack(0);
      type_cast_1330_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1330_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add149_884,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1225_1225_delayed_1_0_1331,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1335_inst
    process(conv137_1305) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv137_1305(31 downto 0);
      type_cast_1335_wire <= tmp_var; -- 
    end process;
    type_cast_1380_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_1380_inst_req_0;
      type_cast_1380_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_1380_inst_req_1;
      type_cast_1380_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  ifx_xthen152_exec_guard_1372(0);
      type_cast_1380_inst_gI: SplitGuardInterface generic map(name => "type_cast_1380_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_1380_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1380_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1379_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv154_1381,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1388_inst
    process(conv154_1381) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv154_1381(31 downto 0);
      type_cast_1388_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1393_inst
    process(ASHR_i32_i32_1392_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1392_wire(31 downto 0);
      shr_1394 <= tmp_var; -- 
    end process;
    type_cast_1402_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_1402_inst_req_0;
      type_cast_1402_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_1402_inst_req_1;
      type_cast_1402_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  ifx_xthen152_exec_guard_1266_delayed_1_0_1397(0);
      type_cast_1402_inst_gI: SplitGuardInterface generic map(name => "type_cast_1402_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_1402_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1402_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1401_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_1403,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1427_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_1427_inst_req_0;
      type_cast_1427_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_1427_inst_req_1;
      type_cast_1427_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  ifx_xelse155_exec_guard_1419(0);
      type_cast_1427_inst_gI: SplitGuardInterface generic map(name => "type_cast_1427_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_1427_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1427_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1426_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv157_1428,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1435_inst
    process(conv157_1428) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv157_1428(31 downto 0);
      type_cast_1435_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1440_inst
    process(ASHR_i32_i32_1439_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1439_wire(31 downto 0);
      shr158_1441 <= tmp_var; -- 
    end process;
    type_cast_1449_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_1449_inst_req_0;
      type_cast_1449_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_1449_inst_req_1;
      type_cast_1449_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  ifx_xelse155_exec_guard_1304_delayed_1_0_1444(0);
      type_cast_1449_inst_gI: SplitGuardInterface generic map(name => "type_cast_1449_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_1449_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1449_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1448_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom159_1450,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1473_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_1473_inst_req_0;
      type_cast_1473_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_1473_inst_req_1;
      type_cast_1473_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  ifx_xelse155_exec_guard_1419(0);
      type_cast_1473_inst_gI: SplitGuardInterface generic map(name => "type_cast_1473_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_1473_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1473_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1472_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv163_1474,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1481_inst
    process(conv163_1474) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv163_1474(31 downto 0);
      type_cast_1481_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1486_inst
    process(ASHR_i32_i32_1485_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1485_wire(31 downto 0);
      shr164_1487 <= tmp_var; -- 
    end process;
    type_cast_1495_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_1495_inst_req_0;
      type_cast_1495_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_1495_inst_req_1;
      type_cast_1495_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  ifx_xelse155_exec_guard_1338_delayed_1_0_1490(0);
      type_cast_1495_inst_gI: SplitGuardInterface generic map(name => "type_cast_1495_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_1495_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1495_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1494_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom165_1496,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_809_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_809_inst_req_0;
      type_cast_809_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_809_inst_req_1;
      type_cast_809_inst_ack_1<= rack(0);
      type_cast_809_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_809_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_792,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv27_810,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_813_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_813_inst_req_0;
      type_cast_813_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_813_inst_req_1;
      type_cast_813_inst_ack_1<= rack(0);
      type_cast_813_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_813_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call1_789,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv29_814,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_817_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_817_inst_req_0;
      type_cast_817_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_817_inst_req_1;
      type_cast_817_inst_ack_1<= rack(0);
      type_cast_817_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_817_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call5_801,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv33_818,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_821_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_821_inst_req_0;
      type_cast_821_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_821_inst_req_1;
      type_cast_821_inst_ack_1<= rack(0);
      type_cast_821_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_821_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call4_798,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv35_822,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_825_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_825_inst_req_0;
      type_cast_825_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_825_inst_req_1;
      type_cast_825_inst_ack_1<= rack(0);
      type_cast_825_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_825_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_792,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv44_826,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_835_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_835_inst_req_0;
      type_cast_835_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_835_inst_req_1;
      type_cast_835_inst_ack_1<= rack(0);
      type_cast_835_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_835_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call1_789,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv58_836,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_839_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_839_inst_req_0;
      type_cast_839_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_839_inst_req_1;
      type_cast_839_inst_ack_1<= rack(0);
      type_cast_839_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_839_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call6_804,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv60_840,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_854_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_854_inst_req_0;
      type_cast_854_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_854_inst_req_1;
      type_cast_854_inst_ack_1<= rack(0);
      type_cast_854_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_854_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_786,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv71_855,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_868_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_868_inst_req_0;
      type_cast_868_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_868_inst_req_1;
      type_cast_868_inst_ack_1<= rack(0);
      type_cast_868_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_868_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call6_804,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv106_869,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_908_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_908_inst_req_0;
      type_cast_908_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_908_inst_req_1;
      type_cast_908_inst_ack_1<= rack(0);
      type_cast_908_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_908_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => kx_x0_1092,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_908_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_913_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_913_inst_req_0;
      type_cast_913_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_913_inst_req_1;
      type_cast_913_inst_ack_1<= rack(0);
      type_cast_913_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_913_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ix_x1_1120,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_913_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_918_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_918_inst_req_0;
      type_cast_918_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_918_inst_req_1;
      type_cast_918_inst_ack_1<= rack(0);
      type_cast_918_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_918_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => jx_x0_1148,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_918_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_923_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_923_inst_req_0;
      type_cast_923_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_923_inst_req_1;
      type_cast_923_inst_ack_1<= rack(0);
      type_cast_923_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_923_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => kx_x1_905,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv47_924,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_927_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_927_inst_req_0;
      type_cast_927_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_927_inst_req_1;
      type_cast_927_inst_ack_1<= rack(0);
      type_cast_927_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_927_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub_832,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_929_929_delayed_2_0_928,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_931_inst
    process(conv47_924) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := conv47_924(31 downto 0);
      type_cast_931_wire <= tmp_var; -- 
    end process;
    type_cast_974_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_974_inst_req_0;
      type_cast_974_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_974_inst_req_1;
      type_cast_974_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  ifx_xelse_exec_guard_960(0);
      type_cast_974_inst_gI: SplitGuardInterface generic map(name => "type_cast_974_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_974_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_974_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc_970,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv56_975,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_991_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_991_inst_req_0;
      type_cast_991_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_991_inst_req_1;
      type_cast_991_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  ifx_xelse_exec_guard_973_delayed_1_0_987(0);
      type_cast_991_inst_gI: SplitGuardInterface generic map(name => "type_cast_991_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_991_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_991_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp62_984,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc67_992,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1408_index_1_rename
    process(R_idxprom_1407_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_1407_resized;
      ov(13 downto 0) := iv;
      R_idxprom_1407_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1408_index_1_resize
    process(idxprom_1403) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_1403;
      ov := iv(13 downto 0);
      R_idxprom_1407_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1408_root_address_inst
    process(array_obj_ref_1408_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1408_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1408_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1455_index_1_rename
    process(R_idxprom159_1454_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom159_1454_resized;
      ov(13 downto 0) := iv;
      R_idxprom159_1454_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1455_index_1_resize
    process(idxprom159_1450) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom159_1450;
      ov := iv(13 downto 0);
      R_idxprom159_1454_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1455_root_address_inst
    process(array_obj_ref_1455_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1455_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1455_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1501_index_1_rename
    process(R_idxprom165_1500_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom165_1500_resized;
      ov(13 downto 0) := iv;
      R_idxprom165_1500_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1501_index_1_resize
    process(idxprom165_1496) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom165_1496;
      ov := iv(13 downto 0);
      R_idxprom165_1500_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1501_root_address_inst
    process(array_obj_ref_1501_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1501_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1501_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1413_addr_0
    process(ptr_deref_1413_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1413_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1413_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1413_base_resize
    process(arrayidx_1410) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_1410;
      ov := iv(13 downto 0);
      ptr_deref_1413_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1413_gather_scatter
    process(type_cast_1415_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_1415_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_1413_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1413_root_address_inst
    process(ptr_deref_1413_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1413_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1413_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1464_addr_0
    process(ptr_deref_1464_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1464_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1464_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1464_base_resize
    process(arrayidx160_1457) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx160_1457;
      ov := iv(13 downto 0);
      ptr_deref_1464_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1464_gather_scatter
    process(ptr_deref_1464_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1464_data_0;
      ov(63 downto 0) := iv;
      tmp161_1465 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1464_root_address_inst
    process(ptr_deref_1464_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1464_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1464_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1512_addr_0
    process(ptr_deref_1512_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1512_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1512_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1512_base_resize
    process(arrayidx166_1352_delayed_6_0_1509) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx166_1352_delayed_6_0_1509;
      ov := iv(13 downto 0);
      ptr_deref_1512_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1512_gather_scatter
    process(tmp161_1465) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp161_1465;
      ov(63 downto 0) := iv;
      ptr_deref_1512_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1512_root_address_inst
    process(ptr_deref_1512_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1512_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1512_root_address <= ov(13 downto 0);
      --
    end process;
    do_while_stmt_903_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tobool_1520;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_903_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_903_branch_req_0,
          ack0 => do_while_stmt_903_branch_ack_0,
          ack1 => do_while_stmt_903_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1527_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= ifx_xend167_whilex_xend_taken_1524;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1527_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1527_branch_req_0,
          ack0 => if_stmt_1527_branch_ack_0,
          ack1 => if_stmt_1527_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1003_inst
    process(inc67_992, ix_x2_981_delayed_3_0_998) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc67_992, ix_x2_981_delayed_3_0_998, tmp_var);
      inc67x_xix_x2_1004 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1187_inst
    process(mul95_1182, kx_x0_1092) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul95_1182, kx_x0_1092, tmp_var);
      add90_1188 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1193_inst
    process(add90_1188, mul89_1176) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add90_1188, mul89_1176, tmp_var);
      add96_1194 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1223_inst
    process(mul117_1218, kx_x0_1092) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul117_1218, kx_x0_1092, tmp_var);
      add109_1224 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1229_inst
    process(add109_1224, mul108_1206) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add109_1224, mul108_1206, tmp_var);
      add118_1230 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_953_inst
    process(kx_x1_944_delayed_1_0_947) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(kx_x1_944_delayed_1_0_947, type_cast_952_wire_constant, tmp_var);
      add_954 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_969_inst
    process(jx_x1_957_delayed_1_0_963) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(jx_x1_957_delayed_1_0_963, type_cast_968_wire_constant, tmp_var);
      inc_970 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_831_inst
    process(conv44_826) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv44_826, type_cast_830_wire_constant, tmp_var);
      sub_832 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_850_inst
    process(shl_846, conv58_836) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shl_846, conv58_836, tmp_var);
      add61_851 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_859_inst
    process(shl_846, conv71_855) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shl_846, conv71_855, tmp_var);
      add75_860 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_878_inst
    process(conv60_840, conv71_855) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv60_840, conv71_855, tmp_var);
      add132_879 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_883_inst
    process(conv60_840, conv58_836) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv60_840, conv58_836, tmp_var);
      add149_884 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1042_inst
    process(ifx_xelse_exec_guard_1004_delayed_3_0_1038, cmp76_1035) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(ifx_xelse_exec_guard_1004_delayed_3_0_1038, cmp76_1035, tmp_var);
      ifx_xelse_ifx_xthen78_taken_1043 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1051_inst
    process(ifx_xelse_exec_guard_1009_delayed_3_0_1046, NOT_u1_u1_1050_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(ifx_xelse_exec_guard_1009_delayed_3_0_1046, NOT_u1_u1_1050_wire, tmp_var);
      ifx_xelse_ifx_xend80_taken_1052 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1276_inst
    process(cmp124x_xnot_1254, cmp133_1268) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(cmp124x_xnot_1254, cmp133_1268, tmp_var);
      orx_xcond_1277 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1284_inst
    process(ifx_xend80_exec_guard_1189_delayed_1_0_1280, orx_xcond_1277) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(ifx_xend80_exec_guard_1189_delayed_1_0_1280, orx_xcond_1277, tmp_var);
      ifx_xend80_lorx_xlhsx_xfalse135_taken_1285 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1293_inst
    process(ifx_xend80_exec_guard_1194_delayed_1_0_1288, NOT_u1_u1_1292_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(ifx_xend80_exec_guard_1194_delayed_1_0_1288, NOT_u1_u1_1292_wire, tmp_var);
      ifx_xend80_ifx_xthen152_taken_1294 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1346_inst
    process(cmp140x_xnot_1324, cmp150_1338) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(cmp140x_xnot_1324, cmp150_1338, tmp_var);
      orx_xcond171_1347 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1354_inst
    process(lorx_xlhsx_xfalse135_exec_guard_1235_delayed_1_0_1350, orx_xcond171_1347) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(lorx_xlhsx_xfalse135_exec_guard_1235_delayed_1_0_1350, orx_xcond171_1347, tmp_var);
      lorx_xlhsx_xfalse135_ifx_xelse155_taken_1355 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1363_inst
    process(lorx_xlhsx_xfalse135_exec_guard_1240_delayed_1_0_1358, NOT_u1_u1_1362_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(lorx_xlhsx_xfalse135_exec_guard_1240_delayed_1_0_1358, NOT_u1_u1_1362_wire, tmp_var);
      lorx_xlhsx_xfalse135_ifx_xthen152_taken_1364 <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1392_inst
    process(type_cast_1388_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1388_wire, type_cast_1391_wire_constant, tmp_var);
      ASHR_i32_i32_1392_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1439_inst
    process(type_cast_1435_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1435_wire, type_cast_1438_wire_constant, tmp_var);
      ASHR_i32_i32_1439_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1485_inst
    process(type_cast_1481_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1481_wire, type_cast_1484_wire_constant, tmp_var);
      ASHR_i32_i32_1485_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_1519_inst
    process(flagx_x0_1170) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(flagx_x0_1170, type_cast_1518_wire_constant, tmp_var);
      tobool_1520 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1034_inst
    process(conv69_1026, add75_860) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv69_1026, add75_860, tmp_var);
      cmp76_1035 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_983_inst
    process(conv56_975, add61_851) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv56_975, add61_851, tmp_var);
      cmp62_984 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1175_inst
    process(jx_x0_1148, conv33_818) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(jx_x0_1148, conv33_818, tmp_var);
      mul89_1176 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1181_inst
    process(mul36_865, ix_x1_1120) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul36_865, ix_x1_1120, tmp_var);
      mul95_1182 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1205_inst
    process(sub107_1200, conv27_810) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(sub107_1200, conv27_810, tmp_var);
      mul108_1206 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1217_inst
    process(mul_874, sub116_1212) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_874, sub116_1212, tmp_var);
      mul117_1218 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_864_inst
    process(conv33_818, conv35_822) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv33_818, conv35_822, tmp_var);
      mul36_865 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_873_inst
    process(conv27_810, conv29_814) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv27_810, conv29_814, tmp_var);
      mul_874 <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_1050_inst
    process(cmp76_1035) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", cmp76_1035, tmp_var);
      NOT_u1_u1_1050_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1292_inst
    process(orx_xcond_1277) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", orx_xcond_1277, tmp_var);
      NOT_u1_u1_1292_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1362_inst
    process(orx_xcond171_1347) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", orx_xcond171_1347, tmp_var);
      NOT_u1_u1_1362_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1523_inst
    process(tobool_1520) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", tobool_1520, tmp_var);
      ifx_xend167_whilex_xend_taken_1524 <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_940_inst
    process(cmp_934) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", cmp_934, tmp_var);
      whilex_xbody_ifx_xthen_taken_941 <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_1066_inst
    process(ifx_xthen_ifx_xend80_taken_1022_delayed_3_0_1061, ifx_xthen78_ifx_xend80_taken_1058) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(ifx_xthen_ifx_xend80_taken_1022_delayed_3_0_1061, ifx_xthen78_ifx_xend80_taken_1058, tmp_var);
      OR_u1_u1_1066_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1067_inst
    process(ifx_xelse_ifx_xend80_taken_1052, OR_u1_u1_1066_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(ifx_xelse_ifx_xend80_taken_1052, OR_u1_u1_1066_wire, tmp_var);
      ifx_xend80_exec_guard_1068 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1371_inst
    process(ifx_xend80_ifx_xthen152_taken_1246_delayed_1_0_1367, lorx_xlhsx_xfalse135_ifx_xthen152_taken_1364) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(ifx_xend80_ifx_xthen152_taken_1246_delayed_1_0_1367, lorx_xlhsx_xfalse135_ifx_xthen152_taken_1364, tmp_var);
      ifx_xthen152_exec_guard_1372 <= tmp_var; --
    end process;
    -- binary operator SGT_i32_u1_933_inst
    process(type_cast_931_wire, type_cast_929_929_delayed_2_0_928) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(type_cast_931_wire, type_cast_929_929_delayed_2_0_928, tmp_var);
      cmp_934 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_845_inst
    process(conv60_840) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv60_840, type_cast_844_wire_constant, tmp_var);
      shl_846 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1267_inst
    process(type_cast_1265_wire, type_cast_1179_1179_delayed_1_0_1261) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1265_wire, type_cast_1179_1179_delayed_1_0_1261, tmp_var);
      cmp133_1268 <= tmp_var; --
    end process;
    -- binary operator SLT_i32_u1_1337_inst
    process(type_cast_1335_wire, type_cast_1225_1225_delayed_1_0_1331) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSlt_proc(type_cast_1335_wire, type_cast_1225_1225_delayed_1_0_1331, tmp_var);
      cmp150_1338 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1199_inst
    process(jx_x0_1148, conv106_869) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(jx_x0_1148, conv106_869, tmp_var);
      sub107_1200 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_1211_inst
    process(ix_x1_1120, conv106_869) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(ix_x1_1120, conv106_869, tmp_var);
      sub116_1212 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_1243_inst
    process(conv121_1235, conv60_840) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(conv121_1235, conv60_840, tmp_var);
      cmp124_1244 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_1313_inst
    process(conv137_1305, conv60_840) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(conv137_1305, conv60_840, tmp_var);
      cmp140_1314 <= tmp_var; --
    end process;
    -- binary operator XOR_u1_u1_1253_inst
    process(cmp124_1244) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntXor_proc(cmp124_1244, type_cast_1252_wire_constant, tmp_var);
      cmp124x_xnot_1254 <= tmp_var; --
    end process;
    -- binary operator XOR_u1_u1_1323_inst
    process(cmp140_1314) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntXor_proc(cmp140_1314, type_cast_1322_wire_constant, tmp_var);
      cmp140x_xnot_1324 <= tmp_var; --
    end process;
    -- shared split operator group (50) : array_obj_ref_1408_index_offset 
    ApIntAdd_group_50: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_1407_scaled;
      array_obj_ref_1408_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1408_index_offset_req_0;
      array_obj_ref_1408_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1408_index_offset_req_1;
      array_obj_ref_1408_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_50_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_50_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_50",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 50
    -- shared split operator group (51) : array_obj_ref_1455_index_offset 
    ApIntAdd_group_51: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom159_1454_scaled;
      array_obj_ref_1455_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1455_index_offset_req_0;
      array_obj_ref_1455_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1455_index_offset_req_1;
      array_obj_ref_1455_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_51_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_51_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_51",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 51
    -- shared split operator group (52) : array_obj_ref_1501_index_offset 
    ApIntAdd_group_52: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom165_1500_scaled;
      array_obj_ref_1501_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1501_index_offset_req_0;
      array_obj_ref_1501_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1501_index_offset_req_1;
      array_obj_ref_1501_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_52_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_52_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_52",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 52
    -- unary operator type_cast_1379_inst
    process(add96_1252_delayed_2_0_1375) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", add96_1252_delayed_2_0_1375, tmp_var);
      type_cast_1379_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1401_inst
    process(shr_1394) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr_1394, tmp_var);
      type_cast_1401_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1426_inst
    process(add118_1290_delayed_2_0_1422) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", add118_1290_delayed_2_0_1422, tmp_var);
      type_cast_1426_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1448_inst
    process(shr158_1441) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr158_1441, tmp_var);
      type_cast_1448_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1472_inst
    process(add96_1324_delayed_2_0_1468) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", add96_1324_delayed_2_0_1468, tmp_var);
      type_cast_1472_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1494_inst
    process(shr164_1487) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr164_1487, tmp_var);
      type_cast_1494_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : ptr_deref_1464_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 6);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1464_load_0_req_0;
      ptr_deref_1464_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1464_load_0_req_1;
      ptr_deref_1464_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= ifx_xelse155_exec_guard_1317_delayed_9_0_1460(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1464_word_address_0;
      ptr_deref_1464_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_1413_store_0 ptr_deref_1512_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(27 downto 0);
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 2, 0 => 2);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 15, 0 => 15);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => true, 1 => true);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 6, 1 => 6);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1413_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1512_store_0_req_0;
      ptr_deref_1413_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1512_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1413_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1512_store_0_req_1;
      ptr_deref_1413_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1512_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= ifx_xelse155_exec_guard_1351_delayed_15_0_1506(0);
      guard_vector(1)  <= ifx_xthen152_exec_guard_1372(0);
      StoreGroup0_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1413_word_address_0 & ptr_deref_1512_word_address_0;
      data_in <= ptr_deref_1413_data_0 & ptr_deref_1512_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(13 downto 0),
          mdata => memory_space_0_sr_data(63 downto 0),
          mtag => memory_space_0_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block0_starting_785_inst RPIPE_Block0_starting_788_inst RPIPE_Block0_starting_791_inst RPIPE_Block0_starting_794_inst RPIPE_Block0_starting_797_inst RPIPE_Block0_starting_800_inst RPIPE_Block0_starting_803_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(55 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 6 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 6 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 6 downto 0);
      signal guard_vector : std_logic_vector( 6 downto 0);
      constant outBUFs : IntegerArray(6 downto 0) := (6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(6 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false);
      constant guardBuffering: IntegerArray(6 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2);
      -- 
    begin -- 
      reqL_unguarded(6) <= RPIPE_Block0_starting_785_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Block0_starting_788_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Block0_starting_791_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Block0_starting_794_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Block0_starting_797_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Block0_starting_800_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Block0_starting_803_inst_req_0;
      RPIPE_Block0_starting_785_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Block0_starting_788_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Block0_starting_791_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Block0_starting_794_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Block0_starting_797_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Block0_starting_800_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Block0_starting_803_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(6) <= RPIPE_Block0_starting_785_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Block0_starting_788_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Block0_starting_791_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Block0_starting_794_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Block0_starting_797_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Block0_starting_800_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Block0_starting_803_inst_req_1;
      RPIPE_Block0_starting_785_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Block0_starting_788_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Block0_starting_791_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Block0_starting_794_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Block0_starting_797_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Block0_starting_800_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Block0_starting_803_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      call_786 <= data_out(55 downto 48);
      call1_789 <= data_out(47 downto 40);
      call2_792 <= data_out(39 downto 32);
      call3_795 <= data_out(31 downto 24);
      call4_798 <= data_out(23 downto 16);
      call5_801 <= data_out(15 downto 8);
      call6_804 <= data_out(7 downto 0);
      Block0_starting_read_0_gI: SplitGuardInterface generic map(name => "Block0_starting_read_0_gI", nreqs => 7, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block0_starting_read_0: InputPortRevised -- 
        generic map ( name => "Block0_starting_read_0", data_width => 8,  num_reqs => 7,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block0_starting_pipe_read_req(0),
          oack => Block0_starting_pipe_read_ack(0),
          odata => Block0_starting_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block0_complete_1533_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block0_complete_1533_inst_req_0;
      WPIPE_Block0_complete_1533_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block0_complete_1533_inst_req_1;
      WPIPE_Block0_complete_1533_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_1535_wire_constant;
      Block0_complete_write_0_gI: SplitGuardInterface generic map(name => "Block0_complete_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block0_complete_write_0: OutputPortRevised -- 
        generic map ( name => "Block0_complete", data_width => 8, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block0_complete_pipe_write_req(0),
          oack => Block0_complete_pipe_write_ack(0),
          odata => Block0_complete_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end zeropad3D_A_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    zeropad_input_pipe_pipe_write_data: in std_logic_vector(7 downto 0);
    zeropad_input_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    zeropad_input_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    zeropad_output_pipe_pipe_read_data: out std_logic_vector(7 downto 0);
    zeropad_output_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    zeropad_output_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(18 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(1 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(17 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(17 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_2_lr_tag : std_logic_vector(0 downto 0);
  signal memory_space_2_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_2_lc_tag :  std_logic_vector(0 downto 0);
  -- declarations related to module sendOutput
  component sendOutput is -- 
    generic (tag_length : integer); 
    port ( -- 
      size : in  std_logic_vector(31 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
      zeropad_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      zeropad_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      zeropad_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module sendOutput
  signal sendOutput_size :  std_logic_vector(31 downto 0);
  signal sendOutput_in_args    : std_logic_vector(31 downto 0);
  signal sendOutput_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal sendOutput_tag_out   : std_logic_vector(1 downto 0);
  signal sendOutput_start_req : std_logic;
  signal sendOutput_start_ack : std_logic;
  signal sendOutput_fin_req   : std_logic;
  signal sendOutput_fin_ack : std_logic;
  -- caller side aggregated signals for module sendOutput
  signal sendOutput_call_reqs: std_logic_vector(0 downto 0);
  signal sendOutput_call_acks: std_logic_vector(0 downto 0);
  signal sendOutput_return_reqs: std_logic_vector(0 downto 0);
  signal sendOutput_return_acks: std_logic_vector(0 downto 0);
  signal sendOutput_call_data: std_logic_vector(31 downto 0);
  signal sendOutput_call_tag: std_logic_vector(0 downto 0);
  signal sendOutput_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module timer
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      c : out  std_logic_vector(63 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timer
  signal timer_c :  std_logic_vector(63 downto 0);
  signal timer_out_args   : std_logic_vector(63 downto 0);
  signal timer_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal timer_tag_out   : std_logic_vector(2 downto 0);
  signal timer_start_req : std_logic;
  signal timer_start_ack : std_logic;
  signal timer_fin_req   : std_logic;
  signal timer_fin_ack : std_logic;
  -- caller side aggregated signals for module timer
  signal timer_call_reqs: std_logic_vector(0 downto 0);
  signal timer_call_acks: std_logic_vector(0 downto 0);
  signal timer_return_reqs: std_logic_vector(0 downto 0);
  signal timer_return_acks: std_logic_vector(0 downto 0);
  signal timer_call_tag: std_logic_vector(1 downto 0);
  signal timer_return_data: std_logic_vector(63 downto 0);
  signal timer_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module zeropad3D
  component zeropad3D is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
      Block0_complete_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block0_complete_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block0_complete_pipe_read_data : in   std_logic_vector(7 downto 0);
      zeropad_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      zeropad_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      zeropad_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      zeropad_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      zeropad_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      zeropad_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      Block0_starting_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block0_starting_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block0_starting_pipe_write_data : out  std_logic_vector(7 downto 0);
      sendOutput_call_reqs : out  std_logic_vector(0 downto 0);
      sendOutput_call_acks : in   std_logic_vector(0 downto 0);
      sendOutput_call_data : out  std_logic_vector(31 downto 0);
      sendOutput_call_tag  :  out  std_logic_vector(0 downto 0);
      sendOutput_return_reqs : out  std_logic_vector(0 downto 0);
      sendOutput_return_acks : in   std_logic_vector(0 downto 0);
      sendOutput_return_tag :  in   std_logic_vector(0 downto 0);
      timer_call_reqs : out  std_logic_vector(0 downto 0);
      timer_call_acks : in   std_logic_vector(0 downto 0);
      timer_call_tag  :  out  std_logic_vector(1 downto 0);
      timer_return_reqs : out  std_logic_vector(0 downto 0);
      timer_return_acks : in   std_logic_vector(0 downto 0);
      timer_return_data : in   std_logic_vector(63 downto 0);
      timer_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module zeropad3D
  signal zeropad3D_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal zeropad3D_tag_out   : std_logic_vector(1 downto 0);
  signal zeropad3D_start_req : std_logic;
  signal zeropad3D_start_ack : std_logic;
  signal zeropad3D_fin_req   : std_logic;
  signal zeropad3D_fin_ack : std_logic;
  -- declarations related to module zeropad3D_A
  component zeropad3D_A is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
      Block0_starting_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block0_starting_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block0_starting_pipe_read_data : in   std_logic_vector(7 downto 0);
      Block0_complete_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block0_complete_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block0_complete_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module zeropad3D_A
  signal zeropad3D_A_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal zeropad3D_A_tag_out   : std_logic_vector(1 downto 0);
  signal zeropad3D_A_start_req : std_logic;
  signal zeropad3D_A_start_ack : std_logic;
  signal zeropad3D_A_fin_req   : std_logic;
  signal zeropad3D_A_fin_ack : std_logic;
  -- aggregate signals for write to pipe Block0_complete
  signal Block0_complete_pipe_write_data: std_logic_vector(7 downto 0);
  signal Block0_complete_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block0_complete_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block0_complete
  signal Block0_complete_pipe_read_data: std_logic_vector(7 downto 0);
  signal Block0_complete_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block0_complete_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block0_starting
  signal Block0_starting_pipe_write_data: std_logic_vector(7 downto 0);
  signal Block0_starting_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block0_starting_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block0_starting
  signal Block0_starting_pipe_read_data: std_logic_vector(7 downto 0);
  signal Block0_starting_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block0_starting_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe zeropad_input_pipe
  signal zeropad_input_pipe_pipe_read_data: std_logic_vector(7 downto 0);
  signal zeropad_input_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal zeropad_input_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe zeropad_output_pipe
  signal zeropad_output_pipe_pipe_write_data: std_logic_vector(15 downto 0);
  signal zeropad_output_pipe_pipe_write_req: std_logic_vector(1 downto 0);
  signal zeropad_output_pipe_pipe_write_ack: std_logic_vector(1 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module sendOutput
  sendOutput_size <= sendOutput_in_args(31 downto 0);
  -- call arbiter for module sendOutput
  sendOutput_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 32,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => sendOutput_call_reqs,
      call_acks => sendOutput_call_acks,
      return_reqs => sendOutput_return_reqs,
      return_acks => sendOutput_return_acks,
      call_data  => sendOutput_call_data,
      call_tag  => sendOutput_call_tag,
      return_tag  => sendOutput_return_tag,
      call_mtag => sendOutput_tag_in,
      return_mtag => sendOutput_tag_out,
      call_mreq => sendOutput_start_req,
      call_mack => sendOutput_start_ack,
      return_mreq => sendOutput_fin_req,
      return_mack => sendOutput_fin_ack,
      call_mdata => sendOutput_in_args,
      clk => clk, 
      reset => reset --
    ); --
  sendOutput_instance:sendOutput-- 
    generic map(tag_length => 2)
    port map(-- 
      size => sendOutput_size,
      start_req => sendOutput_start_req,
      start_ack => sendOutput_start_ack,
      fin_req => sendOutput_fin_req,
      fin_ack => sendOutput_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(13 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(18 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(1 downto 0),
      zeropad_output_pipe_pipe_write_req => zeropad_output_pipe_pipe_write_req(1 downto 1),
      zeropad_output_pipe_pipe_write_ack => zeropad_output_pipe_pipe_write_ack(1 downto 1),
      zeropad_output_pipe_pipe_write_data => zeropad_output_pipe_pipe_write_data(15 downto 8),
      tag_in => sendOutput_tag_in,
      tag_out => sendOutput_tag_out-- 
    ); -- 
  -- module timer
  timer_out_args <= timer_c ;
  -- call arbiter for module timer
  timer_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargs", num_reqs => 1,
      return_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => timer_call_reqs,
      call_acks => timer_call_acks,
      return_reqs => timer_return_reqs,
      return_acks => timer_return_acks,
      call_tag  => timer_call_tag,
      return_tag  => timer_return_tag,
      call_mtag => timer_tag_in,
      return_mtag => timer_tag_out,
      return_data =>timer_return_data,
      call_mreq => timer_start_req,
      call_mack => timer_start_ack,
      return_mreq => timer_fin_req,
      return_mack => timer_fin_ack,
      return_mdata => timer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  timer_instance:timer-- 
    generic map(tag_length => 3)
    port map(-- 
      c => timer_c,
      start_req => timer_start_req,
      start_ack => timer_start_ack,
      fin_req => timer_fin_req,
      fin_ack => timer_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_2_lr_req => memory_space_2_lr_req(0 downto 0),
      memory_space_2_lr_ack => memory_space_2_lr_ack(0 downto 0),
      memory_space_2_lr_addr => memory_space_2_lr_addr(0 downto 0),
      memory_space_2_lr_tag => memory_space_2_lr_tag(0 downto 0),
      memory_space_2_lc_req => memory_space_2_lc_req(0 downto 0),
      memory_space_2_lc_ack => memory_space_2_lc_ack(0 downto 0),
      memory_space_2_lc_data => memory_space_2_lc_data(63 downto 0),
      memory_space_2_lc_tag => memory_space_2_lc_tag(0 downto 0),
      tag_in => timer_tag_in,
      tag_out => timer_tag_out-- 
    ); -- 
  -- module zeropad3D
  zeropad3D_instance:zeropad3D-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => zeropad3D_start_req,
      start_ack => zeropad3D_start_ack,
      fin_req => zeropad3D_fin_req,
      fin_ack => zeropad3D_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(13 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(63 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(17 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(0 downto 0),
      Block0_complete_pipe_read_req => Block0_complete_pipe_read_req(0 downto 0),
      Block0_complete_pipe_read_ack => Block0_complete_pipe_read_ack(0 downto 0),
      Block0_complete_pipe_read_data => Block0_complete_pipe_read_data(7 downto 0),
      zeropad_input_pipe_pipe_read_req => zeropad_input_pipe_pipe_read_req(0 downto 0),
      zeropad_input_pipe_pipe_read_ack => zeropad_input_pipe_pipe_read_ack(0 downto 0),
      zeropad_input_pipe_pipe_read_data => zeropad_input_pipe_pipe_read_data(7 downto 0),
      zeropad_output_pipe_pipe_write_req => zeropad_output_pipe_pipe_write_req(0 downto 0),
      zeropad_output_pipe_pipe_write_ack => zeropad_output_pipe_pipe_write_ack(0 downto 0),
      zeropad_output_pipe_pipe_write_data => zeropad_output_pipe_pipe_write_data(7 downto 0),
      Block0_starting_pipe_write_req => Block0_starting_pipe_write_req(0 downto 0),
      Block0_starting_pipe_write_ack => Block0_starting_pipe_write_ack(0 downto 0),
      Block0_starting_pipe_write_data => Block0_starting_pipe_write_data(7 downto 0),
      sendOutput_call_reqs => sendOutput_call_reqs(0 downto 0),
      sendOutput_call_acks => sendOutput_call_acks(0 downto 0),
      sendOutput_call_data => sendOutput_call_data(31 downto 0),
      sendOutput_call_tag => sendOutput_call_tag(0 downto 0),
      sendOutput_return_reqs => sendOutput_return_reqs(0 downto 0),
      sendOutput_return_acks => sendOutput_return_acks(0 downto 0),
      sendOutput_return_tag => sendOutput_return_tag(0 downto 0),
      timer_call_reqs => timer_call_reqs(0 downto 0),
      timer_call_acks => timer_call_acks(0 downto 0),
      timer_call_tag => timer_call_tag(1 downto 0),
      timer_return_reqs => timer_return_reqs(0 downto 0),
      timer_return_acks => timer_return_acks(0 downto 0),
      timer_return_data => timer_return_data(63 downto 0),
      timer_return_tag => timer_return_tag(1 downto 0),
      tag_in => zeropad3D_tag_in,
      tag_out => zeropad3D_tag_out-- 
    ); -- 
  -- module will be run forever 
  zeropad3D_tag_in <= (others => '0');
  zeropad3D_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => zeropad3D_start_req, start_ack => zeropad3D_start_ack,  fin_req => zeropad3D_fin_req,  fin_ack => zeropad3D_fin_ack);
  -- module zeropad3D_A
  zeropad3D_A_instance:zeropad3D_A-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => zeropad3D_A_start_req,
      start_ack => zeropad3D_A_start_ack,
      fin_req => zeropad3D_A_fin_req,
      fin_ack => zeropad3D_A_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(13 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(17 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(63 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(0 downto 0),
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(13 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(63 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(18 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(1 downto 0),
      Block0_starting_pipe_read_req => Block0_starting_pipe_read_req(0 downto 0),
      Block0_starting_pipe_read_ack => Block0_starting_pipe_read_ack(0 downto 0),
      Block0_starting_pipe_read_data => Block0_starting_pipe_read_data(7 downto 0),
      Block0_complete_pipe_write_req => Block0_complete_pipe_write_req(0 downto 0),
      Block0_complete_pipe_write_ack => Block0_complete_pipe_write_ack(0 downto 0),
      Block0_complete_pipe_write_data => Block0_complete_pipe_write_data(7 downto 0),
      tag_in => zeropad3D_A_tag_in,
      tag_out => zeropad3D_A_tag_out-- 
    ); -- 
  -- module will be run forever 
  zeropad3D_A_tag_in <= (others => '0');
  zeropad3D_A_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => zeropad3D_A_start_req, start_ack => zeropad3D_A_start_ack,  fin_req => zeropad3D_A_fin_req,  fin_ack => zeropad3D_A_fin_ack);
  Block0_complete_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block0_complete",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block0_complete_pipe_read_req,
      read_ack => Block0_complete_pipe_read_ack,
      read_data => Block0_complete_pipe_read_data,
      write_req => Block0_complete_pipe_write_req,
      write_ack => Block0_complete_pipe_write_ack,
      write_data => Block0_complete_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block0_starting_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block0_starting",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block0_starting_pipe_read_req,
      read_ack => Block0_starting_pipe_read_ack,
      read_data => Block0_starting_pipe_read_data,
      write_req => Block0_starting_pipe_write_req,
      write_ack => Block0_starting_pipe_write_ack,
      write_data => Block0_starting_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  zeropad_input_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe zeropad_input_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => zeropad_input_pipe_pipe_read_req,
      read_ack => zeropad_input_pipe_pipe_read_ack,
      read_data => zeropad_input_pipe_pipe_read_data,
      write_req => zeropad_input_pipe_pipe_write_req,
      write_ack => zeropad_input_pipe_pipe_write_ack,
      write_data => zeropad_input_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  zeropad_output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe zeropad_output_pipe",
      num_reads => 1,
      num_writes => 2,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => zeropad_output_pipe_pipe_read_req,
      read_ack => zeropad_output_pipe_pipe_read_ack,
      read_data => zeropad_output_pipe_pipe_read_data,
      write_req => zeropad_output_pipe_pipe_write_req,
      write_ack => zeropad_output_pipe_pipe_write_ack,
      write_data => zeropad_output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  MemorySpace_memory_space_0: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 2,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_1: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  dummyROM_memory_space_2: dummy_read_only_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_2",
      num_loads => 1,
      addr_width => 1,
      data_width => 64,
      tag_width => 1
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_2_lr_addr,
      lr_req_in => memory_space_2_lr_req,
      lr_ack_out => memory_space_2_lr_ack,
      lr_tag_in => memory_space_2_lr_tag,
      lc_req_in => memory_space_2_lc_req,
      lc_ack_out => memory_space_2_lc_ack,
      lc_data_out => memory_space_2_lc_data,
      lc_tag_out => memory_space_2_lc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
