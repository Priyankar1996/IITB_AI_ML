-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity concat is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(15 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(15 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
    Concat_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    Concat_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Concat_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    Concat_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    Concat_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Concat_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    timer_call_reqs : out  std_logic_vector(0 downto 0);
    timer_call_acks : in   std_logic_vector(0 downto 0);
    timer_call_tag  :  out  std_logic_vector(1 downto 0);
    timer_return_reqs : out  std_logic_vector(0 downto 0);
    timer_return_acks : in   std_logic_vector(0 downto 0);
    timer_return_data : in   std_logic_vector(63 downto 0);
    timer_return_tag :  in   std_logic_vector(1 downto 0);
    concat_core_call_reqs : out  std_logic_vector(0 downto 0);
    concat_core_call_acks : in   std_logic_vector(0 downto 0);
    concat_core_call_data : out  std_logic_vector(63 downto 0);
    concat_core_call_tag  :  out  std_logic_vector(0 downto 0);
    concat_core_return_reqs : out  std_logic_vector(0 downto 0);
    concat_core_return_acks : in   std_logic_vector(0 downto 0);
    concat_core_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity concat;
architecture concat_arch of concat is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal concat_CP_664_start: Boolean;
  signal concat_CP_664_symbol: Boolean;
  -- volatile/operator module components. 
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      T : out  std_logic_vector(63 downto 0);
      timer_resp_pipe_read_req : out  std_logic_vector(0 downto 0);
      timer_resp_pipe_read_ack : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_read_data : in   std_logic_vector(63 downto 0);
      timer_req_pipe_write_req : out  std_logic_vector(0 downto 0);
      timer_req_pipe_write_ack : in   std_logic_vector(0 downto 0);
      timer_req_pipe_write_data : out  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component concat_core is -- 
    generic (tag_length : integer); 
    port ( -- 
      input1_count : in  std_logic_vector(15 downto 0);
      input2_count : in  std_logic_vector(15 downto 0);
      output_size : in  std_logic_vector(31 downto 0);
      readModule1_call_reqs : out  std_logic_vector(0 downto 0);
      readModule1_call_acks : in   std_logic_vector(0 downto 0);
      readModule1_call_data : out  std_logic_vector(39 downto 0);
      readModule1_call_tag  :  out  std_logic_vector(1 downto 0);
      readModule1_return_reqs : out  std_logic_vector(0 downto 0);
      readModule1_return_acks : in   std_logic_vector(0 downto 0);
      readModule1_return_data : in   std_logic_vector(63 downto 0);
      readModule1_return_tag :  in   std_logic_vector(1 downto 0);
      writeModule1_call_reqs : out  std_logic_vector(0 downto 0);
      writeModule1_call_acks : in   std_logic_vector(0 downto 0);
      writeModule1_call_data : out  std_logic_vector(103 downto 0);
      writeModule1_call_tag  :  out  std_logic_vector(0 downto 0);
      writeModule1_return_reqs : out  std_logic_vector(0 downto 0);
      writeModule1_return_acks : in   std_logic_vector(0 downto 0);
      writeModule1_return_data : in   std_logic_vector(0 downto 0);
      writeModule1_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal RPIPE_Concat_input_pipe_640_inst_req_0 : boolean;
  signal type_cast_1179_inst_req_0 : boolean;
  signal type_cast_458_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_573_inst_ack_0 : boolean;
  signal type_cast_644_inst_ack_0 : boolean;
  signal type_cast_577_inst_req_1 : boolean;
  signal type_cast_680_inst_req_1 : boolean;
  signal array_obj_ref_1120_index_offset_req_0 : boolean;
  signal addr_of_1121_final_reg_req_0 : boolean;
  signal type_cast_1139_inst_req_0 : boolean;
  signal WPIPE_Concat_output_pipe_1049_inst_req_0 : boolean;
  signal type_cast_1169_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_573_inst_req_1 : boolean;
  signal array_obj_ref_569_index_offset_ack_0 : boolean;
  signal type_cast_698_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_622_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_676_inst_req_0 : boolean;
  signal type_cast_527_inst_req_0 : boolean;
  signal ptr_deref_706_store_0_ack_0 : boolean;
  signal type_cast_680_inst_ack_1 : boolean;
  signal ptr_deref_706_store_0_req_0 : boolean;
  signal type_cast_1139_inst_ack_1 : boolean;
  signal type_cast_1169_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_658_inst_req_1 : boolean;
  signal type_cast_698_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_218_inst_req_0 : boolean;
  signal WPIPE_Concat_output_pipe_1049_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_218_inst_ack_0 : boolean;
  signal type_cast_222_inst_req_0 : boolean;
  signal type_cast_608_inst_ack_0 : boolean;
  signal type_cast_458_inst_req_0 : boolean;
  signal type_cast_458_inst_req_1 : boolean;
  signal type_cast_222_inst_ack_0 : boolean;
  signal type_cast_222_inst_req_1 : boolean;
  signal type_cast_222_inst_ack_1 : boolean;
  signal addr_of_570_final_reg_req_1 : boolean;
  signal if_stmt_498_branch_ack_0 : boolean;
  signal if_stmt_498_branch_ack_1 : boolean;
  signal type_cast_644_inst_ack_1 : boolean;
  signal if_stmt_498_branch_req_0 : boolean;
  signal type_cast_680_inst_req_0 : boolean;
  signal array_obj_ref_569_index_offset_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_658_inst_ack_1 : boolean;
  signal addr_of_570_final_reg_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_640_inst_ack_1 : boolean;
  signal type_cast_698_inst_req_1 : boolean;
  signal type_cast_1199_inst_req_0 : boolean;
  signal type_cast_577_inst_req_0 : boolean;
  signal type_cast_698_inst_ack_1 : boolean;
  signal type_cast_1199_inst_ack_0 : boolean;
  signal ptr_deref_706_store_0_ack_1 : boolean;
  signal if_stmt_513_branch_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_573_inst_req_0 : boolean;
  signal ptr_deref_706_store_0_req_1 : boolean;
  signal if_stmt_513_branch_ack_1 : boolean;
  signal array_obj_ref_1120_index_offset_ack_0 : boolean;
  signal addr_of_570_final_reg_ack_1 : boolean;
  signal if_stmt_513_branch_req_0 : boolean;
  signal type_cast_1139_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_218_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_218_inst_ack_1 : boolean;
  signal type_cast_608_inst_ack_1 : boolean;
  signal type_cast_608_inst_req_1 : boolean;
  signal WPIPE_Concat_output_pipe_1204_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_640_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_658_inst_req_0 : boolean;
  signal array_obj_ref_1120_index_offset_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_658_inst_ack_0 : boolean;
  signal addr_of_570_final_reg_ack_0 : boolean;
  signal type_cast_577_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_676_inst_ack_0 : boolean;
  signal type_cast_458_inst_ack_1 : boolean;
  signal type_cast_644_inst_req_1 : boolean;
  signal type_cast_680_inst_ack_0 : boolean;
  signal type_cast_644_inst_req_0 : boolean;
  signal WPIPE_Concat_output_pipe_1201_inst_req_1 : boolean;
  signal type_cast_1139_inst_ack_0 : boolean;
  signal array_obj_ref_569_index_offset_req_1 : boolean;
  signal array_obj_ref_569_index_offset_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_694_inst_ack_0 : boolean;
  signal type_cast_1169_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_622_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_640_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_694_inst_req_0 : boolean;
  signal type_cast_1169_inst_req_1 : boolean;
  signal addr_of_1121_final_reg_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_573_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_622_inst_req_1 : boolean;
  signal type_cast_577_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_622_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_231_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_231_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_231_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_231_inst_ack_1 : boolean;
  signal type_cast_608_inst_req_0 : boolean;
  signal type_cast_235_inst_req_0 : boolean;
  signal type_cast_235_inst_ack_0 : boolean;
  signal type_cast_235_inst_req_1 : boolean;
  signal type_cast_235_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_243_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_243_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_243_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_243_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_694_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1204_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_604_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_604_inst_req_1 : boolean;
  signal type_cast_247_inst_req_0 : boolean;
  signal type_cast_247_inst_ack_0 : boolean;
  signal WPIPE_Concat_output_pipe_1201_inst_ack_1 : boolean;
  signal type_cast_247_inst_req_1 : boolean;
  signal type_cast_247_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_256_inst_req_0 : boolean;
  signal type_cast_626_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_256_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_256_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_256_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_694_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_604_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_604_inst_req_0 : boolean;
  signal type_cast_662_inst_ack_1 : boolean;
  signal type_cast_260_inst_req_0 : boolean;
  signal type_cast_626_inst_req_1 : boolean;
  signal type_cast_260_inst_ack_0 : boolean;
  signal array_obj_ref_1120_index_offset_req_1 : boolean;
  signal type_cast_260_inst_req_1 : boolean;
  signal WPIPE_Concat_output_pipe_1055_inst_req_0 : boolean;
  signal type_cast_260_inst_ack_1 : boolean;
  signal type_cast_1179_inst_ack_0 : boolean;
  signal WPIPE_Concat_output_pipe_1049_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_268_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_268_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_268_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_268_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1040_inst_ack_1 : boolean;
  signal type_cast_590_inst_ack_1 : boolean;
  signal type_cast_590_inst_req_1 : boolean;
  signal type_cast_662_inst_req_1 : boolean;
  signal type_cast_272_inst_req_0 : boolean;
  signal type_cast_272_inst_ack_0 : boolean;
  signal type_cast_272_inst_req_1 : boolean;
  signal type_cast_626_inst_ack_0 : boolean;
  signal type_cast_272_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_281_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_281_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_676_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_281_inst_req_1 : boolean;
  signal type_cast_626_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_281_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1055_inst_ack_0 : boolean;
  signal type_cast_590_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_676_inst_req_1 : boolean;
  signal type_cast_590_inst_req_0 : boolean;
  signal type_cast_285_inst_req_0 : boolean;
  signal type_cast_285_inst_ack_0 : boolean;
  signal type_cast_285_inst_req_1 : boolean;
  signal type_cast_285_inst_ack_1 : boolean;
  signal type_cast_527_inst_ack_1 : boolean;
  signal type_cast_527_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_586_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_293_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_293_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_293_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_293_inst_ack_1 : boolean;
  signal type_cast_662_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_586_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_586_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_586_inst_req_0 : boolean;
  signal type_cast_662_inst_ack_0 : boolean;
  signal type_cast_297_inst_req_0 : boolean;
  signal type_cast_297_inst_ack_0 : boolean;
  signal type_cast_297_inst_req_1 : boolean;
  signal type_cast_297_inst_ack_1 : boolean;
  signal type_cast_527_inst_ack_0 : boolean;
  signal WPIPE_Concat_output_pipe_1207_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_306_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_306_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_306_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_306_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1049_inst_ack_1 : boolean;
  signal addr_of_1121_final_reg_req_1 : boolean;
  signal addr_of_1121_final_reg_ack_1 : boolean;
  signal type_cast_310_inst_req_0 : boolean;
  signal type_cast_310_inst_ack_0 : boolean;
  signal type_cast_310_inst_req_1 : boolean;
  signal type_cast_1149_inst_req_0 : boolean;
  signal type_cast_310_inst_ack_1 : boolean;
  signal type_cast_1179_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_318_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_318_inst_ack_0 : boolean;
  signal WPIPE_Concat_output_pipe_1207_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_318_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_318_inst_ack_1 : boolean;
  signal type_cast_322_inst_req_0 : boolean;
  signal type_cast_322_inst_ack_0 : boolean;
  signal type_cast_322_inst_req_1 : boolean;
  signal type_cast_322_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_331_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_331_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_331_inst_req_1 : boolean;
  signal type_cast_1149_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_331_inst_ack_1 : boolean;
  signal type_cast_335_inst_req_0 : boolean;
  signal type_cast_335_inst_ack_0 : boolean;
  signal type_cast_335_inst_req_1 : boolean;
  signal type_cast_335_inst_ack_1 : boolean;
  signal type_cast_1179_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_343_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_343_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_343_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_343_inst_ack_1 : boolean;
  signal type_cast_347_inst_req_0 : boolean;
  signal type_cast_1149_inst_req_1 : boolean;
  signal type_cast_347_inst_ack_0 : boolean;
  signal type_cast_347_inst_req_1 : boolean;
  signal type_cast_1149_inst_ack_1 : boolean;
  signal type_cast_347_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1040_inst_req_0 : boolean;
  signal type_cast_1199_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_356_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_356_inst_ack_0 : boolean;
  signal WPIPE_Concat_output_pipe_1043_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_356_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_356_inst_ack_1 : boolean;
  signal type_cast_360_inst_req_0 : boolean;
  signal type_cast_360_inst_ack_0 : boolean;
  signal type_cast_360_inst_req_1 : boolean;
  signal type_cast_360_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1052_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_368_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_368_inst_ack_0 : boolean;
  signal WPIPE_Concat_output_pipe_1052_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_368_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_368_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1052_inst_req_1 : boolean;
  signal type_cast_372_inst_req_0 : boolean;
  signal type_cast_372_inst_ack_0 : boolean;
  signal type_cast_372_inst_req_1 : boolean;
  signal type_cast_372_inst_ack_1 : boolean;
  signal ptr_deref_1125_load_0_req_0 : boolean;
  signal type_cast_1199_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_381_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_381_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_381_inst_req_1 : boolean;
  signal WPIPE_Concat_output_pipe_1052_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_381_inst_ack_1 : boolean;
  signal type_cast_385_inst_req_0 : boolean;
  signal type_cast_385_inst_ack_0 : boolean;
  signal type_cast_385_inst_req_1 : boolean;
  signal type_cast_385_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_393_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_393_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_393_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_393_inst_ack_1 : boolean;
  signal type_cast_397_inst_req_0 : boolean;
  signal type_cast_397_inst_ack_0 : boolean;
  signal type_cast_397_inst_req_1 : boolean;
  signal type_cast_397_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_406_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_406_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_406_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_406_inst_ack_1 : boolean;
  signal type_cast_410_inst_req_0 : boolean;
  signal type_cast_410_inst_ack_0 : boolean;
  signal type_cast_410_inst_req_1 : boolean;
  signal type_cast_410_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_418_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_418_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_418_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_418_inst_ack_1 : boolean;
  signal type_cast_422_inst_req_0 : boolean;
  signal type_cast_422_inst_ack_0 : boolean;
  signal type_cast_422_inst_req_1 : boolean;
  signal type_cast_422_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_431_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_431_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_431_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_431_inst_ack_1 : boolean;
  signal type_cast_435_inst_req_0 : boolean;
  signal type_cast_435_inst_ack_0 : boolean;
  signal type_cast_435_inst_req_1 : boolean;
  signal type_cast_435_inst_ack_1 : boolean;
  signal type_cast_444_inst_req_0 : boolean;
  signal type_cast_444_inst_ack_0 : boolean;
  signal type_cast_444_inst_req_1 : boolean;
  signal type_cast_444_inst_ack_1 : boolean;
  signal if_stmt_720_branch_req_0 : boolean;
  signal if_stmt_720_branch_ack_1 : boolean;
  signal if_stmt_720_branch_ack_0 : boolean;
  signal WPIPE_Concat_output_pipe_1040_inst_req_1 : boolean;
  signal type_cast_734_inst_req_0 : boolean;
  signal type_cast_734_inst_ack_0 : boolean;
  signal WPIPE_Concat_output_pipe_1037_inst_ack_1 : boolean;
  signal type_cast_734_inst_req_1 : boolean;
  signal type_cast_734_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1204_inst_ack_0 : boolean;
  signal WPIPE_Concat_output_pipe_1207_inst_req_1 : boolean;
  signal WPIPE_Concat_output_pipe_1037_inst_req_1 : boolean;
  signal array_obj_ref_776_index_offset_req_0 : boolean;
  signal array_obj_ref_776_index_offset_ack_0 : boolean;
  signal array_obj_ref_776_index_offset_req_1 : boolean;
  signal type_cast_1129_inst_ack_1 : boolean;
  signal array_obj_ref_776_index_offset_ack_1 : boolean;
  signal type_cast_1129_inst_req_1 : boolean;
  signal WPIPE_Concat_output_pipe_1204_inst_req_0 : boolean;
  signal WPIPE_Concat_output_pipe_1201_inst_ack_0 : boolean;
  signal addr_of_777_final_reg_req_0 : boolean;
  signal addr_of_777_final_reg_ack_0 : boolean;
  signal addr_of_777_final_reg_req_1 : boolean;
  signal type_cast_1129_inst_ack_0 : boolean;
  signal addr_of_777_final_reg_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1046_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1046_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_780_inst_req_0 : boolean;
  signal type_cast_1129_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_780_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_780_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_780_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1207_inst_ack_1 : boolean;
  signal if_stmt_1068_branch_ack_0 : boolean;
  signal WPIPE_Concat_output_pipe_1201_inst_req_0 : boolean;
  signal type_cast_784_inst_req_0 : boolean;
  signal type_cast_784_inst_ack_0 : boolean;
  signal type_cast_784_inst_req_1 : boolean;
  signal type_cast_784_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1046_inst_ack_0 : boolean;
  signal type_cast_1159_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_793_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_793_inst_ack_0 : boolean;
  signal WPIPE_Concat_output_pipe_1046_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_793_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_793_inst_ack_1 : boolean;
  signal if_stmt_1068_branch_ack_1 : boolean;
  signal if_stmt_1068_branch_req_0 : boolean;
  signal type_cast_797_inst_req_0 : boolean;
  signal type_cast_797_inst_ack_0 : boolean;
  signal type_cast_797_inst_req_1 : boolean;
  signal type_cast_797_inst_ack_1 : boolean;
  signal type_cast_1159_inst_req_1 : boolean;
  signal type_cast_1189_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_811_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_811_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_811_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_811_inst_ack_1 : boolean;
  signal type_cast_815_inst_req_0 : boolean;
  signal type_cast_815_inst_ack_0 : boolean;
  signal type_cast_815_inst_req_1 : boolean;
  signal ptr_deref_1125_load_0_ack_1 : boolean;
  signal type_cast_815_inst_ack_1 : boolean;
  signal type_cast_1159_inst_ack_0 : boolean;
  signal type_cast_1189_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_829_inst_req_0 : boolean;
  signal ptr_deref_1125_load_0_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_829_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_829_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_829_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1058_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1058_inst_req_1 : boolean;
  signal WPIPE_Concat_output_pipe_1058_inst_ack_0 : boolean;
  signal WPIPE_Concat_output_pipe_1058_inst_req_0 : boolean;
  signal type_cast_833_inst_req_0 : boolean;
  signal type_cast_833_inst_ack_0 : boolean;
  signal type_cast_833_inst_req_1 : boolean;
  signal type_cast_833_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1043_inst_ack_1 : boolean;
  signal type_cast_1159_inst_req_0 : boolean;
  signal WPIPE_Concat_output_pipe_1043_inst_req_1 : boolean;
  signal type_cast_1189_inst_ack_0 : boolean;
  signal type_cast_1189_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_847_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_847_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_847_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_847_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1055_inst_ack_1 : boolean;
  signal type_cast_851_inst_req_0 : boolean;
  signal type_cast_851_inst_ack_0 : boolean;
  signal type_cast_851_inst_req_1 : boolean;
  signal type_cast_851_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_865_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_865_inst_ack_0 : boolean;
  signal WPIPE_Concat_output_pipe_1043_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_865_inst_req_1 : boolean;
  signal ptr_deref_1125_load_0_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_865_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1055_inst_req_1 : boolean;
  signal WPIPE_Concat_output_pipe_1040_inst_ack_0 : boolean;
  signal type_cast_869_inst_req_0 : boolean;
  signal type_cast_869_inst_ack_0 : boolean;
  signal type_cast_869_inst_req_1 : boolean;
  signal type_cast_869_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_883_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_883_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_883_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_883_inst_ack_1 : boolean;
  signal type_cast_887_inst_req_0 : boolean;
  signal type_cast_887_inst_ack_0 : boolean;
  signal type_cast_887_inst_req_1 : boolean;
  signal type_cast_887_inst_ack_1 : boolean;
  signal RPIPE_Concat_input_pipe_901_inst_req_0 : boolean;
  signal RPIPE_Concat_input_pipe_901_inst_ack_0 : boolean;
  signal RPIPE_Concat_input_pipe_901_inst_req_1 : boolean;
  signal RPIPE_Concat_input_pipe_901_inst_ack_1 : boolean;
  signal type_cast_905_inst_req_0 : boolean;
  signal type_cast_905_inst_ack_0 : boolean;
  signal type_cast_905_inst_req_1 : boolean;
  signal type_cast_905_inst_ack_1 : boolean;
  signal ptr_deref_913_store_0_req_0 : boolean;
  signal ptr_deref_913_store_0_ack_0 : boolean;
  signal ptr_deref_913_store_0_req_1 : boolean;
  signal ptr_deref_913_store_0_ack_1 : boolean;
  signal if_stmt_927_branch_req_0 : boolean;
  signal if_stmt_927_branch_ack_1 : boolean;
  signal if_stmt_927_branch_ack_0 : boolean;
  signal call_stmt_938_call_req_0 : boolean;
  signal call_stmt_938_call_ack_0 : boolean;
  signal call_stmt_938_call_req_1 : boolean;
  signal call_stmt_938_call_ack_1 : boolean;
  signal type_cast_943_inst_req_0 : boolean;
  signal type_cast_943_inst_ack_0 : boolean;
  signal type_cast_943_inst_req_1 : boolean;
  signal type_cast_943_inst_ack_1 : boolean;
  signal call_stmt_949_call_req_0 : boolean;
  signal call_stmt_949_call_ack_0 : boolean;
  signal call_stmt_949_call_req_1 : boolean;
  signal call_stmt_949_call_ack_1 : boolean;
  signal call_stmt_952_call_req_0 : boolean;
  signal call_stmt_952_call_ack_0 : boolean;
  signal call_stmt_952_call_req_1 : boolean;
  signal call_stmt_952_call_ack_1 : boolean;
  signal type_cast_956_inst_req_0 : boolean;
  signal type_cast_956_inst_ack_0 : boolean;
  signal type_cast_956_inst_req_1 : boolean;
  signal type_cast_956_inst_ack_1 : boolean;
  signal type_cast_965_inst_req_0 : boolean;
  signal type_cast_965_inst_ack_0 : boolean;
  signal type_cast_965_inst_req_1 : boolean;
  signal type_cast_965_inst_ack_1 : boolean;
  signal type_cast_975_inst_req_0 : boolean;
  signal type_cast_975_inst_ack_0 : boolean;
  signal type_cast_975_inst_req_1 : boolean;
  signal type_cast_975_inst_ack_1 : boolean;
  signal type_cast_985_inst_req_0 : boolean;
  signal type_cast_985_inst_ack_0 : boolean;
  signal type_cast_985_inst_req_1 : boolean;
  signal type_cast_985_inst_ack_1 : boolean;
  signal type_cast_995_inst_req_0 : boolean;
  signal type_cast_995_inst_ack_0 : boolean;
  signal type_cast_995_inst_req_1 : boolean;
  signal type_cast_995_inst_ack_1 : boolean;
  signal type_cast_1005_inst_req_0 : boolean;
  signal type_cast_1005_inst_ack_0 : boolean;
  signal type_cast_1005_inst_req_1 : boolean;
  signal type_cast_1005_inst_ack_1 : boolean;
  signal type_cast_1015_inst_req_0 : boolean;
  signal type_cast_1015_inst_ack_0 : boolean;
  signal type_cast_1015_inst_req_1 : boolean;
  signal type_cast_1015_inst_ack_1 : boolean;
  signal type_cast_1025_inst_req_0 : boolean;
  signal type_cast_1025_inst_ack_0 : boolean;
  signal type_cast_1025_inst_req_1 : boolean;
  signal type_cast_1025_inst_ack_1 : boolean;
  signal type_cast_1035_inst_req_0 : boolean;
  signal type_cast_1035_inst_ack_0 : boolean;
  signal type_cast_1035_inst_req_1 : boolean;
  signal type_cast_1035_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1037_inst_req_0 : boolean;
  signal WPIPE_Concat_output_pipe_1037_inst_ack_0 : boolean;
  signal WPIPE_Concat_output_pipe_1210_inst_req_0 : boolean;
  signal WPIPE_Concat_output_pipe_1210_inst_ack_0 : boolean;
  signal WPIPE_Concat_output_pipe_1210_inst_req_1 : boolean;
  signal WPIPE_Concat_output_pipe_1210_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1213_inst_req_0 : boolean;
  signal WPIPE_Concat_output_pipe_1213_inst_ack_0 : boolean;
  signal WPIPE_Concat_output_pipe_1213_inst_req_1 : boolean;
  signal WPIPE_Concat_output_pipe_1213_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1216_inst_req_0 : boolean;
  signal WPIPE_Concat_output_pipe_1216_inst_ack_0 : boolean;
  signal WPIPE_Concat_output_pipe_1216_inst_req_1 : boolean;
  signal WPIPE_Concat_output_pipe_1216_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1219_inst_req_0 : boolean;
  signal WPIPE_Concat_output_pipe_1219_inst_ack_0 : boolean;
  signal WPIPE_Concat_output_pipe_1219_inst_req_1 : boolean;
  signal WPIPE_Concat_output_pipe_1219_inst_ack_1 : boolean;
  signal WPIPE_Concat_output_pipe_1222_inst_req_0 : boolean;
  signal WPIPE_Concat_output_pipe_1222_inst_ack_0 : boolean;
  signal WPIPE_Concat_output_pipe_1222_inst_req_1 : boolean;
  signal WPIPE_Concat_output_pipe_1222_inst_ack_1 : boolean;
  signal if_stmt_1236_branch_req_0 : boolean;
  signal if_stmt_1236_branch_ack_1 : boolean;
  signal if_stmt_1236_branch_ack_0 : boolean;
  signal phi_stmt_555_req_0 : boolean;
  signal type_cast_561_inst_req_0 : boolean;
  signal type_cast_561_inst_ack_0 : boolean;
  signal type_cast_561_inst_req_1 : boolean;
  signal type_cast_561_inst_ack_1 : boolean;
  signal phi_stmt_555_req_1 : boolean;
  signal phi_stmt_555_ack_0 : boolean;
  signal phi_stmt_762_req_0 : boolean;
  signal type_cast_768_inst_req_0 : boolean;
  signal type_cast_768_inst_ack_0 : boolean;
  signal type_cast_768_inst_req_1 : boolean;
  signal type_cast_768_inst_ack_1 : boolean;
  signal phi_stmt_762_req_1 : boolean;
  signal phi_stmt_762_ack_0 : boolean;
  signal phi_stmt_1106_req_0 : boolean;
  signal type_cast_1112_inst_req_0 : boolean;
  signal type_cast_1112_inst_ack_0 : boolean;
  signal type_cast_1112_inst_req_1 : boolean;
  signal type_cast_1112_inst_ack_1 : boolean;
  signal phi_stmt_1106_req_1 : boolean;
  signal phi_stmt_1106_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "concat_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  concat_CP_664_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "concat_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= concat_CP_664_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= concat_CP_664_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= concat_CP_664_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  concat_CP_664: Block -- control-path 
    signal concat_CP_664_elements: BooleanArray(291 downto 0);
    -- 
  begin -- 
    concat_CP_664_elements(0) <= concat_CP_664_start;
    concat_CP_664_symbol <= concat_CP_664_elements(291);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	56 
    -- CP-element group 0: 	72 
    -- CP-element group 0: 	75 
    -- CP-element group 0: 	78 
    -- CP-element group 0: 	36 
    -- CP-element group 0: 	44 
    -- CP-element group 0: 	52 
    -- CP-element group 0: 	48 
    -- CP-element group 0: 	40 
    -- CP-element group 0: 	60 
    -- CP-element group 0: 	64 
    -- CP-element group 0: 	68 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	8 
    -- CP-element group 0: 	12 
    -- CP-element group 0: 	16 
    -- CP-element group 0: 	20 
    -- CP-element group 0: 	24 
    -- CP-element group 0: 	28 
    -- CP-element group 0: 	32 
    -- CP-element group 0:  members (68) 
      -- CP-element group 0: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_458_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_216/branch_block_stmt_216__entry__
      -- CP-element group 0: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_458_update_start_
      -- CP-element group 0: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_218_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_458_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_222_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_222_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/$entry
      -- CP-element group 0: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497__entry__
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_218_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_222_update_start_
      -- CP-element group 0: 	 branch_block_stmt_216/$entry
      -- CP-element group 0: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_218_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_235_update_start_
      -- CP-element group 0: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_235_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_235_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_247_update_start_
      -- CP-element group 0: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_247_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_247_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_260_update_start_
      -- CP-element group 0: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_260_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_260_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_272_update_start_
      -- CP-element group 0: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_272_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_272_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_285_update_start_
      -- CP-element group 0: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_285_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_285_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_297_update_start_
      -- CP-element group 0: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_297_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_297_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_310_update_start_
      -- CP-element group 0: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_310_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_310_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_322_update_start_
      -- CP-element group 0: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_322_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_322_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_335_update_start_
      -- CP-element group 0: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_335_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_335_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_347_update_start_
      -- CP-element group 0: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_347_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_347_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_360_update_start_
      -- CP-element group 0: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_360_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_360_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_372_update_start_
      -- CP-element group 0: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_372_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_372_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_385_update_start_
      -- CP-element group 0: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_385_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_385_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_397_update_start_
      -- CP-element group 0: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_397_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_397_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_410_update_start_
      -- CP-element group 0: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_410_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_410_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_422_update_start_
      -- CP-element group 0: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_422_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_422_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_435_update_start_
      -- CP-element group 0: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_435_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_435_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_444_update_start_
      -- CP-element group 0: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_444_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_444_Update/cr
      -- 
    rr_744_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_744_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(0), ack => RPIPE_Concat_input_pipe_218_inst_req_0); -- 
    cr_1267_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1267_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(0), ack => type_cast_458_inst_req_1); -- 
    cr_763_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_763_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(0), ack => type_cast_222_inst_req_1); -- 
    cr_791_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_791_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(0), ack => type_cast_235_inst_req_1); -- 
    cr_819_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_819_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(0), ack => type_cast_247_inst_req_1); -- 
    cr_847_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_847_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(0), ack => type_cast_260_inst_req_1); -- 
    cr_875_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_875_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(0), ack => type_cast_272_inst_req_1); -- 
    cr_903_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_903_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(0), ack => type_cast_285_inst_req_1); -- 
    cr_931_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_931_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(0), ack => type_cast_297_inst_req_1); -- 
    cr_959_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_959_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(0), ack => type_cast_310_inst_req_1); -- 
    cr_987_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_987_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(0), ack => type_cast_322_inst_req_1); -- 
    cr_1015_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1015_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(0), ack => type_cast_335_inst_req_1); -- 
    cr_1043_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1043_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(0), ack => type_cast_347_inst_req_1); -- 
    cr_1071_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1071_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(0), ack => type_cast_360_inst_req_1); -- 
    cr_1099_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1099_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(0), ack => type_cast_372_inst_req_1); -- 
    cr_1127_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1127_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(0), ack => type_cast_385_inst_req_1); -- 
    cr_1155_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1155_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(0), ack => type_cast_397_inst_req_1); -- 
    cr_1183_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1183_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(0), ack => type_cast_410_inst_req_1); -- 
    cr_1211_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1211_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(0), ack => type_cast_422_inst_req_1); -- 
    cr_1239_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1239_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(0), ack => type_cast_435_inst_req_1); -- 
    cr_1253_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1253_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(0), ack => type_cast_444_inst_req_1); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_218_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_218_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_218_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_218_Update/cr
      -- CP-element group 1: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_218_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_218_update_start_
      -- 
    ra_745_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_218_inst_ack_0, ack => concat_CP_664_elements(1)); -- 
    cr_749_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_749_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(1), ack => RPIPE_Concat_input_pipe_218_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (9) 
      -- CP-element group 2: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_222_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_222_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_218_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_218_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_218_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_222_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_231_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_231_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_231_Sample/rr
      -- 
    ca_750_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_218_inst_ack_1, ack => concat_CP_664_elements(2)); -- 
    rr_758_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_758_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(2), ack => type_cast_222_inst_req_0); -- 
    rr_772_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_772_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(2), ack => RPIPE_Concat_input_pipe_231_inst_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_222_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_222_Sample/ra
      -- CP-element group 3: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_222_sample_completed_
      -- 
    ra_759_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_222_inst_ack_0, ack => concat_CP_664_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	79 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_222_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_222_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_222_Update/ca
      -- 
    ca_764_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_222_inst_ack_1, ack => concat_CP_664_elements(4)); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_231_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_231_update_start_
      -- CP-element group 5: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_231_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_231_Sample/ra
      -- CP-element group 5: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_231_Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_231_Update/cr
      -- 
    ra_773_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_231_inst_ack_0, ack => concat_CP_664_elements(5)); -- 
    cr_777_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_777_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(5), ack => RPIPE_Concat_input_pipe_231_inst_req_1); -- 
    -- CP-element group 6:  fork  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6: 	9 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_231_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_231_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_231_Update/ca
      -- CP-element group 6: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_235_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_235_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_235_Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_243_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_243_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_243_Sample/rr
      -- 
    ca_778_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_231_inst_ack_1, ack => concat_CP_664_elements(6)); -- 
    rr_786_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_786_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(6), ack => type_cast_235_inst_req_0); -- 
    rr_800_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_800_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(6), ack => RPIPE_Concat_input_pipe_243_inst_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_235_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_235_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_235_Sample/ra
      -- 
    ra_787_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_235_inst_ack_0, ack => concat_CP_664_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	0 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	79 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_235_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_235_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_235_Update/ca
      -- 
    ca_792_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_235_inst_ack_1, ack => concat_CP_664_elements(8)); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	6 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_243_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_243_update_start_
      -- CP-element group 9: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_243_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_243_Sample/ra
      -- CP-element group 9: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_243_Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_243_Update/cr
      -- 
    ra_801_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_243_inst_ack_0, ack => concat_CP_664_elements(9)); -- 
    cr_805_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_805_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(9), ack => RPIPE_Concat_input_pipe_243_inst_req_1); -- 
    -- CP-element group 10:  fork  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10: 	13 
    -- CP-element group 10:  members (9) 
      -- CP-element group 10: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_243_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_243_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_243_Update/ca
      -- CP-element group 10: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_247_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_247_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_247_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_256_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_256_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_256_Sample/rr
      -- 
    ca_806_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_243_inst_ack_1, ack => concat_CP_664_elements(10)); -- 
    rr_814_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_814_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(10), ack => type_cast_247_inst_req_0); -- 
    rr_828_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_828_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(10), ack => RPIPE_Concat_input_pipe_256_inst_req_0); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_247_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_247_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_247_Sample/ra
      -- 
    ra_815_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_247_inst_ack_0, ack => concat_CP_664_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	0 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	79 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_247_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_247_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_247_Update/ca
      -- 
    ca_820_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_247_inst_ack_1, ack => concat_CP_664_elements(12)); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	10 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_256_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_256_update_start_
      -- CP-element group 13: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_256_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_256_Sample/ra
      -- CP-element group 13: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_256_Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_256_Update/cr
      -- 
    ra_829_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_256_inst_ack_0, ack => concat_CP_664_elements(13)); -- 
    cr_833_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_833_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(13), ack => RPIPE_Concat_input_pipe_256_inst_req_1); -- 
    -- CP-element group 14:  fork  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14: 	17 
    -- CP-element group 14:  members (9) 
      -- CP-element group 14: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_256_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_256_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_256_Update/ca
      -- CP-element group 14: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_260_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_260_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_260_Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_268_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_268_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_268_Sample/rr
      -- 
    ca_834_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_256_inst_ack_1, ack => concat_CP_664_elements(14)); -- 
    rr_842_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_842_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(14), ack => type_cast_260_inst_req_0); -- 
    rr_856_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_856_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(14), ack => RPIPE_Concat_input_pipe_268_inst_req_0); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_260_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_260_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_260_Sample/ra
      -- 
    ra_843_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_260_inst_ack_0, ack => concat_CP_664_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	0 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	79 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_260_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_260_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_260_Update/ca
      -- 
    ca_848_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_260_inst_ack_1, ack => concat_CP_664_elements(16)); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	14 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_268_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_268_update_start_
      -- CP-element group 17: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_268_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_268_Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_268_Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_268_Update/cr
      -- 
    ra_857_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_268_inst_ack_0, ack => concat_CP_664_elements(17)); -- 
    cr_861_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_861_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(17), ack => RPIPE_Concat_input_pipe_268_inst_req_1); -- 
    -- CP-element group 18:  fork  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18: 	21 
    -- CP-element group 18:  members (9) 
      -- CP-element group 18: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_268_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_268_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_268_Update/ca
      -- CP-element group 18: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_272_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_272_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_272_Sample/rr
      -- CP-element group 18: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_281_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_281_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_281_Sample/rr
      -- 
    ca_862_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_268_inst_ack_1, ack => concat_CP_664_elements(18)); -- 
    rr_870_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_870_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(18), ack => type_cast_272_inst_req_0); -- 
    rr_884_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_884_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(18), ack => RPIPE_Concat_input_pipe_281_inst_req_0); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_272_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_272_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_272_Sample/ra
      -- 
    ra_871_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_272_inst_ack_0, ack => concat_CP_664_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	0 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	73 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_272_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_272_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_272_Update/ca
      -- 
    ca_876_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_272_inst_ack_1, ack => concat_CP_664_elements(20)); -- 
    -- CP-element group 21:  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	18 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (6) 
      -- CP-element group 21: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_281_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_281_update_start_
      -- CP-element group 21: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_281_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_281_Sample/ra
      -- CP-element group 21: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_281_Update/$entry
      -- CP-element group 21: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_281_Update/cr
      -- 
    ra_885_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_281_inst_ack_0, ack => concat_CP_664_elements(21)); -- 
    cr_889_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_889_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(21), ack => RPIPE_Concat_input_pipe_281_inst_req_1); -- 
    -- CP-element group 22:  fork  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22: 	25 
    -- CP-element group 22:  members (9) 
      -- CP-element group 22: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_281_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_281_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_281_Update/ca
      -- CP-element group 22: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_285_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_285_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_285_Sample/rr
      -- CP-element group 22: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_293_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_293_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_293_Sample/rr
      -- 
    ca_890_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_281_inst_ack_1, ack => concat_CP_664_elements(22)); -- 
    rr_898_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_898_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(22), ack => type_cast_285_inst_req_0); -- 
    rr_912_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_912_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(22), ack => RPIPE_Concat_input_pipe_293_inst_req_0); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_285_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_285_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_285_Sample/ra
      -- 
    ra_899_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_285_inst_ack_0, ack => concat_CP_664_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	0 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	73 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_285_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_285_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_285_Update/ca
      -- 
    ca_904_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_285_inst_ack_1, ack => concat_CP_664_elements(24)); -- 
    -- CP-element group 25:  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	22 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25:  members (6) 
      -- CP-element group 25: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_293_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_293_update_start_
      -- CP-element group 25: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_293_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_293_Sample/ra
      -- CP-element group 25: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_293_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_293_Update/cr
      -- 
    ra_913_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_293_inst_ack_0, ack => concat_CP_664_elements(25)); -- 
    cr_917_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_917_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(25), ack => RPIPE_Concat_input_pipe_293_inst_req_1); -- 
    -- CP-element group 26:  fork  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: 	29 
    -- CP-element group 26:  members (9) 
      -- CP-element group 26: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_293_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_293_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_293_Update/ca
      -- CP-element group 26: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_297_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_297_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_297_Sample/rr
      -- CP-element group 26: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_306_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_306_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_306_Sample/rr
      -- 
    ca_918_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_293_inst_ack_1, ack => concat_CP_664_elements(26)); -- 
    rr_926_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_926_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(26), ack => type_cast_297_inst_req_0); -- 
    rr_940_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_940_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(26), ack => RPIPE_Concat_input_pipe_306_inst_req_0); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_297_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_297_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_297_Sample/ra
      -- 
    ra_927_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_297_inst_ack_0, ack => concat_CP_664_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	0 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	79 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_297_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_297_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_297_Update/ca
      -- 
    ca_932_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_297_inst_ack_1, ack => concat_CP_664_elements(28)); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	26 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_306_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_306_update_start_
      -- CP-element group 29: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_306_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_306_Sample/ra
      -- CP-element group 29: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_306_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_306_Update/cr
      -- 
    ra_941_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_306_inst_ack_0, ack => concat_CP_664_elements(29)); -- 
    cr_945_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_945_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(29), ack => RPIPE_Concat_input_pipe_306_inst_req_1); -- 
    -- CP-element group 30:  fork  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30: 	33 
    -- CP-element group 30:  members (9) 
      -- CP-element group 30: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_306_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_306_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_306_Update/ca
      -- CP-element group 30: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_310_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_310_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_310_Sample/rr
      -- CP-element group 30: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_318_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_318_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_318_Sample/rr
      -- 
    ca_946_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_306_inst_ack_1, ack => concat_CP_664_elements(30)); -- 
    rr_954_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_954_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(30), ack => type_cast_310_inst_req_0); -- 
    rr_968_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_968_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(30), ack => RPIPE_Concat_input_pipe_318_inst_req_0); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_310_sample_completed_
      -- CP-element group 31: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_310_Sample/$exit
      -- CP-element group 31: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_310_Sample/ra
      -- 
    ra_955_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_310_inst_ack_0, ack => concat_CP_664_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	0 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	79 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_310_update_completed_
      -- CP-element group 32: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_310_Update/$exit
      -- CP-element group 32: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_310_Update/ca
      -- 
    ca_960_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_310_inst_ack_1, ack => concat_CP_664_elements(32)); -- 
    -- CP-element group 33:  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	30 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (6) 
      -- CP-element group 33: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_318_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_318_update_start_
      -- CP-element group 33: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_318_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_318_Sample/ra
      -- CP-element group 33: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_318_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_318_Update/cr
      -- 
    ra_969_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_318_inst_ack_0, ack => concat_CP_664_elements(33)); -- 
    cr_973_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_973_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(33), ack => RPIPE_Concat_input_pipe_318_inst_req_1); -- 
    -- CP-element group 34:  fork  transition  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	37 
    -- CP-element group 34: 	35 
    -- CP-element group 34:  members (9) 
      -- CP-element group 34: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_318_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_318_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_318_Update/ca
      -- CP-element group 34: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_322_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_322_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_322_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_331_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_331_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_331_Sample/rr
      -- 
    ca_974_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_318_inst_ack_1, ack => concat_CP_664_elements(34)); -- 
    rr_982_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_982_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(34), ack => type_cast_322_inst_req_0); -- 
    rr_996_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_996_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(34), ack => RPIPE_Concat_input_pipe_331_inst_req_0); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_322_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_322_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_322_Sample/ra
      -- 
    ra_983_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_322_inst_ack_0, ack => concat_CP_664_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	0 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	79 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_322_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_322_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_322_Update/ca
      -- 
    ca_988_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_322_inst_ack_1, ack => concat_CP_664_elements(36)); -- 
    -- CP-element group 37:  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (6) 
      -- CP-element group 37: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_331_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_331_update_start_
      -- CP-element group 37: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_331_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_331_Sample/ra
      -- CP-element group 37: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_331_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_331_Update/cr
      -- 
    ra_997_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_331_inst_ack_0, ack => concat_CP_664_elements(37)); -- 
    cr_1001_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1001_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(37), ack => RPIPE_Concat_input_pipe_331_inst_req_1); -- 
    -- CP-element group 38:  fork  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38: 	41 
    -- CP-element group 38:  members (9) 
      -- CP-element group 38: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_331_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_331_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_331_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_335_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_335_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_335_Sample/rr
      -- CP-element group 38: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_343_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_343_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_343_Sample/rr
      -- 
    ca_1002_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_331_inst_ack_1, ack => concat_CP_664_elements(38)); -- 
    rr_1024_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1024_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(38), ack => RPIPE_Concat_input_pipe_343_inst_req_0); -- 
    rr_1010_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1010_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(38), ack => type_cast_335_inst_req_0); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_335_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_335_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_335_Sample/ra
      -- 
    ra_1011_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_335_inst_ack_0, ack => concat_CP_664_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	0 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	79 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_335_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_335_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_335_Update/ca
      -- 
    ca_1016_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_335_inst_ack_1, ack => concat_CP_664_elements(40)); -- 
    -- CP-element group 41:  transition  input  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	38 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (6) 
      -- CP-element group 41: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_343_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_343_update_start_
      -- CP-element group 41: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_343_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_343_Sample/ra
      -- CP-element group 41: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_343_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_343_Update/cr
      -- 
    ra_1025_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_343_inst_ack_0, ack => concat_CP_664_elements(41)); -- 
    cr_1029_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1029_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(41), ack => RPIPE_Concat_input_pipe_343_inst_req_1); -- 
    -- CP-element group 42:  fork  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	45 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (9) 
      -- CP-element group 42: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_343_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_343_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_343_Update/ca
      -- CP-element group 42: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_347_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_347_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_347_Sample/rr
      -- CP-element group 42: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_356_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_356_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_356_Sample/rr
      -- 
    ca_1030_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_343_inst_ack_1, ack => concat_CP_664_elements(42)); -- 
    rr_1038_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1038_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(42), ack => type_cast_347_inst_req_0); -- 
    rr_1052_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1052_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(42), ack => RPIPE_Concat_input_pipe_356_inst_req_0); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_347_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_347_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_347_Sample/ra
      -- 
    ra_1039_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_347_inst_ack_0, ack => concat_CP_664_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	0 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	76 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_347_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_347_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_347_Update/ca
      -- 
    ca_1044_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_347_inst_ack_1, ack => concat_CP_664_elements(44)); -- 
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	42 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (6) 
      -- CP-element group 45: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_356_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_356_update_start_
      -- CP-element group 45: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_356_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_356_Sample/ra
      -- CP-element group 45: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_356_Update/$entry
      -- CP-element group 45: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_356_Update/cr
      -- 
    ra_1053_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_356_inst_ack_0, ack => concat_CP_664_elements(45)); -- 
    cr_1057_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1057_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(45), ack => RPIPE_Concat_input_pipe_356_inst_req_1); -- 
    -- CP-element group 46:  fork  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46: 	49 
    -- CP-element group 46:  members (9) 
      -- CP-element group 46: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_356_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_356_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_356_Update/ca
      -- CP-element group 46: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_360_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_360_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_360_Sample/rr
      -- CP-element group 46: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_368_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_368_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_368_Sample/rr
      -- 
    ca_1058_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_356_inst_ack_1, ack => concat_CP_664_elements(46)); -- 
    rr_1080_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1080_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(46), ack => RPIPE_Concat_input_pipe_368_inst_req_0); -- 
    rr_1066_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1066_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(46), ack => type_cast_360_inst_req_0); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_360_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_360_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_360_Sample/ra
      -- 
    ra_1067_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_360_inst_ack_0, ack => concat_CP_664_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	0 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	76 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_360_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_360_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_360_Update/ca
      -- 
    ca_1072_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_360_inst_ack_1, ack => concat_CP_664_elements(48)); -- 
    -- CP-element group 49:  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	46 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (6) 
      -- CP-element group 49: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_368_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_368_update_start_
      -- CP-element group 49: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_368_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_368_Sample/ra
      -- CP-element group 49: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_368_Update/$entry
      -- CP-element group 49: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_368_Update/cr
      -- 
    ra_1081_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_368_inst_ack_0, ack => concat_CP_664_elements(49)); -- 
    cr_1085_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1085_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(49), ack => RPIPE_Concat_input_pipe_368_inst_req_1); -- 
    -- CP-element group 50:  fork  transition  input  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	53 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (9) 
      -- CP-element group 50: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_368_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_368_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_368_Update/ca
      -- CP-element group 50: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_372_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_372_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_372_Sample/rr
      -- CP-element group 50: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_381_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_381_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_381_Sample/rr
      -- 
    ca_1086_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_368_inst_ack_1, ack => concat_CP_664_elements(50)); -- 
    rr_1094_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1094_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(50), ack => type_cast_372_inst_req_0); -- 
    rr_1108_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1108_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(50), ack => RPIPE_Concat_input_pipe_381_inst_req_0); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_372_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_372_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_372_Sample/ra
      -- 
    ra_1095_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_372_inst_ack_0, ack => concat_CP_664_elements(51)); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	0 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	79 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_372_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_372_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_372_Update/ca
      -- 
    ca_1100_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_372_inst_ack_1, ack => concat_CP_664_elements(52)); -- 
    -- CP-element group 53:  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	50 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (6) 
      -- CP-element group 53: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_381_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_381_update_start_
      -- CP-element group 53: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_381_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_381_Sample/ra
      -- CP-element group 53: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_381_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_381_Update/cr
      -- 
    ra_1109_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_381_inst_ack_0, ack => concat_CP_664_elements(53)); -- 
    cr_1113_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1113_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(53), ack => RPIPE_Concat_input_pipe_381_inst_req_1); -- 
    -- CP-element group 54:  fork  transition  input  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	57 
    -- CP-element group 54: 	55 
    -- CP-element group 54:  members (9) 
      -- CP-element group 54: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_381_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_381_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_381_Update/ca
      -- CP-element group 54: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_385_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_385_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_385_Sample/rr
      -- CP-element group 54: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_393_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_393_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_393_Sample/rr
      -- 
    ca_1114_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_381_inst_ack_1, ack => concat_CP_664_elements(54)); -- 
    rr_1136_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1136_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(54), ack => RPIPE_Concat_input_pipe_393_inst_req_0); -- 
    rr_1122_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1122_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(54), ack => type_cast_385_inst_req_0); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_385_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_385_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_385_Sample/ra
      -- 
    ra_1123_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_385_inst_ack_0, ack => concat_CP_664_elements(55)); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	0 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	79 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_385_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_385_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_385_Update/ca
      -- 
    ca_1128_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_385_inst_ack_1, ack => concat_CP_664_elements(56)); -- 
    -- CP-element group 57:  transition  input  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	54 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (6) 
      -- CP-element group 57: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_393_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_393_update_start_
      -- CP-element group 57: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_393_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_393_Sample/ra
      -- CP-element group 57: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_393_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_393_Update/cr
      -- 
    ra_1137_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_393_inst_ack_0, ack => concat_CP_664_elements(57)); -- 
    cr_1141_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1141_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(57), ack => RPIPE_Concat_input_pipe_393_inst_req_1); -- 
    -- CP-element group 58:  fork  transition  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58: 	61 
    -- CP-element group 58:  members (9) 
      -- CP-element group 58: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_393_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_393_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_393_Update/ca
      -- CP-element group 58: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_397_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_397_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_397_Sample/rr
      -- CP-element group 58: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_406_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_406_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_406_Sample/rr
      -- 
    ca_1142_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_393_inst_ack_1, ack => concat_CP_664_elements(58)); -- 
    rr_1150_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1150_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(58), ack => type_cast_397_inst_req_0); -- 
    rr_1164_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1164_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(58), ack => RPIPE_Concat_input_pipe_406_inst_req_0); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_397_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_397_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_397_Sample/ra
      -- 
    ra_1151_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_397_inst_ack_0, ack => concat_CP_664_elements(59)); -- 
    -- CP-element group 60:  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	0 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	79 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_397_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_397_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_397_Update/ca
      -- 
    ca_1156_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_397_inst_ack_1, ack => concat_CP_664_elements(60)); -- 
    -- CP-element group 61:  transition  input  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	58 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61:  members (6) 
      -- CP-element group 61: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_406_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_406_update_start_
      -- CP-element group 61: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_406_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_406_Sample/ra
      -- CP-element group 61: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_406_Update/$entry
      -- CP-element group 61: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_406_Update/cr
      -- 
    ra_1165_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_406_inst_ack_0, ack => concat_CP_664_elements(61)); -- 
    cr_1169_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1169_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(61), ack => RPIPE_Concat_input_pipe_406_inst_req_1); -- 
    -- CP-element group 62:  fork  transition  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62: 	65 
    -- CP-element group 62:  members (9) 
      -- CP-element group 62: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_406_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_406_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_406_Update/ca
      -- CP-element group 62: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_410_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_410_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_410_Sample/rr
      -- CP-element group 62: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_418_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_418_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_418_Sample/rr
      -- 
    ca_1170_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_406_inst_ack_1, ack => concat_CP_664_elements(62)); -- 
    rr_1178_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1178_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(62), ack => type_cast_410_inst_req_0); -- 
    rr_1192_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1192_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(62), ack => RPIPE_Concat_input_pipe_418_inst_req_0); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_410_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_410_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_410_Sample/ra
      -- 
    ra_1179_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_410_inst_ack_0, ack => concat_CP_664_elements(63)); -- 
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	0 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	79 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_410_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_410_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_410_Update/ca
      -- 
    ca_1184_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_410_inst_ack_1, ack => concat_CP_664_elements(64)); -- 
    -- CP-element group 65:  transition  input  output  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	62 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65:  members (6) 
      -- CP-element group 65: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_418_sample_completed_
      -- CP-element group 65: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_418_update_start_
      -- CP-element group 65: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_418_Sample/$exit
      -- CP-element group 65: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_418_Sample/ra
      -- CP-element group 65: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_418_Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_418_Update/cr
      -- 
    ra_1193_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_418_inst_ack_0, ack => concat_CP_664_elements(65)); -- 
    cr_1197_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1197_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(65), ack => RPIPE_Concat_input_pipe_418_inst_req_1); -- 
    -- CP-element group 66:  fork  transition  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	65 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	69 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (9) 
      -- CP-element group 66: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_418_update_completed_
      -- CP-element group 66: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_418_Update/$exit
      -- CP-element group 66: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_418_Update/ca
      -- CP-element group 66: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_422_sample_start_
      -- CP-element group 66: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_422_Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_422_Sample/rr
      -- CP-element group 66: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_431_sample_start_
      -- CP-element group 66: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_431_Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_431_Sample/rr
      -- 
    ca_1198_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_418_inst_ack_1, ack => concat_CP_664_elements(66)); -- 
    rr_1220_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1220_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(66), ack => RPIPE_Concat_input_pipe_431_inst_req_0); -- 
    rr_1206_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1206_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(66), ack => type_cast_422_inst_req_0); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_422_sample_completed_
      -- CP-element group 67: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_422_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_422_Sample/ra
      -- 
    ra_1207_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_422_inst_ack_0, ack => concat_CP_664_elements(67)); -- 
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	0 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	79 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_422_update_completed_
      -- CP-element group 68: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_422_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_422_Update/ca
      -- 
    ca_1212_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_422_inst_ack_1, ack => concat_CP_664_elements(68)); -- 
    -- CP-element group 69:  transition  input  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	66 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69:  members (6) 
      -- CP-element group 69: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_431_sample_completed_
      -- CP-element group 69: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_431_update_start_
      -- CP-element group 69: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_431_Sample/$exit
      -- CP-element group 69: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_431_Sample/ra
      -- CP-element group 69: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_431_Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_431_Update/cr
      -- 
    ra_1221_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_431_inst_ack_0, ack => concat_CP_664_elements(69)); -- 
    cr_1225_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1225_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(69), ack => RPIPE_Concat_input_pipe_431_inst_req_1); -- 
    -- CP-element group 70:  transition  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70:  members (6) 
      -- CP-element group 70: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_431_update_completed_
      -- CP-element group 70: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_431_Update/$exit
      -- CP-element group 70: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/RPIPE_Concat_input_pipe_431_Update/ca
      -- CP-element group 70: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_435_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_435_Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_435_Sample/rr
      -- 
    ca_1226_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_431_inst_ack_1, ack => concat_CP_664_elements(70)); -- 
    rr_1234_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1234_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(70), ack => type_cast_435_inst_req_0); -- 
    -- CP-element group 71:  transition  input  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_435_sample_completed_
      -- CP-element group 71: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_435_Sample/$exit
      -- CP-element group 71: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_435_Sample/ra
      -- 
    ra_1235_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_435_inst_ack_0, ack => concat_CP_664_elements(71)); -- 
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	0 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	79 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_435_update_completed_
      -- CP-element group 72: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_435_Update/$exit
      -- CP-element group 72: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_435_Update/ca
      -- 
    ca_1240_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_435_inst_ack_1, ack => concat_CP_664_elements(72)); -- 
    -- CP-element group 73:  join  transition  output  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	20 
    -- CP-element group 73: 	24 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_444_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_444_Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_444_Sample/rr
      -- 
    rr_1248_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1248_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(73), ack => type_cast_444_inst_req_0); -- 
    concat_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 26) := "concat_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_664_elements(20) & concat_CP_664_elements(24);
      gj_concat_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_664_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_444_sample_completed_
      -- CP-element group 74: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_444_Sample/$exit
      -- CP-element group 74: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_444_Sample/ra
      -- 
    ra_1249_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_444_inst_ack_0, ack => concat_CP_664_elements(74)); -- 
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	0 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	79 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_444_update_completed_
      -- CP-element group 75: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_444_Update/$exit
      -- CP-element group 75: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_444_Update/ca
      -- 
    ca_1254_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_444_inst_ack_1, ack => concat_CP_664_elements(75)); -- 
    -- CP-element group 76:  join  transition  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	44 
    -- CP-element group 76: 	48 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_458_Sample/rr
      -- CP-element group 76: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_458_Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_458_sample_start_
      -- 
    rr_1262_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1262_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(76), ack => type_cast_458_inst_req_0); -- 
    concat_cp_element_group_76: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 26) := "concat_cp_element_group_76"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_664_elements(44) & concat_CP_664_elements(48);
      gj_concat_cp_element_group_76 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_664_elements(76), clk => clk, reset => reset); --
    end block;
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	76 
    -- CP-element group 77: successors 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_458_Sample/ra
      -- CP-element group 77: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_458_Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_458_sample_completed_
      -- 
    ra_1263_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_458_inst_ack_0, ack => concat_CP_664_elements(77)); -- 
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	0 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_458_update_completed_
      -- CP-element group 78: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_458_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/type_cast_458_Update/ca
      -- 
    ca_1268_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_458_inst_ack_1, ack => concat_CP_664_elements(78)); -- 
    -- CP-element group 79:  branch  join  transition  place  output  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	56 
    -- CP-element group 79: 	72 
    -- CP-element group 79: 	75 
    -- CP-element group 79: 	78 
    -- CP-element group 79: 	36 
    -- CP-element group 79: 	52 
    -- CP-element group 79: 	40 
    -- CP-element group 79: 	60 
    -- CP-element group 79: 	64 
    -- CP-element group 79: 	68 
    -- CP-element group 79: 	4 
    -- CP-element group 79: 	8 
    -- CP-element group 79: 	12 
    -- CP-element group 79: 	16 
    -- CP-element group 79: 	28 
    -- CP-element group 79: 	32 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79: 	81 
    -- CP-element group 79:  members (10) 
      -- CP-element group 79: 	 branch_block_stmt_216/if_stmt_498_eval_test/$entry
      -- CP-element group 79: 	 branch_block_stmt_216/if_stmt_498_else_link/$entry
      -- CP-element group 79: 	 branch_block_stmt_216/R_cmp388_499_place
      -- CP-element group 79: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497/$exit
      -- CP-element group 79: 	 branch_block_stmt_216/if_stmt_498_eval_test/branch_req
      -- CP-element group 79: 	 branch_block_stmt_216/if_stmt_498_eval_test/$exit
      -- CP-element group 79: 	 branch_block_stmt_216/if_stmt_498__entry__
      -- CP-element group 79: 	 branch_block_stmt_216/assign_stmt_219_to_assign_stmt_497__exit__
      -- CP-element group 79: 	 branch_block_stmt_216/if_stmt_498_dead_link/$entry
      -- CP-element group 79: 	 branch_block_stmt_216/if_stmt_498_if_link/$entry
      -- 
    branch_req_1276_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1276_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(79), ack => if_stmt_498_branch_req_0); -- 
    concat_cp_element_group_79: block -- 
      constant place_capacities: IntegerArray(0 to 15) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1);
      constant place_markings: IntegerArray(0 to 15)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0);
      constant place_delays: IntegerArray(0 to 15) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0);
      constant joinName: string(1 to 26) := "concat_cp_element_group_79"; 
      signal preds: BooleanArray(1 to 16); -- 
    begin -- 
      preds <= concat_CP_664_elements(56) & concat_CP_664_elements(72) & concat_CP_664_elements(75) & concat_CP_664_elements(78) & concat_CP_664_elements(36) & concat_CP_664_elements(52) & concat_CP_664_elements(40) & concat_CP_664_elements(60) & concat_CP_664_elements(64) & concat_CP_664_elements(68) & concat_CP_664_elements(4) & concat_CP_664_elements(8) & concat_CP_664_elements(12) & concat_CP_664_elements(16) & concat_CP_664_elements(28) & concat_CP_664_elements(32);
      gj_concat_cp_element_group_79 : generic_join generic map(name => joinName, number_of_predecessors => 16, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_664_elements(79), clk => clk, reset => reset); --
    end block;
    -- CP-element group 80:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	84 
    -- CP-element group 80: 	85 
    -- CP-element group 80:  members (18) 
      -- CP-element group 80: 	 branch_block_stmt_216/assign_stmt_524_to_assign_stmt_552/$entry
      -- CP-element group 80: 	 branch_block_stmt_216/assign_stmt_524_to_assign_stmt_552/type_cast_527_Sample/rr
      -- CP-element group 80: 	 branch_block_stmt_216/if_stmt_498_if_link/if_choice_transition
      -- CP-element group 80: 	 branch_block_stmt_216/assign_stmt_524_to_assign_stmt_552/type_cast_527_update_start_
      -- CP-element group 80: 	 branch_block_stmt_216/if_stmt_498_if_link/$exit
      -- CP-element group 80: 	 branch_block_stmt_216/assign_stmt_524_to_assign_stmt_552__entry__
      -- CP-element group 80: 	 branch_block_stmt_216/entry_bbx_xnph390
      -- CP-element group 80: 	 branch_block_stmt_216/assign_stmt_524_to_assign_stmt_552/type_cast_527_Sample/$entry
      -- CP-element group 80: 	 branch_block_stmt_216/assign_stmt_524_to_assign_stmt_552/type_cast_527_sample_start_
      -- CP-element group 80: 	 branch_block_stmt_216/merge_stmt_519__exit__
      -- CP-element group 80: 	 branch_block_stmt_216/assign_stmt_524_to_assign_stmt_552/type_cast_527_Update/cr
      -- CP-element group 80: 	 branch_block_stmt_216/assign_stmt_524_to_assign_stmt_552/type_cast_527_Update/$entry
      -- CP-element group 80: 	 branch_block_stmt_216/entry_bbx_xnph390_PhiReq/$entry
      -- CP-element group 80: 	 branch_block_stmt_216/entry_bbx_xnph390_PhiReq/$exit
      -- CP-element group 80: 	 branch_block_stmt_216/merge_stmt_519_PhiReqMerge
      -- CP-element group 80: 	 branch_block_stmt_216/merge_stmt_519_PhiAck/$entry
      -- CP-element group 80: 	 branch_block_stmt_216/merge_stmt_519_PhiAck/$exit
      -- CP-element group 80: 	 branch_block_stmt_216/merge_stmt_519_PhiAck/dummy
      -- 
    if_choice_transition_1281_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_498_branch_ack_1, ack => concat_CP_664_elements(80)); -- 
    rr_1320_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1320_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(80), ack => type_cast_527_inst_req_0); -- 
    cr_1325_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1325_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(80), ack => type_cast_527_inst_req_1); -- 
    -- CP-element group 81:  transition  place  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	79 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	271 
    -- CP-element group 81:  members (5) 
      -- CP-element group 81: 	 branch_block_stmt_216/if_stmt_498_else_link/else_choice_transition
      -- CP-element group 81: 	 branch_block_stmt_216/if_stmt_498_else_link/$exit
      -- CP-element group 81: 	 branch_block_stmt_216/entry_forx_xcond165x_xpreheader
      -- CP-element group 81: 	 branch_block_stmt_216/entry_forx_xcond165x_xpreheader_PhiReq/$entry
      -- CP-element group 81: 	 branch_block_stmt_216/entry_forx_xcond165x_xpreheader_PhiReq/$exit
      -- 
    else_choice_transition_1285_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_498_branch_ack_0, ack => concat_CP_664_elements(81)); -- 
    -- CP-element group 82:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	271 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	128 
    -- CP-element group 82: 	129 
    -- CP-element group 82:  members (18) 
      -- CP-element group 82: 	 branch_block_stmt_216/merge_stmt_726__exit__
      -- CP-element group 82: 	 branch_block_stmt_216/if_stmt_513_if_link/if_choice_transition
      -- CP-element group 82: 	 branch_block_stmt_216/forx_xcond165x_xpreheader_bbx_xnph386
      -- CP-element group 82: 	 branch_block_stmt_216/assign_stmt_731_to_assign_stmt_759__entry__
      -- CP-element group 82: 	 branch_block_stmt_216/if_stmt_513_if_link/$exit
      -- CP-element group 82: 	 branch_block_stmt_216/assign_stmt_731_to_assign_stmt_759/$entry
      -- CP-element group 82: 	 branch_block_stmt_216/assign_stmt_731_to_assign_stmt_759/type_cast_734_sample_start_
      -- CP-element group 82: 	 branch_block_stmt_216/assign_stmt_731_to_assign_stmt_759/type_cast_734_update_start_
      -- CP-element group 82: 	 branch_block_stmt_216/assign_stmt_731_to_assign_stmt_759/type_cast_734_Sample/$entry
      -- CP-element group 82: 	 branch_block_stmt_216/assign_stmt_731_to_assign_stmt_759/type_cast_734_Sample/rr
      -- CP-element group 82: 	 branch_block_stmt_216/assign_stmt_731_to_assign_stmt_759/type_cast_734_Update/$entry
      -- CP-element group 82: 	 branch_block_stmt_216/assign_stmt_731_to_assign_stmt_759/type_cast_734_Update/cr
      -- CP-element group 82: 	 branch_block_stmt_216/forx_xcond165x_xpreheader_bbx_xnph386_PhiReq/$entry
      -- CP-element group 82: 	 branch_block_stmt_216/forx_xcond165x_xpreheader_bbx_xnph386_PhiReq/$exit
      -- CP-element group 82: 	 branch_block_stmt_216/merge_stmt_726_PhiReqMerge
      -- CP-element group 82: 	 branch_block_stmt_216/merge_stmt_726_PhiAck/$entry
      -- CP-element group 82: 	 branch_block_stmt_216/merge_stmt_726_PhiAck/$exit
      -- CP-element group 82: 	 branch_block_stmt_216/merge_stmt_726_PhiAck/dummy
      -- 
    if_choice_transition_1303_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_513_branch_ack_1, ack => concat_CP_664_elements(82)); -- 
    rr_1679_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1679_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(82), ack => type_cast_734_inst_req_0); -- 
    cr_1684_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1684_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(82), ack => type_cast_734_inst_req_1); -- 
    -- CP-element group 83:  transition  place  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	271 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	284 
    -- CP-element group 83:  members (5) 
      -- CP-element group 83: 	 branch_block_stmt_216/if_stmt_513_else_link/$exit
      -- CP-element group 83: 	 branch_block_stmt_216/forx_xcond165x_xpreheader_forx_xend224
      -- CP-element group 83: 	 branch_block_stmt_216/if_stmt_513_else_link/else_choice_transition
      -- CP-element group 83: 	 branch_block_stmt_216/forx_xcond165x_xpreheader_forx_xend224_PhiReq/$entry
      -- CP-element group 83: 	 branch_block_stmt_216/forx_xcond165x_xpreheader_forx_xend224_PhiReq/$exit
      -- 
    else_choice_transition_1307_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_513_branch_ack_0, ack => concat_CP_664_elements(83)); -- 
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	80 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_216/assign_stmt_524_to_assign_stmt_552/type_cast_527_sample_completed_
      -- CP-element group 84: 	 branch_block_stmt_216/assign_stmt_524_to_assign_stmt_552/type_cast_527_Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_216/assign_stmt_524_to_assign_stmt_552/type_cast_527_Sample/ra
      -- 
    ra_1321_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_527_inst_ack_0, ack => concat_CP_664_elements(84)); -- 
    -- CP-element group 85:  transition  place  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	80 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	272 
    -- CP-element group 85:  members (9) 
      -- CP-element group 85: 	 branch_block_stmt_216/assign_stmt_524_to_assign_stmt_552/type_cast_527_update_completed_
      -- CP-element group 85: 	 branch_block_stmt_216/assign_stmt_524_to_assign_stmt_552/$exit
      -- CP-element group 85: 	 branch_block_stmt_216/bbx_xnph390_forx_xbody
      -- CP-element group 85: 	 branch_block_stmt_216/assign_stmt_524_to_assign_stmt_552__exit__
      -- CP-element group 85: 	 branch_block_stmt_216/assign_stmt_524_to_assign_stmt_552/type_cast_527_Update/ca
      -- CP-element group 85: 	 branch_block_stmt_216/assign_stmt_524_to_assign_stmt_552/type_cast_527_Update/$exit
      -- CP-element group 85: 	 branch_block_stmt_216/bbx_xnph390_forx_xbody_PhiReq/$entry
      -- CP-element group 85: 	 branch_block_stmt_216/bbx_xnph390_forx_xbody_PhiReq/phi_stmt_555/$entry
      -- CP-element group 85: 	 branch_block_stmt_216/bbx_xnph390_forx_xbody_PhiReq/phi_stmt_555/phi_stmt_555_sources/$entry
      -- 
    ca_1326_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_527_inst_ack_1, ack => concat_CP_664_elements(85)); -- 
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	277 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	125 
    -- CP-element group 86:  members (3) 
      -- CP-element group 86: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/array_obj_ref_569_final_index_sum_regn_Sample/ack
      -- CP-element group 86: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/array_obj_ref_569_final_index_sum_regn_Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/array_obj_ref_569_final_index_sum_regn_sample_complete
      -- 
    ack_1355_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_569_index_offset_ack_0, ack => concat_CP_664_elements(86)); -- 
    -- CP-element group 87:  transition  input  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	277 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (11) 
      -- CP-element group 87: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/array_obj_ref_569_base_plus_offset/sum_rename_req
      -- CP-element group 87: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/array_obj_ref_569_base_plus_offset/$entry
      -- CP-element group 87: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/array_obj_ref_569_base_plus_offset/sum_rename_ack
      -- CP-element group 87: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/addr_of_570_request/$entry
      -- CP-element group 87: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/array_obj_ref_569_final_index_sum_regn_Update/ack
      -- CP-element group 87: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/addr_of_570_request/req
      -- CP-element group 87: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/array_obj_ref_569_final_index_sum_regn_Update/$exit
      -- CP-element group 87: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/array_obj_ref_569_base_plus_offset/$exit
      -- CP-element group 87: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/array_obj_ref_569_offset_calculated
      -- CP-element group 87: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/array_obj_ref_569_root_address_calculated
      -- CP-element group 87: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/addr_of_570_sample_start_
      -- 
    ack_1360_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_569_index_offset_ack_1, ack => concat_CP_664_elements(87)); -- 
    req_1369_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1369_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(87), ack => addr_of_570_final_reg_req_0); -- 
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/addr_of_570_request/$exit
      -- CP-element group 88: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/addr_of_570_request/ack
      -- CP-element group 88: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/addr_of_570_sample_completed_
      -- 
    ack_1370_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_570_final_reg_ack_0, ack => concat_CP_664_elements(88)); -- 
    -- CP-element group 89:  fork  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	277 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	122 
    -- CP-element group 89:  members (19) 
      -- CP-element group 89: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/ptr_deref_706_base_address_resized
      -- CP-element group 89: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/ptr_deref_706_base_plus_offset/$entry
      -- CP-element group 89: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/ptr_deref_706_base_addr_resize/$entry
      -- CP-element group 89: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/ptr_deref_706_root_address_calculated
      -- CP-element group 89: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/addr_of_570_complete/$exit
      -- CP-element group 89: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/ptr_deref_706_base_addr_resize/$exit
      -- CP-element group 89: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/ptr_deref_706_base_address_calculated
      -- CP-element group 89: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/ptr_deref_706_base_plus_offset/sum_rename_ack
      -- CP-element group 89: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/ptr_deref_706_base_addr_resize/base_resize_req
      -- CP-element group 89: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/ptr_deref_706_base_plus_offset/$exit
      -- CP-element group 89: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/ptr_deref_706_word_address_calculated
      -- CP-element group 89: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/addr_of_570_complete/ack
      -- CP-element group 89: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/ptr_deref_706_base_plus_offset/sum_rename_req
      -- CP-element group 89: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/ptr_deref_706_word_addrgen/root_register_ack
      -- CP-element group 89: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/ptr_deref_706_base_addr_resize/base_resize_ack
      -- CP-element group 89: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/addr_of_570_update_completed_
      -- CP-element group 89: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/ptr_deref_706_word_addrgen/root_register_req
      -- CP-element group 89: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/ptr_deref_706_word_addrgen/$entry
      -- CP-element group 89: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/ptr_deref_706_word_addrgen/$exit
      -- 
    ack_1375_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_570_final_reg_ack_1, ack => concat_CP_664_elements(89)); -- 
    -- CP-element group 90:  transition  input  output  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	277 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (6) 
      -- CP-element group 90: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_573_Sample/ra
      -- CP-element group 90: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_573_Update/cr
      -- CP-element group 90: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_573_Update/$entry
      -- CP-element group 90: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_573_Sample/$exit
      -- CP-element group 90: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_573_sample_completed_
      -- CP-element group 90: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_573_update_start_
      -- 
    ra_1384_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_573_inst_ack_0, ack => concat_CP_664_elements(90)); -- 
    cr_1388_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1388_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(90), ack => RPIPE_Concat_input_pipe_573_inst_req_1); -- 
    -- CP-element group 91:  fork  transition  input  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91: 	94 
    -- CP-element group 91:  members (9) 
      -- CP-element group 91: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_577_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_573_update_completed_
      -- CP-element group 91: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_573_Update/$exit
      -- CP-element group 91: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_577_Sample/rr
      -- CP-element group 91: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_577_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_573_Update/ca
      -- CP-element group 91: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_586_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_586_Sample/rr
      -- CP-element group 91: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_586_Sample/$entry
      -- 
    ca_1389_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_573_inst_ack_1, ack => concat_CP_664_elements(91)); -- 
    rr_1397_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1397_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(91), ack => type_cast_577_inst_req_0); -- 
    rr_1411_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1411_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(91), ack => RPIPE_Concat_input_pipe_586_inst_req_0); -- 
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92:  members (3) 
      -- CP-element group 92: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_577_Sample/$exit
      -- CP-element group 92: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_577_Sample/ra
      -- CP-element group 92: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_577_sample_completed_
      -- 
    ra_1398_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_577_inst_ack_0, ack => concat_CP_664_elements(92)); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	277 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	122 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_577_update_completed_
      -- CP-element group 93: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_577_Update/$exit
      -- CP-element group 93: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_577_Update/ca
      -- 
    ca_1403_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_577_inst_ack_1, ack => concat_CP_664_elements(93)); -- 
    -- CP-element group 94:  transition  input  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	91 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94:  members (6) 
      -- CP-element group 94: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_586_sample_completed_
      -- CP-element group 94: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_586_Update/cr
      -- CP-element group 94: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_586_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_586_Sample/ra
      -- CP-element group 94: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_586_Sample/$exit
      -- CP-element group 94: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_586_update_start_
      -- 
    ra_1412_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_586_inst_ack_0, ack => concat_CP_664_elements(94)); -- 
    cr_1416_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1416_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(94), ack => RPIPE_Concat_input_pipe_586_inst_req_1); -- 
    -- CP-element group 95:  fork  transition  input  output  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95: 	98 
    -- CP-element group 95:  members (9) 
      -- CP-element group 95: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_604_Sample/rr
      -- CP-element group 95: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_604_Sample/$entry
      -- CP-element group 95: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_604_sample_start_
      -- CP-element group 95: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_590_Sample/rr
      -- CP-element group 95: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_590_Sample/$entry
      -- CP-element group 95: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_590_sample_start_
      -- CP-element group 95: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_586_Update/ca
      -- CP-element group 95: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_586_Update/$exit
      -- CP-element group 95: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_586_update_completed_
      -- 
    ca_1417_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_586_inst_ack_1, ack => concat_CP_664_elements(95)); -- 
    rr_1425_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1425_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(95), ack => type_cast_590_inst_req_0); -- 
    rr_1439_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1439_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(95), ack => RPIPE_Concat_input_pipe_604_inst_req_0); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_590_Sample/ra
      -- CP-element group 96: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_590_Sample/$exit
      -- CP-element group 96: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_590_sample_completed_
      -- 
    ra_1426_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_590_inst_ack_0, ack => concat_CP_664_elements(96)); -- 
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	277 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	122 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_590_Update/ca
      -- CP-element group 97: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_590_Update/$exit
      -- CP-element group 97: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_590_update_completed_
      -- 
    ca_1431_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_590_inst_ack_1, ack => concat_CP_664_elements(97)); -- 
    -- CP-element group 98:  transition  input  output  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	95 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (6) 
      -- CP-element group 98: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_604_Update/cr
      -- CP-element group 98: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_604_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_604_Sample/ra
      -- CP-element group 98: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_604_Sample/$exit
      -- CP-element group 98: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_604_update_start_
      -- CP-element group 98: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_604_sample_completed_
      -- 
    ra_1440_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_604_inst_ack_0, ack => concat_CP_664_elements(98)); -- 
    cr_1444_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1444_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(98), ack => RPIPE_Concat_input_pipe_604_inst_req_1); -- 
    -- CP-element group 99:  fork  transition  input  output  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	98 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99: 	102 
    -- CP-element group 99:  members (9) 
      -- CP-element group 99: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_622_Sample/$entry
      -- CP-element group 99: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_622_sample_start_
      -- CP-element group 99: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_622_Sample/rr
      -- CP-element group 99: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_608_Sample/rr
      -- CP-element group 99: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_608_Sample/$entry
      -- CP-element group 99: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_608_sample_start_
      -- CP-element group 99: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_604_Update/ca
      -- CP-element group 99: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_604_Update/$exit
      -- CP-element group 99: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_604_update_completed_
      -- 
    ca_1445_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_604_inst_ack_1, ack => concat_CP_664_elements(99)); -- 
    rr_1453_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1453_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(99), ack => type_cast_608_inst_req_0); -- 
    rr_1467_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1467_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(99), ack => RPIPE_Concat_input_pipe_622_inst_req_0); -- 
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100:  members (3) 
      -- CP-element group 100: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_608_Sample/ra
      -- CP-element group 100: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_608_Sample/$exit
      -- CP-element group 100: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_608_sample_completed_
      -- 
    ra_1454_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_608_inst_ack_0, ack => concat_CP_664_elements(100)); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	277 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	122 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_608_Update/$exit
      -- CP-element group 101: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_608_Update/ca
      -- CP-element group 101: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_608_update_completed_
      -- 
    ca_1459_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_608_inst_ack_1, ack => concat_CP_664_elements(101)); -- 
    -- CP-element group 102:  transition  input  output  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	99 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	103 
    -- CP-element group 102:  members (6) 
      -- CP-element group 102: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_622_update_start_
      -- CP-element group 102: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_622_Sample/ra
      -- CP-element group 102: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_622_sample_completed_
      -- CP-element group 102: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_622_Sample/$exit
      -- CP-element group 102: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_622_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_622_Update/cr
      -- 
    ra_1468_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_622_inst_ack_0, ack => concat_CP_664_elements(102)); -- 
    cr_1472_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1472_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(102), ack => RPIPE_Concat_input_pipe_622_inst_req_1); -- 
    -- CP-element group 103:  fork  transition  input  output  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	102 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103: 	106 
    -- CP-element group 103:  members (9) 
      -- CP-element group 103: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_640_Sample/rr
      -- CP-element group 103: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_640_Sample/$entry
      -- CP-element group 103: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_626_sample_start_
      -- CP-element group 103: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_640_sample_start_
      -- CP-element group 103: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_622_update_completed_
      -- CP-element group 103: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_622_Update/$exit
      -- CP-element group 103: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_622_Update/ca
      -- CP-element group 103: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_626_Sample/rr
      -- CP-element group 103: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_626_Sample/$entry
      -- 
    ca_1473_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_622_inst_ack_1, ack => concat_CP_664_elements(103)); -- 
    rr_1481_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1481_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(103), ack => type_cast_626_inst_req_0); -- 
    rr_1495_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1495_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(103), ack => RPIPE_Concat_input_pipe_640_inst_req_0); -- 
    -- CP-element group 104:  transition  input  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (3) 
      -- CP-element group 104: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_626_sample_completed_
      -- CP-element group 104: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_626_Sample/ra
      -- CP-element group 104: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_626_Sample/$exit
      -- 
    ra_1482_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_626_inst_ack_0, ack => concat_CP_664_elements(104)); -- 
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	277 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	122 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_626_Update/ca
      -- CP-element group 105: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_626_Update/$exit
      -- CP-element group 105: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_626_update_completed_
      -- 
    ca_1487_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_626_inst_ack_1, ack => concat_CP_664_elements(105)); -- 
    -- CP-element group 106:  transition  input  output  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	103 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106:  members (6) 
      -- CP-element group 106: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_640_Update/$entry
      -- CP-element group 106: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_640_sample_completed_
      -- CP-element group 106: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_640_update_start_
      -- CP-element group 106: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_640_Sample/ra
      -- CP-element group 106: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_640_Sample/$exit
      -- CP-element group 106: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_640_Update/cr
      -- 
    ra_1496_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_640_inst_ack_0, ack => concat_CP_664_elements(106)); -- 
    cr_1500_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1500_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(106), ack => RPIPE_Concat_input_pipe_640_inst_req_1); -- 
    -- CP-element group 107:  fork  transition  input  output  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	106 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107: 	110 
    -- CP-element group 107:  members (9) 
      -- CP-element group 107: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_644_Sample/$entry
      -- CP-element group 107: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_640_Update/$exit
      -- CP-element group 107: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_640_update_completed_
      -- CP-element group 107: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_640_Update/ca
      -- CP-element group 107: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_658_Sample/rr
      -- CP-element group 107: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_644_Sample/rr
      -- CP-element group 107: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_658_Sample/$entry
      -- CP-element group 107: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_644_sample_start_
      -- CP-element group 107: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_658_sample_start_
      -- 
    ca_1501_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_640_inst_ack_1, ack => concat_CP_664_elements(107)); -- 
    rr_1509_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1509_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(107), ack => type_cast_644_inst_req_0); -- 
    rr_1523_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1523_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(107), ack => RPIPE_Concat_input_pipe_658_inst_req_0); -- 
    -- CP-element group 108:  transition  input  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108:  members (3) 
      -- CP-element group 108: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_644_Sample/ra
      -- CP-element group 108: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_644_Sample/$exit
      -- CP-element group 108: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_644_sample_completed_
      -- 
    ra_1510_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_644_inst_ack_0, ack => concat_CP_664_elements(108)); -- 
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	277 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	122 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_644_Update/$exit
      -- CP-element group 109: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_644_update_completed_
      -- CP-element group 109: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_644_Update/ca
      -- 
    ca_1515_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_644_inst_ack_1, ack => concat_CP_664_elements(109)); -- 
    -- CP-element group 110:  transition  input  output  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	107 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (6) 
      -- CP-element group 110: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_658_Update/$entry
      -- CP-element group 110: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_658_Update/cr
      -- CP-element group 110: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_658_Sample/ra
      -- CP-element group 110: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_658_Sample/$exit
      -- CP-element group 110: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_658_update_start_
      -- CP-element group 110: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_658_sample_completed_
      -- 
    ra_1524_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_658_inst_ack_0, ack => concat_CP_664_elements(110)); -- 
    cr_1528_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1528_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(110), ack => RPIPE_Concat_input_pipe_658_inst_req_1); -- 
    -- CP-element group 111:  fork  transition  input  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111: 	114 
    -- CP-element group 111:  members (9) 
      -- CP-element group 111: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_676_Sample/rr
      -- CP-element group 111: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_662_sample_start_
      -- CP-element group 111: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_658_Update/$exit
      -- CP-element group 111: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_658_Update/ca
      -- CP-element group 111: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_676_sample_start_
      -- CP-element group 111: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_662_Sample/$entry
      -- CP-element group 111: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_676_Sample/$entry
      -- CP-element group 111: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_658_update_completed_
      -- CP-element group 111: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_662_Sample/rr
      -- 
    ca_1529_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_658_inst_ack_1, ack => concat_CP_664_elements(111)); -- 
    rr_1537_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1537_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(111), ack => type_cast_662_inst_req_0); -- 
    rr_1551_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1551_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(111), ack => RPIPE_Concat_input_pipe_676_inst_req_0); -- 
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112:  members (3) 
      -- CP-element group 112: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_662_sample_completed_
      -- CP-element group 112: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_662_Sample/$exit
      -- CP-element group 112: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_662_Sample/ra
      -- 
    ra_1538_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_662_inst_ack_0, ack => concat_CP_664_elements(112)); -- 
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	277 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	122 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_662_update_completed_
      -- CP-element group 113: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_662_Update/ca
      -- CP-element group 113: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_662_Update/$exit
      -- 
    ca_1543_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_662_inst_ack_1, ack => concat_CP_664_elements(113)); -- 
    -- CP-element group 114:  transition  input  output  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	111 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (6) 
      -- CP-element group 114: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_676_Sample/$exit
      -- CP-element group 114: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_676_update_start_
      -- CP-element group 114: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_676_sample_completed_
      -- CP-element group 114: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_676_Sample/ra
      -- CP-element group 114: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_676_Update/cr
      -- CP-element group 114: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_676_Update/$entry
      -- 
    ra_1552_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_676_inst_ack_0, ack => concat_CP_664_elements(114)); -- 
    cr_1556_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1556_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(114), ack => RPIPE_Concat_input_pipe_676_inst_req_1); -- 
    -- CP-element group 115:  fork  transition  input  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	116 
    -- CP-element group 115: 	118 
    -- CP-element group 115:  members (9) 
      -- CP-element group 115: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_694_sample_start_
      -- CP-element group 115: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_680_sample_start_
      -- CP-element group 115: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_694_Sample/$entry
      -- CP-element group 115: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_680_Sample/rr
      -- CP-element group 115: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_676_update_completed_
      -- CP-element group 115: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_680_Sample/$entry
      -- CP-element group 115: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_694_Sample/rr
      -- CP-element group 115: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_676_Update/ca
      -- CP-element group 115: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_676_Update/$exit
      -- 
    ca_1557_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_676_inst_ack_1, ack => concat_CP_664_elements(115)); -- 
    rr_1565_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1565_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(115), ack => type_cast_680_inst_req_0); -- 
    rr_1579_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1579_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(115), ack => RPIPE_Concat_input_pipe_694_inst_req_0); -- 
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	115 
    -- CP-element group 116: successors 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_680_Sample/$exit
      -- CP-element group 116: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_680_sample_completed_
      -- CP-element group 116: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_680_Sample/ra
      -- 
    ra_1566_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_680_inst_ack_0, ack => concat_CP_664_elements(116)); -- 
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	277 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	122 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_680_Update/$exit
      -- CP-element group 117: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_680_Update/ca
      -- CP-element group 117: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_680_update_completed_
      -- 
    ca_1571_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_680_inst_ack_1, ack => concat_CP_664_elements(117)); -- 
    -- CP-element group 118:  transition  input  output  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	115 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	119 
    -- CP-element group 118:  members (6) 
      -- CP-element group 118: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_694_Update/$entry
      -- CP-element group 118: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_694_sample_completed_
      -- CP-element group 118: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_694_Sample/$exit
      -- CP-element group 118: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_694_update_start_
      -- CP-element group 118: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_694_Sample/ra
      -- CP-element group 118: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_694_Update/cr
      -- 
    ra_1580_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_694_inst_ack_0, ack => concat_CP_664_elements(118)); -- 
    cr_1584_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1584_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(118), ack => RPIPE_Concat_input_pipe_694_inst_req_1); -- 
    -- CP-element group 119:  transition  input  output  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	118 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	120 
    -- CP-element group 119:  members (6) 
      -- CP-element group 119: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_698_Sample/rr
      -- CP-element group 119: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_694_update_completed_
      -- CP-element group 119: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_694_Update/$exit
      -- CP-element group 119: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_698_Sample/$entry
      -- CP-element group 119: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_694_Update/ca
      -- CP-element group 119: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_698_sample_start_
      -- 
    ca_1585_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_694_inst_ack_1, ack => concat_CP_664_elements(119)); -- 
    rr_1593_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1593_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(119), ack => type_cast_698_inst_req_0); -- 
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	119 
    -- CP-element group 120: successors 
    -- CP-element group 120:  members (3) 
      -- CP-element group 120: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_698_Sample/ra
      -- CP-element group 120: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_698_Sample/$exit
      -- CP-element group 120: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_698_sample_completed_
      -- 
    ra_1594_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_698_inst_ack_0, ack => concat_CP_664_elements(120)); -- 
    -- CP-element group 121:  transition  input  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	277 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121:  members (3) 
      -- CP-element group 121: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_698_Update/$exit
      -- CP-element group 121: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_698_Update/ca
      -- CP-element group 121: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_698_update_completed_
      -- 
    ca_1599_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_698_inst_ack_1, ack => concat_CP_664_elements(121)); -- 
    -- CP-element group 122:  join  transition  output  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	89 
    -- CP-element group 122: 	93 
    -- CP-element group 122: 	97 
    -- CP-element group 122: 	101 
    -- CP-element group 122: 	105 
    -- CP-element group 122: 	109 
    -- CP-element group 122: 	113 
    -- CP-element group 122: 	117 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	123 
    -- CP-element group 122:  members (9) 
      -- CP-element group 122: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/ptr_deref_706_Sample/word_access_start/word_0/rr
      -- CP-element group 122: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/ptr_deref_706_Sample/ptr_deref_706_Split/split_ack
      -- CP-element group 122: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/ptr_deref_706_sample_start_
      -- CP-element group 122: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/ptr_deref_706_Sample/$entry
      -- CP-element group 122: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/ptr_deref_706_Sample/ptr_deref_706_Split/$entry
      -- CP-element group 122: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/ptr_deref_706_Sample/ptr_deref_706_Split/$exit
      -- CP-element group 122: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/ptr_deref_706_Sample/word_access_start/$entry
      -- CP-element group 122: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/ptr_deref_706_Sample/ptr_deref_706_Split/split_req
      -- CP-element group 122: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/ptr_deref_706_Sample/word_access_start/word_0/$entry
      -- 
    rr_1637_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1637_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(122), ack => ptr_deref_706_store_0_req_0); -- 
    concat_cp_element_group_122: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_122"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= concat_CP_664_elements(89) & concat_CP_664_elements(93) & concat_CP_664_elements(97) & concat_CP_664_elements(101) & concat_CP_664_elements(105) & concat_CP_664_elements(109) & concat_CP_664_elements(113) & concat_CP_664_elements(117) & concat_CP_664_elements(121);
      gj_concat_cp_element_group_122 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_664_elements(122), clk => clk, reset => reset); --
    end block;
    -- CP-element group 123:  transition  input  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	122 
    -- CP-element group 123: successors 
    -- CP-element group 123:  members (5) 
      -- CP-element group 123: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/ptr_deref_706_Sample/word_access_start/word_0/ra
      -- CP-element group 123: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/ptr_deref_706_Sample/$exit
      -- CP-element group 123: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/ptr_deref_706_Sample/word_access_start/word_0/$exit
      -- CP-element group 123: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/ptr_deref_706_sample_completed_
      -- CP-element group 123: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/ptr_deref_706_Sample/word_access_start/$exit
      -- 
    ra_1638_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_706_store_0_ack_0, ack => concat_CP_664_elements(123)); -- 
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	277 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	125 
    -- CP-element group 124:  members (5) 
      -- CP-element group 124: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/ptr_deref_706_update_completed_
      -- CP-element group 124: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/ptr_deref_706_Update/word_access_complete/$exit
      -- CP-element group 124: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/ptr_deref_706_Update/word_access_complete/word_0/$exit
      -- CP-element group 124: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/ptr_deref_706_Update/word_access_complete/word_0/ca
      -- CP-element group 124: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/ptr_deref_706_Update/$exit
      -- 
    ca_1649_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_706_store_0_ack_1, ack => concat_CP_664_elements(124)); -- 
    -- CP-element group 125:  branch  join  transition  place  output  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	86 
    -- CP-element group 125: 	124 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	126 
    -- CP-element group 125: 	127 
    -- CP-element group 125:  members (10) 
      -- CP-element group 125: 	 branch_block_stmt_216/if_stmt_720__entry__
      -- CP-element group 125: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719__exit__
      -- CP-element group 125: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/$exit
      -- CP-element group 125: 	 branch_block_stmt_216/if_stmt_720_dead_link/$entry
      -- CP-element group 125: 	 branch_block_stmt_216/if_stmt_720_eval_test/$entry
      -- CP-element group 125: 	 branch_block_stmt_216/if_stmt_720_eval_test/$exit
      -- CP-element group 125: 	 branch_block_stmt_216/if_stmt_720_eval_test/branch_req
      -- CP-element group 125: 	 branch_block_stmt_216/R_exitcond17_721_place
      -- CP-element group 125: 	 branch_block_stmt_216/if_stmt_720_if_link/$entry
      -- CP-element group 125: 	 branch_block_stmt_216/if_stmt_720_else_link/$entry
      -- 
    branch_req_1657_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1657_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(125), ack => if_stmt_720_branch_req_0); -- 
    concat_cp_element_group_125: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_125"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_664_elements(86) & concat_CP_664_elements(124);
      gj_concat_cp_element_group_125 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_664_elements(125), clk => clk, reset => reset); --
    end block;
    -- CP-element group 126:  merge  transition  place  input  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	125 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	271 
    -- CP-element group 126:  members (13) 
      -- CP-element group 126: 	 branch_block_stmt_216/merge_stmt_504__exit__
      -- CP-element group 126: 	 branch_block_stmt_216/forx_xcond165x_xpreheaderx_xloopexit_forx_xcond165x_xpreheader
      -- CP-element group 126: 	 branch_block_stmt_216/if_stmt_720_if_link/$exit
      -- CP-element group 126: 	 branch_block_stmt_216/if_stmt_720_if_link/if_choice_transition
      -- CP-element group 126: 	 branch_block_stmt_216/forx_xbody_forx_xcond165x_xpreheaderx_xloopexit
      -- CP-element group 126: 	 branch_block_stmt_216/forx_xbody_forx_xcond165x_xpreheaderx_xloopexit_PhiReq/$entry
      -- CP-element group 126: 	 branch_block_stmt_216/forx_xbody_forx_xcond165x_xpreheaderx_xloopexit_PhiReq/$exit
      -- CP-element group 126: 	 branch_block_stmt_216/merge_stmt_504_PhiReqMerge
      -- CP-element group 126: 	 branch_block_stmt_216/merge_stmt_504_PhiAck/$entry
      -- CP-element group 126: 	 branch_block_stmt_216/merge_stmt_504_PhiAck/$exit
      -- CP-element group 126: 	 branch_block_stmt_216/merge_stmt_504_PhiAck/dummy
      -- CP-element group 126: 	 branch_block_stmt_216/forx_xcond165x_xpreheaderx_xloopexit_forx_xcond165x_xpreheader_PhiReq/$entry
      -- CP-element group 126: 	 branch_block_stmt_216/forx_xcond165x_xpreheaderx_xloopexit_forx_xcond165x_xpreheader_PhiReq/$exit
      -- 
    if_choice_transition_1662_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_720_branch_ack_1, ack => concat_CP_664_elements(126)); -- 
    -- CP-element group 127:  fork  transition  place  input  output  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	125 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	273 
    -- CP-element group 127: 	274 
    -- CP-element group 127:  members (12) 
      -- CP-element group 127: 	 branch_block_stmt_216/if_stmt_720_else_link/$exit
      -- CP-element group 127: 	 branch_block_stmt_216/if_stmt_720_else_link/else_choice_transition
      -- CP-element group 127: 	 branch_block_stmt_216/forx_xbody_forx_xbody
      -- CP-element group 127: 	 branch_block_stmt_216/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 127: 	 branch_block_stmt_216/forx_xbody_forx_xbody_PhiReq/phi_stmt_555/$entry
      -- CP-element group 127: 	 branch_block_stmt_216/forx_xbody_forx_xbody_PhiReq/phi_stmt_555/phi_stmt_555_sources/$entry
      -- CP-element group 127: 	 branch_block_stmt_216/forx_xbody_forx_xbody_PhiReq/phi_stmt_555/phi_stmt_555_sources/type_cast_561/$entry
      -- CP-element group 127: 	 branch_block_stmt_216/forx_xbody_forx_xbody_PhiReq/phi_stmt_555/phi_stmt_555_sources/type_cast_561/SplitProtocol/$entry
      -- CP-element group 127: 	 branch_block_stmt_216/forx_xbody_forx_xbody_PhiReq/phi_stmt_555/phi_stmt_555_sources/type_cast_561/SplitProtocol/Sample/$entry
      -- CP-element group 127: 	 branch_block_stmt_216/forx_xbody_forx_xbody_PhiReq/phi_stmt_555/phi_stmt_555_sources/type_cast_561/SplitProtocol/Sample/rr
      -- CP-element group 127: 	 branch_block_stmt_216/forx_xbody_forx_xbody_PhiReq/phi_stmt_555/phi_stmt_555_sources/type_cast_561/SplitProtocol/Update/$entry
      -- CP-element group 127: 	 branch_block_stmt_216/forx_xbody_forx_xbody_PhiReq/phi_stmt_555/phi_stmt_555_sources/type_cast_561/SplitProtocol/Update/cr
      -- 
    else_choice_transition_1666_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_720_branch_ack_0, ack => concat_CP_664_elements(127)); -- 
    rr_2762_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2762_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(127), ack => type_cast_561_inst_req_0); -- 
    cr_2767_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2767_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(127), ack => type_cast_561_inst_req_1); -- 
    -- CP-element group 128:  transition  input  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	82 
    -- CP-element group 128: successors 
    -- CP-element group 128:  members (3) 
      -- CP-element group 128: 	 branch_block_stmt_216/assign_stmt_731_to_assign_stmt_759/type_cast_734_sample_completed_
      -- CP-element group 128: 	 branch_block_stmt_216/assign_stmt_731_to_assign_stmt_759/type_cast_734_Sample/$exit
      -- CP-element group 128: 	 branch_block_stmt_216/assign_stmt_731_to_assign_stmt_759/type_cast_734_Sample/ra
      -- 
    ra_1680_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_734_inst_ack_0, ack => concat_CP_664_elements(128)); -- 
    -- CP-element group 129:  transition  place  input  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	82 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	278 
    -- CP-element group 129:  members (9) 
      -- CP-element group 129: 	 branch_block_stmt_216/bbx_xnph386_forx_xbody171
      -- CP-element group 129: 	 branch_block_stmt_216/assign_stmt_731_to_assign_stmt_759__exit__
      -- CP-element group 129: 	 branch_block_stmt_216/assign_stmt_731_to_assign_stmt_759/$exit
      -- CP-element group 129: 	 branch_block_stmt_216/assign_stmt_731_to_assign_stmt_759/type_cast_734_update_completed_
      -- CP-element group 129: 	 branch_block_stmt_216/assign_stmt_731_to_assign_stmt_759/type_cast_734_Update/$exit
      -- CP-element group 129: 	 branch_block_stmt_216/assign_stmt_731_to_assign_stmt_759/type_cast_734_Update/ca
      -- CP-element group 129: 	 branch_block_stmt_216/bbx_xnph386_forx_xbody171_PhiReq/$entry
      -- CP-element group 129: 	 branch_block_stmt_216/bbx_xnph386_forx_xbody171_PhiReq/phi_stmt_762/$entry
      -- CP-element group 129: 	 branch_block_stmt_216/bbx_xnph386_forx_xbody171_PhiReq/phi_stmt_762/phi_stmt_762_sources/$entry
      -- 
    ca_1685_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_734_inst_ack_1, ack => concat_CP_664_elements(129)); -- 
    -- CP-element group 130:  transition  input  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	283 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	169 
    -- CP-element group 130:  members (3) 
      -- CP-element group 130: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/array_obj_ref_776_final_index_sum_regn_sample_complete
      -- CP-element group 130: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/array_obj_ref_776_final_index_sum_regn_Sample/$exit
      -- CP-element group 130: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/array_obj_ref_776_final_index_sum_regn_Sample/ack
      -- 
    ack_1714_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_776_index_offset_ack_0, ack => concat_CP_664_elements(130)); -- 
    -- CP-element group 131:  transition  input  output  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	283 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	132 
    -- CP-element group 131:  members (11) 
      -- CP-element group 131: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/addr_of_777_sample_start_
      -- CP-element group 131: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/array_obj_ref_776_root_address_calculated
      -- CP-element group 131: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/array_obj_ref_776_offset_calculated
      -- CP-element group 131: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/array_obj_ref_776_final_index_sum_regn_Update/$exit
      -- CP-element group 131: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/array_obj_ref_776_final_index_sum_regn_Update/ack
      -- CP-element group 131: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/array_obj_ref_776_base_plus_offset/$entry
      -- CP-element group 131: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/array_obj_ref_776_base_plus_offset/$exit
      -- CP-element group 131: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/array_obj_ref_776_base_plus_offset/sum_rename_req
      -- CP-element group 131: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/array_obj_ref_776_base_plus_offset/sum_rename_ack
      -- CP-element group 131: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/addr_of_777_request/$entry
      -- CP-element group 131: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/addr_of_777_request/req
      -- 
    ack_1719_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_776_index_offset_ack_1, ack => concat_CP_664_elements(131)); -- 
    req_1728_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1728_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(131), ack => addr_of_777_final_reg_req_0); -- 
    -- CP-element group 132:  transition  input  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	131 
    -- CP-element group 132: successors 
    -- CP-element group 132:  members (3) 
      -- CP-element group 132: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/addr_of_777_sample_completed_
      -- CP-element group 132: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/addr_of_777_request/$exit
      -- CP-element group 132: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/addr_of_777_request/ack
      -- 
    ack_1729_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_777_final_reg_ack_0, ack => concat_CP_664_elements(132)); -- 
    -- CP-element group 133:  fork  transition  input  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	283 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	166 
    -- CP-element group 133:  members (19) 
      -- CP-element group 133: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/addr_of_777_update_completed_
      -- CP-element group 133: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/addr_of_777_complete/$exit
      -- CP-element group 133: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/addr_of_777_complete/ack
      -- CP-element group 133: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_base_address_calculated
      -- CP-element group 133: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_word_address_calculated
      -- CP-element group 133: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_root_address_calculated
      -- CP-element group 133: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_base_address_resized
      -- CP-element group 133: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_base_addr_resize/$entry
      -- CP-element group 133: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_base_addr_resize/$exit
      -- CP-element group 133: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_base_addr_resize/base_resize_req
      -- CP-element group 133: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_base_addr_resize/base_resize_ack
      -- CP-element group 133: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_base_plus_offset/$entry
      -- CP-element group 133: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_base_plus_offset/$exit
      -- CP-element group 133: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_base_plus_offset/sum_rename_req
      -- CP-element group 133: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_base_plus_offset/sum_rename_ack
      -- CP-element group 133: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_word_addrgen/$entry
      -- CP-element group 133: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_word_addrgen/$exit
      -- CP-element group 133: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_word_addrgen/root_register_req
      -- CP-element group 133: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_word_addrgen/root_register_ack
      -- 
    ack_1734_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_777_final_reg_ack_1, ack => concat_CP_664_elements(133)); -- 
    -- CP-element group 134:  transition  input  output  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	283 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	135 
    -- CP-element group 134:  members (6) 
      -- CP-element group 134: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_780_sample_completed_
      -- CP-element group 134: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_780_update_start_
      -- CP-element group 134: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_780_Sample/$exit
      -- CP-element group 134: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_780_Sample/ra
      -- CP-element group 134: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_780_Update/$entry
      -- CP-element group 134: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_780_Update/cr
      -- 
    ra_1743_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_780_inst_ack_0, ack => concat_CP_664_elements(134)); -- 
    cr_1747_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1747_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(134), ack => RPIPE_Concat_input_pipe_780_inst_req_1); -- 
    -- CP-element group 135:  fork  transition  input  output  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	134 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	136 
    -- CP-element group 135: 	138 
    -- CP-element group 135:  members (9) 
      -- CP-element group 135: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_780_update_completed_
      -- CP-element group 135: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_780_Update/$exit
      -- CP-element group 135: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_780_Update/ca
      -- CP-element group 135: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_784_sample_start_
      -- CP-element group 135: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_784_Sample/$entry
      -- CP-element group 135: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_784_Sample/rr
      -- CP-element group 135: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_793_sample_start_
      -- CP-element group 135: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_793_Sample/$entry
      -- CP-element group 135: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_793_Sample/rr
      -- 
    ca_1748_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_780_inst_ack_1, ack => concat_CP_664_elements(135)); -- 
    rr_1756_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1756_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(135), ack => type_cast_784_inst_req_0); -- 
    rr_1770_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1770_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(135), ack => RPIPE_Concat_input_pipe_793_inst_req_0); -- 
    -- CP-element group 136:  transition  input  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	135 
    -- CP-element group 136: successors 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_784_sample_completed_
      -- CP-element group 136: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_784_Sample/$exit
      -- CP-element group 136: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_784_Sample/ra
      -- 
    ra_1757_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_784_inst_ack_0, ack => concat_CP_664_elements(136)); -- 
    -- CP-element group 137:  transition  input  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	283 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	166 
    -- CP-element group 137:  members (3) 
      -- CP-element group 137: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_784_update_completed_
      -- CP-element group 137: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_784_Update/$exit
      -- CP-element group 137: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_784_Update/ca
      -- 
    ca_1762_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_784_inst_ack_1, ack => concat_CP_664_elements(137)); -- 
    -- CP-element group 138:  transition  input  output  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	135 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	139 
    -- CP-element group 138:  members (6) 
      -- CP-element group 138: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_793_sample_completed_
      -- CP-element group 138: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_793_update_start_
      -- CP-element group 138: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_793_Sample/$exit
      -- CP-element group 138: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_793_Sample/ra
      -- CP-element group 138: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_793_Update/$entry
      -- CP-element group 138: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_793_Update/cr
      -- 
    ra_1771_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_793_inst_ack_0, ack => concat_CP_664_elements(138)); -- 
    cr_1775_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1775_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(138), ack => RPIPE_Concat_input_pipe_793_inst_req_1); -- 
    -- CP-element group 139:  fork  transition  input  output  bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	138 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	140 
    -- CP-element group 139: 	142 
    -- CP-element group 139:  members (9) 
      -- CP-element group 139: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_793_update_completed_
      -- CP-element group 139: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_793_Update/$exit
      -- CP-element group 139: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_793_Update/ca
      -- CP-element group 139: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_797_sample_start_
      -- CP-element group 139: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_797_Sample/$entry
      -- CP-element group 139: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_797_Sample/rr
      -- CP-element group 139: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_811_sample_start_
      -- CP-element group 139: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_811_Sample/$entry
      -- CP-element group 139: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_811_Sample/rr
      -- 
    ca_1776_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_793_inst_ack_1, ack => concat_CP_664_elements(139)); -- 
    rr_1784_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1784_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(139), ack => type_cast_797_inst_req_0); -- 
    rr_1798_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1798_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(139), ack => RPIPE_Concat_input_pipe_811_inst_req_0); -- 
    -- CP-element group 140:  transition  input  bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	139 
    -- CP-element group 140: successors 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_797_sample_completed_
      -- CP-element group 140: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_797_Sample/$exit
      -- CP-element group 140: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_797_Sample/ra
      -- 
    ra_1785_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_797_inst_ack_0, ack => concat_CP_664_elements(140)); -- 
    -- CP-element group 141:  transition  input  bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	283 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	166 
    -- CP-element group 141:  members (3) 
      -- CP-element group 141: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_797_update_completed_
      -- CP-element group 141: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_797_Update/$exit
      -- CP-element group 141: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_797_Update/ca
      -- 
    ca_1790_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_797_inst_ack_1, ack => concat_CP_664_elements(141)); -- 
    -- CP-element group 142:  transition  input  output  bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	139 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	143 
    -- CP-element group 142:  members (6) 
      -- CP-element group 142: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_811_sample_completed_
      -- CP-element group 142: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_811_update_start_
      -- CP-element group 142: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_811_Sample/$exit
      -- CP-element group 142: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_811_Sample/ra
      -- CP-element group 142: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_811_Update/$entry
      -- CP-element group 142: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_811_Update/cr
      -- 
    ra_1799_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_811_inst_ack_0, ack => concat_CP_664_elements(142)); -- 
    cr_1803_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1803_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(142), ack => RPIPE_Concat_input_pipe_811_inst_req_1); -- 
    -- CP-element group 143:  fork  transition  input  output  bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	142 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	144 
    -- CP-element group 143: 	146 
    -- CP-element group 143:  members (9) 
      -- CP-element group 143: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_811_update_completed_
      -- CP-element group 143: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_811_Update/$exit
      -- CP-element group 143: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_811_Update/ca
      -- CP-element group 143: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_815_sample_start_
      -- CP-element group 143: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_815_Sample/$entry
      -- CP-element group 143: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_815_Sample/rr
      -- CP-element group 143: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_829_sample_start_
      -- CP-element group 143: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_829_Sample/$entry
      -- CP-element group 143: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_829_Sample/rr
      -- 
    ca_1804_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_811_inst_ack_1, ack => concat_CP_664_elements(143)); -- 
    rr_1812_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1812_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(143), ack => type_cast_815_inst_req_0); -- 
    rr_1826_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1826_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(143), ack => RPIPE_Concat_input_pipe_829_inst_req_0); -- 
    -- CP-element group 144:  transition  input  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	143 
    -- CP-element group 144: successors 
    -- CP-element group 144:  members (3) 
      -- CP-element group 144: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_815_sample_completed_
      -- CP-element group 144: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_815_Sample/$exit
      -- CP-element group 144: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_815_Sample/ra
      -- 
    ra_1813_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_815_inst_ack_0, ack => concat_CP_664_elements(144)); -- 
    -- CP-element group 145:  transition  input  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	283 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	166 
    -- CP-element group 145:  members (3) 
      -- CP-element group 145: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_815_update_completed_
      -- CP-element group 145: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_815_Update/$exit
      -- CP-element group 145: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_815_Update/ca
      -- 
    ca_1818_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_815_inst_ack_1, ack => concat_CP_664_elements(145)); -- 
    -- CP-element group 146:  transition  input  output  bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	143 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	147 
    -- CP-element group 146:  members (6) 
      -- CP-element group 146: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_829_sample_completed_
      -- CP-element group 146: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_829_update_start_
      -- CP-element group 146: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_829_Sample/$exit
      -- CP-element group 146: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_829_Sample/ra
      -- CP-element group 146: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_829_Update/$entry
      -- CP-element group 146: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_829_Update/cr
      -- 
    ra_1827_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_829_inst_ack_0, ack => concat_CP_664_elements(146)); -- 
    cr_1831_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1831_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(146), ack => RPIPE_Concat_input_pipe_829_inst_req_1); -- 
    -- CP-element group 147:  fork  transition  input  output  bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	146 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	148 
    -- CP-element group 147: 	150 
    -- CP-element group 147:  members (9) 
      -- CP-element group 147: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_829_update_completed_
      -- CP-element group 147: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_829_Update/$exit
      -- CP-element group 147: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_829_Update/ca
      -- CP-element group 147: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_833_sample_start_
      -- CP-element group 147: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_833_Sample/$entry
      -- CP-element group 147: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_833_Sample/rr
      -- CP-element group 147: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_847_sample_start_
      -- CP-element group 147: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_847_Sample/$entry
      -- CP-element group 147: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_847_Sample/rr
      -- 
    ca_1832_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_829_inst_ack_1, ack => concat_CP_664_elements(147)); -- 
    rr_1840_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1840_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(147), ack => type_cast_833_inst_req_0); -- 
    rr_1854_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1854_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(147), ack => RPIPE_Concat_input_pipe_847_inst_req_0); -- 
    -- CP-element group 148:  transition  input  bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	147 
    -- CP-element group 148: successors 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_833_sample_completed_
      -- CP-element group 148: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_833_Sample/$exit
      -- CP-element group 148: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_833_Sample/ra
      -- 
    ra_1841_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_833_inst_ack_0, ack => concat_CP_664_elements(148)); -- 
    -- CP-element group 149:  transition  input  bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	283 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	166 
    -- CP-element group 149:  members (3) 
      -- CP-element group 149: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_833_update_completed_
      -- CP-element group 149: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_833_Update/$exit
      -- CP-element group 149: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_833_Update/ca
      -- 
    ca_1846_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_833_inst_ack_1, ack => concat_CP_664_elements(149)); -- 
    -- CP-element group 150:  transition  input  output  bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	147 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	151 
    -- CP-element group 150:  members (6) 
      -- CP-element group 150: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_847_sample_completed_
      -- CP-element group 150: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_847_update_start_
      -- CP-element group 150: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_847_Sample/$exit
      -- CP-element group 150: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_847_Sample/ra
      -- CP-element group 150: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_847_Update/$entry
      -- CP-element group 150: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_847_Update/cr
      -- 
    ra_1855_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_847_inst_ack_0, ack => concat_CP_664_elements(150)); -- 
    cr_1859_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1859_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(150), ack => RPIPE_Concat_input_pipe_847_inst_req_1); -- 
    -- CP-element group 151:  fork  transition  input  output  bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	150 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	152 
    -- CP-element group 151: 	154 
    -- CP-element group 151:  members (9) 
      -- CP-element group 151: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_847_update_completed_
      -- CP-element group 151: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_847_Update/$exit
      -- CP-element group 151: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_847_Update/ca
      -- CP-element group 151: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_851_sample_start_
      -- CP-element group 151: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_851_Sample/$entry
      -- CP-element group 151: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_851_Sample/rr
      -- CP-element group 151: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_865_sample_start_
      -- CP-element group 151: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_865_Sample/$entry
      -- CP-element group 151: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_865_Sample/rr
      -- 
    ca_1860_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_847_inst_ack_1, ack => concat_CP_664_elements(151)); -- 
    rr_1868_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1868_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(151), ack => type_cast_851_inst_req_0); -- 
    rr_1882_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1882_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(151), ack => RPIPE_Concat_input_pipe_865_inst_req_0); -- 
    -- CP-element group 152:  transition  input  bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	151 
    -- CP-element group 152: successors 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_851_sample_completed_
      -- CP-element group 152: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_851_Sample/$exit
      -- CP-element group 152: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_851_Sample/ra
      -- 
    ra_1869_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_851_inst_ack_0, ack => concat_CP_664_elements(152)); -- 
    -- CP-element group 153:  transition  input  bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	283 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	166 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_851_update_completed_
      -- CP-element group 153: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_851_Update/$exit
      -- CP-element group 153: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_851_Update/ca
      -- 
    ca_1874_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_851_inst_ack_1, ack => concat_CP_664_elements(153)); -- 
    -- CP-element group 154:  transition  input  output  bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	151 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	155 
    -- CP-element group 154:  members (6) 
      -- CP-element group 154: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_865_sample_completed_
      -- CP-element group 154: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_865_update_start_
      -- CP-element group 154: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_865_Sample/$exit
      -- CP-element group 154: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_865_Sample/ra
      -- CP-element group 154: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_865_Update/$entry
      -- CP-element group 154: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_865_Update/cr
      -- 
    ra_1883_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_865_inst_ack_0, ack => concat_CP_664_elements(154)); -- 
    cr_1887_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1887_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(154), ack => RPIPE_Concat_input_pipe_865_inst_req_1); -- 
    -- CP-element group 155:  fork  transition  input  output  bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	154 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	156 
    -- CP-element group 155: 	158 
    -- CP-element group 155:  members (9) 
      -- CP-element group 155: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_865_update_completed_
      -- CP-element group 155: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_865_Update/$exit
      -- CP-element group 155: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_865_Update/ca
      -- CP-element group 155: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_869_sample_start_
      -- CP-element group 155: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_869_Sample/$entry
      -- CP-element group 155: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_869_Sample/rr
      -- CP-element group 155: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_883_sample_start_
      -- CP-element group 155: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_883_Sample/$entry
      -- CP-element group 155: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_883_Sample/rr
      -- 
    ca_1888_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_865_inst_ack_1, ack => concat_CP_664_elements(155)); -- 
    rr_1896_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1896_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(155), ack => type_cast_869_inst_req_0); -- 
    rr_1910_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1910_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(155), ack => RPIPE_Concat_input_pipe_883_inst_req_0); -- 
    -- CP-element group 156:  transition  input  bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	155 
    -- CP-element group 156: successors 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_869_sample_completed_
      -- CP-element group 156: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_869_Sample/$exit
      -- CP-element group 156: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_869_Sample/ra
      -- 
    ra_1897_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_869_inst_ack_0, ack => concat_CP_664_elements(156)); -- 
    -- CP-element group 157:  transition  input  bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	283 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	166 
    -- CP-element group 157:  members (3) 
      -- CP-element group 157: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_869_update_completed_
      -- CP-element group 157: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_869_Update/$exit
      -- CP-element group 157: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_869_Update/ca
      -- 
    ca_1902_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_869_inst_ack_1, ack => concat_CP_664_elements(157)); -- 
    -- CP-element group 158:  transition  input  output  bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	155 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	159 
    -- CP-element group 158:  members (6) 
      -- CP-element group 158: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_883_sample_completed_
      -- CP-element group 158: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_883_update_start_
      -- CP-element group 158: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_883_Sample/$exit
      -- CP-element group 158: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_883_Sample/ra
      -- CP-element group 158: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_883_Update/$entry
      -- CP-element group 158: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_883_Update/cr
      -- 
    ra_1911_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_883_inst_ack_0, ack => concat_CP_664_elements(158)); -- 
    cr_1915_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1915_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(158), ack => RPIPE_Concat_input_pipe_883_inst_req_1); -- 
    -- CP-element group 159:  fork  transition  input  output  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	158 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	160 
    -- CP-element group 159: 	162 
    -- CP-element group 159:  members (9) 
      -- CP-element group 159: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_883_update_completed_
      -- CP-element group 159: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_883_Update/$exit
      -- CP-element group 159: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_883_Update/ca
      -- CP-element group 159: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_887_sample_start_
      -- CP-element group 159: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_887_Sample/$entry
      -- CP-element group 159: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_887_Sample/rr
      -- CP-element group 159: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_901_sample_start_
      -- CP-element group 159: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_901_Sample/$entry
      -- CP-element group 159: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_901_Sample/rr
      -- 
    ca_1916_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_883_inst_ack_1, ack => concat_CP_664_elements(159)); -- 
    rr_1924_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1924_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(159), ack => type_cast_887_inst_req_0); -- 
    rr_1938_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1938_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(159), ack => RPIPE_Concat_input_pipe_901_inst_req_0); -- 
    -- CP-element group 160:  transition  input  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	159 
    -- CP-element group 160: successors 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_887_sample_completed_
      -- CP-element group 160: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_887_Sample/$exit
      -- CP-element group 160: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_887_Sample/ra
      -- 
    ra_1925_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_887_inst_ack_0, ack => concat_CP_664_elements(160)); -- 
    -- CP-element group 161:  transition  input  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	283 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	166 
    -- CP-element group 161:  members (3) 
      -- CP-element group 161: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_887_update_completed_
      -- CP-element group 161: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_887_Update/$exit
      -- CP-element group 161: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_887_Update/ca
      -- 
    ca_1930_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_887_inst_ack_1, ack => concat_CP_664_elements(161)); -- 
    -- CP-element group 162:  transition  input  output  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	159 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	163 
    -- CP-element group 162:  members (6) 
      -- CP-element group 162: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_901_sample_completed_
      -- CP-element group 162: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_901_update_start_
      -- CP-element group 162: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_901_Sample/$exit
      -- CP-element group 162: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_901_Sample/ra
      -- CP-element group 162: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_901_Update/$entry
      -- CP-element group 162: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_901_Update/cr
      -- 
    ra_1939_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_901_inst_ack_0, ack => concat_CP_664_elements(162)); -- 
    cr_1943_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1943_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(162), ack => RPIPE_Concat_input_pipe_901_inst_req_1); -- 
    -- CP-element group 163:  transition  input  output  bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	162 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	164 
    -- CP-element group 163:  members (6) 
      -- CP-element group 163: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_901_update_completed_
      -- CP-element group 163: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_901_Update/$exit
      -- CP-element group 163: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_901_Update/ca
      -- CP-element group 163: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_905_sample_start_
      -- CP-element group 163: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_905_Sample/$entry
      -- CP-element group 163: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_905_Sample/rr
      -- 
    ca_1944_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Concat_input_pipe_901_inst_ack_1, ack => concat_CP_664_elements(163)); -- 
    rr_1952_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1952_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(163), ack => type_cast_905_inst_req_0); -- 
    -- CP-element group 164:  transition  input  bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	163 
    -- CP-element group 164: successors 
    -- CP-element group 164:  members (3) 
      -- CP-element group 164: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_905_sample_completed_
      -- CP-element group 164: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_905_Sample/$exit
      -- CP-element group 164: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_905_Sample/ra
      -- 
    ra_1953_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_905_inst_ack_0, ack => concat_CP_664_elements(164)); -- 
    -- CP-element group 165:  transition  input  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	283 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	166 
    -- CP-element group 165:  members (3) 
      -- CP-element group 165: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_905_update_completed_
      -- CP-element group 165: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_905_Update/$exit
      -- CP-element group 165: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_905_Update/ca
      -- 
    ca_1958_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_905_inst_ack_1, ack => concat_CP_664_elements(165)); -- 
    -- CP-element group 166:  join  transition  output  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	133 
    -- CP-element group 166: 	137 
    -- CP-element group 166: 	141 
    -- CP-element group 166: 	145 
    -- CP-element group 166: 	149 
    -- CP-element group 166: 	153 
    -- CP-element group 166: 	157 
    -- CP-element group 166: 	161 
    -- CP-element group 166: 	165 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	167 
    -- CP-element group 166:  members (9) 
      -- CP-element group 166: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_sample_start_
      -- CP-element group 166: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_Sample/$entry
      -- CP-element group 166: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_Sample/ptr_deref_913_Split/$entry
      -- CP-element group 166: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_Sample/ptr_deref_913_Split/$exit
      -- CP-element group 166: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_Sample/ptr_deref_913_Split/split_req
      -- CP-element group 166: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_Sample/ptr_deref_913_Split/split_ack
      -- CP-element group 166: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_Sample/word_access_start/$entry
      -- CP-element group 166: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_Sample/word_access_start/word_0/$entry
      -- CP-element group 166: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_Sample/word_access_start/word_0/rr
      -- 
    rr_1996_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1996_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(166), ack => ptr_deref_913_store_0_req_0); -- 
    concat_cp_element_group_166: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_166"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= concat_CP_664_elements(133) & concat_CP_664_elements(137) & concat_CP_664_elements(141) & concat_CP_664_elements(145) & concat_CP_664_elements(149) & concat_CP_664_elements(153) & concat_CP_664_elements(157) & concat_CP_664_elements(161) & concat_CP_664_elements(165);
      gj_concat_cp_element_group_166 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_664_elements(166), clk => clk, reset => reset); --
    end block;
    -- CP-element group 167:  transition  input  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	166 
    -- CP-element group 167: successors 
    -- CP-element group 167:  members (5) 
      -- CP-element group 167: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_sample_completed_
      -- CP-element group 167: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_Sample/$exit
      -- CP-element group 167: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_Sample/word_access_start/$exit
      -- CP-element group 167: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_Sample/word_access_start/word_0/$exit
      -- CP-element group 167: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_Sample/word_access_start/word_0/ra
      -- 
    ra_1997_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_913_store_0_ack_0, ack => concat_CP_664_elements(167)); -- 
    -- CP-element group 168:  transition  input  bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	283 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	169 
    -- CP-element group 168:  members (5) 
      -- CP-element group 168: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_update_completed_
      -- CP-element group 168: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_Update/$exit
      -- CP-element group 168: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_Update/word_access_complete/$exit
      -- CP-element group 168: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_Update/word_access_complete/word_0/$exit
      -- CP-element group 168: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_Update/word_access_complete/word_0/ca
      -- 
    ca_2008_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_913_store_0_ack_1, ack => concat_CP_664_elements(168)); -- 
    -- CP-element group 169:  branch  join  transition  place  output  bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	130 
    -- CP-element group 169: 	168 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	170 
    -- CP-element group 169: 	171 
    -- CP-element group 169:  members (10) 
      -- CP-element group 169: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926__exit__
      -- CP-element group 169: 	 branch_block_stmt_216/if_stmt_927__entry__
      -- CP-element group 169: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/$exit
      -- CP-element group 169: 	 branch_block_stmt_216/if_stmt_927_dead_link/$entry
      -- CP-element group 169: 	 branch_block_stmt_216/if_stmt_927_eval_test/$entry
      -- CP-element group 169: 	 branch_block_stmt_216/if_stmt_927_eval_test/$exit
      -- CP-element group 169: 	 branch_block_stmt_216/if_stmt_927_eval_test/branch_req
      -- CP-element group 169: 	 branch_block_stmt_216/R_exitcond_928_place
      -- CP-element group 169: 	 branch_block_stmt_216/if_stmt_927_if_link/$entry
      -- CP-element group 169: 	 branch_block_stmt_216/if_stmt_927_else_link/$entry
      -- 
    branch_req_2016_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2016_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(169), ack => if_stmt_927_branch_req_0); -- 
    concat_cp_element_group_169: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_169"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_664_elements(130) & concat_CP_664_elements(168);
      gj_concat_cp_element_group_169 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_664_elements(169), clk => clk, reset => reset); --
    end block;
    -- CP-element group 170:  merge  transition  place  input  bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	169 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	284 
    -- CP-element group 170:  members (13) 
      -- CP-element group 170: 	 branch_block_stmt_216/merge_stmt_933__exit__
      -- CP-element group 170: 	 branch_block_stmt_216/forx_xend224x_xloopexit_forx_xend224
      -- CP-element group 170: 	 branch_block_stmt_216/if_stmt_927_if_link/$exit
      -- CP-element group 170: 	 branch_block_stmt_216/if_stmt_927_if_link/if_choice_transition
      -- CP-element group 170: 	 branch_block_stmt_216/forx_xbody171_forx_xend224x_xloopexit
      -- CP-element group 170: 	 branch_block_stmt_216/forx_xbody171_forx_xend224x_xloopexit_PhiReq/$entry
      -- CP-element group 170: 	 branch_block_stmt_216/forx_xbody171_forx_xend224x_xloopexit_PhiReq/$exit
      -- CP-element group 170: 	 branch_block_stmt_216/merge_stmt_933_PhiReqMerge
      -- CP-element group 170: 	 branch_block_stmt_216/merge_stmt_933_PhiAck/$entry
      -- CP-element group 170: 	 branch_block_stmt_216/merge_stmt_933_PhiAck/$exit
      -- CP-element group 170: 	 branch_block_stmt_216/merge_stmt_933_PhiAck/dummy
      -- CP-element group 170: 	 branch_block_stmt_216/forx_xend224x_xloopexit_forx_xend224_PhiReq/$entry
      -- CP-element group 170: 	 branch_block_stmt_216/forx_xend224x_xloopexit_forx_xend224_PhiReq/$exit
      -- 
    if_choice_transition_2021_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_927_branch_ack_1, ack => concat_CP_664_elements(170)); -- 
    -- CP-element group 171:  fork  transition  place  input  output  bypass 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	169 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	279 
    -- CP-element group 171: 	280 
    -- CP-element group 171:  members (12) 
      -- CP-element group 171: 	 branch_block_stmt_216/if_stmt_927_else_link/$exit
      -- CP-element group 171: 	 branch_block_stmt_216/if_stmt_927_else_link/else_choice_transition
      -- CP-element group 171: 	 branch_block_stmt_216/forx_xbody171_forx_xbody171
      -- CP-element group 171: 	 branch_block_stmt_216/forx_xbody171_forx_xbody171_PhiReq/$entry
      -- CP-element group 171: 	 branch_block_stmt_216/forx_xbody171_forx_xbody171_PhiReq/phi_stmt_762/$entry
      -- CP-element group 171: 	 branch_block_stmt_216/forx_xbody171_forx_xbody171_PhiReq/phi_stmt_762/phi_stmt_762_sources/$entry
      -- CP-element group 171: 	 branch_block_stmt_216/forx_xbody171_forx_xbody171_PhiReq/phi_stmt_762/phi_stmt_762_sources/type_cast_768/$entry
      -- CP-element group 171: 	 branch_block_stmt_216/forx_xbody171_forx_xbody171_PhiReq/phi_stmt_762/phi_stmt_762_sources/type_cast_768/SplitProtocol/$entry
      -- CP-element group 171: 	 branch_block_stmt_216/forx_xbody171_forx_xbody171_PhiReq/phi_stmt_762/phi_stmt_762_sources/type_cast_768/SplitProtocol/Sample/$entry
      -- CP-element group 171: 	 branch_block_stmt_216/forx_xbody171_forx_xbody171_PhiReq/phi_stmt_762/phi_stmt_762_sources/type_cast_768/SplitProtocol/Sample/rr
      -- CP-element group 171: 	 branch_block_stmt_216/forx_xbody171_forx_xbody171_PhiReq/phi_stmt_762/phi_stmt_762_sources/type_cast_768/SplitProtocol/Update/$entry
      -- CP-element group 171: 	 branch_block_stmt_216/forx_xbody171_forx_xbody171_PhiReq/phi_stmt_762/phi_stmt_762_sources/type_cast_768/SplitProtocol/Update/cr
      -- 
    else_choice_transition_2025_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_927_branch_ack_0, ack => concat_CP_664_elements(171)); -- 
    rr_2816_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2816_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(171), ack => type_cast_768_inst_req_0); -- 
    cr_2821_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2821_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(171), ack => type_cast_768_inst_req_1); -- 
    -- CP-element group 172:  transition  input  bypass 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	284 
    -- CP-element group 172: successors 
    -- CP-element group 172:  members (3) 
      -- CP-element group 172: 	 branch_block_stmt_216/call_stmt_938_to_assign_stmt_944/call_stmt_938_sample_completed_
      -- CP-element group 172: 	 branch_block_stmt_216/call_stmt_938_to_assign_stmt_944/call_stmt_938_Sample/$exit
      -- CP-element group 172: 	 branch_block_stmt_216/call_stmt_938_to_assign_stmt_944/call_stmt_938_Sample/cra
      -- 
    cra_2039_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_938_call_ack_0, ack => concat_CP_664_elements(172)); -- 
    -- CP-element group 173:  transition  input  output  bypass 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	284 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	174 
    -- CP-element group 173:  members (6) 
      -- CP-element group 173: 	 branch_block_stmt_216/call_stmt_938_to_assign_stmt_944/call_stmt_938_update_completed_
      -- CP-element group 173: 	 branch_block_stmt_216/call_stmt_938_to_assign_stmt_944/call_stmt_938_Update/$exit
      -- CP-element group 173: 	 branch_block_stmt_216/call_stmt_938_to_assign_stmt_944/call_stmt_938_Update/cca
      -- CP-element group 173: 	 branch_block_stmt_216/call_stmt_938_to_assign_stmt_944/type_cast_943_sample_start_
      -- CP-element group 173: 	 branch_block_stmt_216/call_stmt_938_to_assign_stmt_944/type_cast_943_Sample/$entry
      -- CP-element group 173: 	 branch_block_stmt_216/call_stmt_938_to_assign_stmt_944/type_cast_943_Sample/rr
      -- 
    cca_2044_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_938_call_ack_1, ack => concat_CP_664_elements(173)); -- 
    rr_2052_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2052_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(173), ack => type_cast_943_inst_req_0); -- 
    -- CP-element group 174:  transition  input  bypass 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	173 
    -- CP-element group 174: successors 
    -- CP-element group 174:  members (3) 
      -- CP-element group 174: 	 branch_block_stmt_216/call_stmt_938_to_assign_stmt_944/type_cast_943_sample_completed_
      -- CP-element group 174: 	 branch_block_stmt_216/call_stmt_938_to_assign_stmt_944/type_cast_943_Sample/$exit
      -- CP-element group 174: 	 branch_block_stmt_216/call_stmt_938_to_assign_stmt_944/type_cast_943_Sample/ra
      -- 
    ra_2053_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_943_inst_ack_0, ack => concat_CP_664_elements(174)); -- 
    -- CP-element group 175:  fork  transition  place  input  output  bypass 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	284 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	176 
    -- CP-element group 175: 	177 
    -- CP-element group 175:  members (13) 
      -- CP-element group 175: 	 branch_block_stmt_216/call_stmt_938_to_assign_stmt_944__exit__
      -- CP-element group 175: 	 branch_block_stmt_216/call_stmt_949__entry__
      -- CP-element group 175: 	 branch_block_stmt_216/call_stmt_938_to_assign_stmt_944/$exit
      -- CP-element group 175: 	 branch_block_stmt_216/call_stmt_938_to_assign_stmt_944/type_cast_943_update_completed_
      -- CP-element group 175: 	 branch_block_stmt_216/call_stmt_938_to_assign_stmt_944/type_cast_943_Update/$exit
      -- CP-element group 175: 	 branch_block_stmt_216/call_stmt_938_to_assign_stmt_944/type_cast_943_Update/ca
      -- CP-element group 175: 	 branch_block_stmt_216/call_stmt_949/$entry
      -- CP-element group 175: 	 branch_block_stmt_216/call_stmt_949/call_stmt_949_sample_start_
      -- CP-element group 175: 	 branch_block_stmt_216/call_stmt_949/call_stmt_949_update_start_
      -- CP-element group 175: 	 branch_block_stmt_216/call_stmt_949/call_stmt_949_Sample/$entry
      -- CP-element group 175: 	 branch_block_stmt_216/call_stmt_949/call_stmt_949_Sample/crr
      -- CP-element group 175: 	 branch_block_stmt_216/call_stmt_949/call_stmt_949_Update/$entry
      -- CP-element group 175: 	 branch_block_stmt_216/call_stmt_949/call_stmt_949_Update/ccr
      -- 
    ca_2058_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_943_inst_ack_1, ack => concat_CP_664_elements(175)); -- 
    crr_2069_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2069_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(175), ack => call_stmt_949_call_req_0); -- 
    ccr_2074_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2074_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(175), ack => call_stmt_949_call_req_1); -- 
    -- CP-element group 176:  transition  input  bypass 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	175 
    -- CP-element group 176: successors 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 branch_block_stmt_216/call_stmt_949/call_stmt_949_sample_completed_
      -- CP-element group 176: 	 branch_block_stmt_216/call_stmt_949/call_stmt_949_Sample/$exit
      -- CP-element group 176: 	 branch_block_stmt_216/call_stmt_949/call_stmt_949_Sample/cra
      -- 
    cra_2070_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_949_call_ack_0, ack => concat_CP_664_elements(176)); -- 
    -- CP-element group 177:  fork  transition  place  input  output  bypass 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	175 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	178 
    -- CP-element group 177: 	179 
    -- CP-element group 177: 	181 
    -- CP-element group 177: 	183 
    -- CP-element group 177: 	185 
    -- CP-element group 177: 	187 
    -- CP-element group 177: 	189 
    -- CP-element group 177: 	191 
    -- CP-element group 177: 	193 
    -- CP-element group 177: 	195 
    -- CP-element group 177: 	197 
    -- CP-element group 177:  members (40) 
      -- CP-element group 177: 	 branch_block_stmt_216/call_stmt_949__exit__
      -- CP-element group 177: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060__entry__
      -- CP-element group 177: 	 branch_block_stmt_216/call_stmt_949/$exit
      -- CP-element group 177: 	 branch_block_stmt_216/call_stmt_949/call_stmt_949_update_completed_
      -- CP-element group 177: 	 branch_block_stmt_216/call_stmt_949/call_stmt_949_Update/$exit
      -- CP-element group 177: 	 branch_block_stmt_216/call_stmt_949/call_stmt_949_Update/cca
      -- CP-element group 177: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/$entry
      -- CP-element group 177: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/call_stmt_952_sample_start_
      -- CP-element group 177: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/call_stmt_952_update_start_
      -- CP-element group 177: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/call_stmt_952_Sample/$entry
      -- CP-element group 177: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/call_stmt_952_Sample/crr
      -- CP-element group 177: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/call_stmt_952_Update/$entry
      -- CP-element group 177: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/call_stmt_952_Update/ccr
      -- CP-element group 177: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_956_update_start_
      -- CP-element group 177: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_956_Update/$entry
      -- CP-element group 177: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_956_Update/cr
      -- CP-element group 177: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_965_update_start_
      -- CP-element group 177: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_965_Update/$entry
      -- CP-element group 177: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_965_Update/cr
      -- CP-element group 177: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_975_update_start_
      -- CP-element group 177: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_975_Update/$entry
      -- CP-element group 177: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_975_Update/cr
      -- CP-element group 177: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_985_update_start_
      -- CP-element group 177: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_985_Update/$entry
      -- CP-element group 177: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_985_Update/cr
      -- CP-element group 177: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_995_update_start_
      -- CP-element group 177: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_995_Update/$entry
      -- CP-element group 177: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_995_Update/cr
      -- CP-element group 177: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_1005_update_start_
      -- CP-element group 177: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_1005_Update/$entry
      -- CP-element group 177: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_1005_Update/cr
      -- CP-element group 177: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_1015_update_start_
      -- CP-element group 177: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_1015_Update/$entry
      -- CP-element group 177: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_1015_Update/cr
      -- CP-element group 177: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_1025_update_start_
      -- CP-element group 177: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_1025_Update/$entry
      -- CP-element group 177: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_1025_Update/cr
      -- CP-element group 177: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_1035_update_start_
      -- CP-element group 177: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_1035_Update/$entry
      -- CP-element group 177: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_1035_Update/cr
      -- 
    cca_2075_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_949_call_ack_1, ack => concat_CP_664_elements(177)); -- 
    crr_2086_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2086_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(177), ack => call_stmt_952_call_req_0); -- 
    ccr_2091_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2091_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(177), ack => call_stmt_952_call_req_1); -- 
    cr_2105_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2105_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(177), ack => type_cast_956_inst_req_1); -- 
    cr_2119_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2119_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(177), ack => type_cast_965_inst_req_1); -- 
    cr_2133_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2133_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(177), ack => type_cast_975_inst_req_1); -- 
    cr_2147_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2147_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(177), ack => type_cast_985_inst_req_1); -- 
    cr_2161_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2161_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(177), ack => type_cast_995_inst_req_1); -- 
    cr_2175_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2175_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(177), ack => type_cast_1005_inst_req_1); -- 
    cr_2189_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2189_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(177), ack => type_cast_1015_inst_req_1); -- 
    cr_2203_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2203_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(177), ack => type_cast_1025_inst_req_1); -- 
    cr_2217_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2217_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(177), ack => type_cast_1035_inst_req_1); -- 
    -- CP-element group 178:  transition  input  bypass 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	177 
    -- CP-element group 178: successors 
    -- CP-element group 178:  members (3) 
      -- CP-element group 178: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/call_stmt_952_sample_completed_
      -- CP-element group 178: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/call_stmt_952_Sample/$exit
      -- CP-element group 178: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/call_stmt_952_Sample/cra
      -- 
    cra_2087_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_952_call_ack_0, ack => concat_CP_664_elements(178)); -- 
    -- CP-element group 179:  transition  input  output  bypass 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	177 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	180 
    -- CP-element group 179:  members (6) 
      -- CP-element group 179: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/call_stmt_952_update_completed_
      -- CP-element group 179: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/call_stmt_952_Update/$exit
      -- CP-element group 179: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/call_stmt_952_Update/cca
      -- CP-element group 179: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_956_sample_start_
      -- CP-element group 179: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_956_Sample/$entry
      -- CP-element group 179: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_956_Sample/rr
      -- 
    cca_2092_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_952_call_ack_1, ack => concat_CP_664_elements(179)); -- 
    rr_2100_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2100_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(179), ack => type_cast_956_inst_req_0); -- 
    -- CP-element group 180:  transition  input  bypass 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	179 
    -- CP-element group 180: successors 
    -- CP-element group 180:  members (3) 
      -- CP-element group 180: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_956_sample_completed_
      -- CP-element group 180: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_956_Sample/$exit
      -- CP-element group 180: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_956_Sample/ra
      -- 
    ra_2101_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_956_inst_ack_0, ack => concat_CP_664_elements(180)); -- 
    -- CP-element group 181:  fork  transition  input  output  bypass 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	177 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	182 
    -- CP-element group 181: 	184 
    -- CP-element group 181: 	186 
    -- CP-element group 181: 	188 
    -- CP-element group 181: 	190 
    -- CP-element group 181: 	192 
    -- CP-element group 181: 	194 
    -- CP-element group 181: 	196 
    -- CP-element group 181:  members (27) 
      -- CP-element group 181: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_956_update_completed_
      -- CP-element group 181: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_956_Update/$exit
      -- CP-element group 181: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_956_Update/ca
      -- CP-element group 181: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_965_sample_start_
      -- CP-element group 181: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_965_Sample/$entry
      -- CP-element group 181: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_965_Sample/rr
      -- CP-element group 181: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_975_sample_start_
      -- CP-element group 181: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_975_Sample/$entry
      -- CP-element group 181: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_975_Sample/rr
      -- CP-element group 181: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_985_sample_start_
      -- CP-element group 181: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_985_Sample/$entry
      -- CP-element group 181: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_985_Sample/rr
      -- CP-element group 181: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_995_sample_start_
      -- CP-element group 181: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_995_Sample/$entry
      -- CP-element group 181: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_995_Sample/rr
      -- CP-element group 181: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_1005_sample_start_
      -- CP-element group 181: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_1005_Sample/$entry
      -- CP-element group 181: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_1005_Sample/rr
      -- CP-element group 181: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_1015_sample_start_
      -- CP-element group 181: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_1015_Sample/$entry
      -- CP-element group 181: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_1015_Sample/rr
      -- CP-element group 181: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_1025_sample_start_
      -- CP-element group 181: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_1025_Sample/$entry
      -- CP-element group 181: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_1025_Sample/rr
      -- CP-element group 181: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_1035_sample_start_
      -- CP-element group 181: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_1035_Sample/$entry
      -- CP-element group 181: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_1035_Sample/rr
      -- 
    ca_2106_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_956_inst_ack_1, ack => concat_CP_664_elements(181)); -- 
    rr_2114_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2114_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(181), ack => type_cast_965_inst_req_0); -- 
    rr_2128_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2128_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(181), ack => type_cast_975_inst_req_0); -- 
    rr_2142_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2142_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(181), ack => type_cast_985_inst_req_0); -- 
    rr_2156_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2156_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(181), ack => type_cast_995_inst_req_0); -- 
    rr_2170_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2170_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(181), ack => type_cast_1005_inst_req_0); -- 
    rr_2184_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2184_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(181), ack => type_cast_1015_inst_req_0); -- 
    rr_2198_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2198_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(181), ack => type_cast_1025_inst_req_0); -- 
    rr_2212_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2212_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(181), ack => type_cast_1035_inst_req_0); -- 
    -- CP-element group 182:  transition  input  bypass 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	181 
    -- CP-element group 182: successors 
    -- CP-element group 182:  members (3) 
      -- CP-element group 182: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_965_sample_completed_
      -- CP-element group 182: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_965_Sample/$exit
      -- CP-element group 182: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_965_Sample/ra
      -- 
    ra_2115_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_965_inst_ack_0, ack => concat_CP_664_elements(182)); -- 
    -- CP-element group 183:  transition  input  bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	177 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	218 
    -- CP-element group 183:  members (3) 
      -- CP-element group 183: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_965_update_completed_
      -- CP-element group 183: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_965_Update/$exit
      -- CP-element group 183: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_965_Update/ca
      -- 
    ca_2120_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_965_inst_ack_1, ack => concat_CP_664_elements(183)); -- 
    -- CP-element group 184:  transition  input  bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	181 
    -- CP-element group 184: successors 
    -- CP-element group 184:  members (3) 
      -- CP-element group 184: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_975_sample_completed_
      -- CP-element group 184: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_975_Sample/$exit
      -- CP-element group 184: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_975_Sample/ra
      -- 
    ra_2129_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_975_inst_ack_0, ack => concat_CP_664_elements(184)); -- 
    -- CP-element group 185:  transition  input  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	177 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	215 
    -- CP-element group 185:  members (3) 
      -- CP-element group 185: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_975_update_completed_
      -- CP-element group 185: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_975_Update/$exit
      -- CP-element group 185: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_975_Update/ca
      -- 
    ca_2134_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_975_inst_ack_1, ack => concat_CP_664_elements(185)); -- 
    -- CP-element group 186:  transition  input  bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	181 
    -- CP-element group 186: successors 
    -- CP-element group 186:  members (3) 
      -- CP-element group 186: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_985_sample_completed_
      -- CP-element group 186: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_985_Sample/$exit
      -- CP-element group 186: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_985_Sample/ra
      -- 
    ra_2143_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_985_inst_ack_0, ack => concat_CP_664_elements(186)); -- 
    -- CP-element group 187:  transition  input  bypass 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	177 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	212 
    -- CP-element group 187:  members (3) 
      -- CP-element group 187: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_985_update_completed_
      -- CP-element group 187: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_985_Update/$exit
      -- CP-element group 187: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_985_Update/ca
      -- 
    ca_2148_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_985_inst_ack_1, ack => concat_CP_664_elements(187)); -- 
    -- CP-element group 188:  transition  input  bypass 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	181 
    -- CP-element group 188: successors 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_995_sample_completed_
      -- CP-element group 188: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_995_Sample/$exit
      -- CP-element group 188: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_995_Sample/ra
      -- 
    ra_2157_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_995_inst_ack_0, ack => concat_CP_664_elements(188)); -- 
    -- CP-element group 189:  transition  input  bypass 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	177 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	209 
    -- CP-element group 189:  members (3) 
      -- CP-element group 189: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_995_update_completed_
      -- CP-element group 189: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_995_Update/$exit
      -- CP-element group 189: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_995_Update/ca
      -- 
    ca_2162_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_995_inst_ack_1, ack => concat_CP_664_elements(189)); -- 
    -- CP-element group 190:  transition  input  bypass 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	181 
    -- CP-element group 190: successors 
    -- CP-element group 190:  members (3) 
      -- CP-element group 190: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_1005_sample_completed_
      -- CP-element group 190: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_1005_Sample/$exit
      -- CP-element group 190: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_1005_Sample/ra
      -- 
    ra_2171_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1005_inst_ack_0, ack => concat_CP_664_elements(190)); -- 
    -- CP-element group 191:  transition  input  bypass 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	177 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	206 
    -- CP-element group 191:  members (3) 
      -- CP-element group 191: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_1005_update_completed_
      -- CP-element group 191: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_1005_Update/$exit
      -- CP-element group 191: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_1005_Update/ca
      -- 
    ca_2176_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1005_inst_ack_1, ack => concat_CP_664_elements(191)); -- 
    -- CP-element group 192:  transition  input  bypass 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	181 
    -- CP-element group 192: successors 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_1015_sample_completed_
      -- CP-element group 192: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_1015_Sample/$exit
      -- CP-element group 192: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_1015_Sample/ra
      -- 
    ra_2185_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1015_inst_ack_0, ack => concat_CP_664_elements(192)); -- 
    -- CP-element group 193:  transition  input  bypass 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	177 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	203 
    -- CP-element group 193:  members (3) 
      -- CP-element group 193: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_1015_update_completed_
      -- CP-element group 193: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_1015_Update/$exit
      -- CP-element group 193: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_1015_Update/ca
      -- 
    ca_2190_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1015_inst_ack_1, ack => concat_CP_664_elements(193)); -- 
    -- CP-element group 194:  transition  input  bypass 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	181 
    -- CP-element group 194: successors 
    -- CP-element group 194:  members (3) 
      -- CP-element group 194: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_1025_sample_completed_
      -- CP-element group 194: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_1025_Sample/$exit
      -- CP-element group 194: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_1025_Sample/ra
      -- 
    ra_2199_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1025_inst_ack_0, ack => concat_CP_664_elements(194)); -- 
    -- CP-element group 195:  transition  input  bypass 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	177 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	200 
    -- CP-element group 195:  members (3) 
      -- CP-element group 195: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_1025_update_completed_
      -- CP-element group 195: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_1025_Update/$exit
      -- CP-element group 195: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_1025_Update/ca
      -- 
    ca_2204_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1025_inst_ack_1, ack => concat_CP_664_elements(195)); -- 
    -- CP-element group 196:  transition  input  bypass 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	181 
    -- CP-element group 196: successors 
    -- CP-element group 196:  members (3) 
      -- CP-element group 196: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_1035_sample_completed_
      -- CP-element group 196: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_1035_Sample/$exit
      -- CP-element group 196: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_1035_Sample/ra
      -- 
    ra_2213_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1035_inst_ack_0, ack => concat_CP_664_elements(196)); -- 
    -- CP-element group 197:  transition  input  output  bypass 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	177 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	198 
    -- CP-element group 197:  members (6) 
      -- CP-element group 197: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_1035_update_completed_
      -- CP-element group 197: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_1035_Update/$exit
      -- CP-element group 197: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/type_cast_1035_Update/ca
      -- CP-element group 197: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1037_sample_start_
      -- CP-element group 197: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1037_Sample/$entry
      -- CP-element group 197: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1037_Sample/req
      -- 
    ca_2218_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1035_inst_ack_1, ack => concat_CP_664_elements(197)); -- 
    req_2226_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2226_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(197), ack => WPIPE_Concat_output_pipe_1037_inst_req_0); -- 
    -- CP-element group 198:  transition  input  output  bypass 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	197 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	199 
    -- CP-element group 198:  members (6) 
      -- CP-element group 198: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1037_Update/req
      -- CP-element group 198: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1037_Update/$entry
      -- CP-element group 198: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1037_sample_completed_
      -- CP-element group 198: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1037_update_start_
      -- CP-element group 198: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1037_Sample/$exit
      -- CP-element group 198: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1037_Sample/ack
      -- 
    ack_2227_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1037_inst_ack_0, ack => concat_CP_664_elements(198)); -- 
    req_2231_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2231_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(198), ack => WPIPE_Concat_output_pipe_1037_inst_req_1); -- 
    -- CP-element group 199:  transition  input  bypass 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	198 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	200 
    -- CP-element group 199:  members (3) 
      -- CP-element group 199: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1037_Update/ack
      -- CP-element group 199: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1037_Update/$exit
      -- CP-element group 199: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1037_update_completed_
      -- 
    ack_2232_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1037_inst_ack_1, ack => concat_CP_664_elements(199)); -- 
    -- CP-element group 200:  join  transition  output  bypass 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	195 
    -- CP-element group 200: 	199 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	201 
    -- CP-element group 200:  members (3) 
      -- CP-element group 200: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1040_Sample/$entry
      -- CP-element group 200: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1040_Sample/req
      -- CP-element group 200: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1040_sample_start_
      -- 
    req_2240_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2240_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(200), ack => WPIPE_Concat_output_pipe_1040_inst_req_0); -- 
    concat_cp_element_group_200: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_200"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_664_elements(195) & concat_CP_664_elements(199);
      gj_concat_cp_element_group_200 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_664_elements(200), clk => clk, reset => reset); --
    end block;
    -- CP-element group 201:  transition  input  output  bypass 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	200 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	202 
    -- CP-element group 201:  members (6) 
      -- CP-element group 201: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1040_sample_completed_
      -- CP-element group 201: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1040_update_start_
      -- CP-element group 201: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1040_Sample/$exit
      -- CP-element group 201: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1040_Update/req
      -- CP-element group 201: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1040_Update/$entry
      -- CP-element group 201: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1040_Sample/ack
      -- 
    ack_2241_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1040_inst_ack_0, ack => concat_CP_664_elements(201)); -- 
    req_2245_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2245_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(201), ack => WPIPE_Concat_output_pipe_1040_inst_req_1); -- 
    -- CP-element group 202:  transition  input  bypass 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	201 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	203 
    -- CP-element group 202:  members (3) 
      -- CP-element group 202: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1040_update_completed_
      -- CP-element group 202: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1040_Update/ack
      -- CP-element group 202: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1040_Update/$exit
      -- 
    ack_2246_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1040_inst_ack_1, ack => concat_CP_664_elements(202)); -- 
    -- CP-element group 203:  join  transition  output  bypass 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	193 
    -- CP-element group 203: 	202 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	204 
    -- CP-element group 203:  members (3) 
      -- CP-element group 203: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1043_sample_start_
      -- CP-element group 203: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1043_Sample/$entry
      -- CP-element group 203: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1043_Sample/req
      -- 
    req_2254_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2254_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(203), ack => WPIPE_Concat_output_pipe_1043_inst_req_0); -- 
    concat_cp_element_group_203: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_203"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_664_elements(193) & concat_CP_664_elements(202);
      gj_concat_cp_element_group_203 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_664_elements(203), clk => clk, reset => reset); --
    end block;
    -- CP-element group 204:  transition  input  output  bypass 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	203 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	205 
    -- CP-element group 204:  members (6) 
      -- CP-element group 204: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1043_sample_completed_
      -- CP-element group 204: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1043_update_start_
      -- CP-element group 204: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1043_Sample/$exit
      -- CP-element group 204: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1043_Update/req
      -- CP-element group 204: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1043_Update/$entry
      -- CP-element group 204: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1043_Sample/ack
      -- 
    ack_2255_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 204_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1043_inst_ack_0, ack => concat_CP_664_elements(204)); -- 
    req_2259_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2259_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(204), ack => WPIPE_Concat_output_pipe_1043_inst_req_1); -- 
    -- CP-element group 205:  transition  input  bypass 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	204 
    -- CP-element group 205: successors 
    -- CP-element group 205: 	206 
    -- CP-element group 205:  members (3) 
      -- CP-element group 205: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1043_update_completed_
      -- CP-element group 205: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1043_Update/ack
      -- CP-element group 205: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1043_Update/$exit
      -- 
    ack_2260_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1043_inst_ack_1, ack => concat_CP_664_elements(205)); -- 
    -- CP-element group 206:  join  transition  output  bypass 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	191 
    -- CP-element group 206: 	205 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	207 
    -- CP-element group 206:  members (3) 
      -- CP-element group 206: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1046_Sample/req
      -- CP-element group 206: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1046_Sample/$entry
      -- CP-element group 206: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1046_sample_start_
      -- 
    req_2268_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2268_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(206), ack => WPIPE_Concat_output_pipe_1046_inst_req_0); -- 
    concat_cp_element_group_206: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_206"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_664_elements(191) & concat_CP_664_elements(205);
      gj_concat_cp_element_group_206 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_664_elements(206), clk => clk, reset => reset); --
    end block;
    -- CP-element group 207:  transition  input  output  bypass 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	206 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	208 
    -- CP-element group 207:  members (6) 
      -- CP-element group 207: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1046_Update/req
      -- CP-element group 207: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1046_Update/$entry
      -- CP-element group 207: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1046_Sample/ack
      -- CP-element group 207: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1046_Sample/$exit
      -- CP-element group 207: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1046_update_start_
      -- CP-element group 207: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1046_sample_completed_
      -- 
    ack_2269_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 207_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1046_inst_ack_0, ack => concat_CP_664_elements(207)); -- 
    req_2273_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2273_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(207), ack => WPIPE_Concat_output_pipe_1046_inst_req_1); -- 
    -- CP-element group 208:  transition  input  bypass 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	207 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	209 
    -- CP-element group 208:  members (3) 
      -- CP-element group 208: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1046_Update/ack
      -- CP-element group 208: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1046_Update/$exit
      -- CP-element group 208: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1046_update_completed_
      -- 
    ack_2274_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 208_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1046_inst_ack_1, ack => concat_CP_664_elements(208)); -- 
    -- CP-element group 209:  join  transition  output  bypass 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	189 
    -- CP-element group 209: 	208 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	210 
    -- CP-element group 209:  members (3) 
      -- CP-element group 209: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1049_Sample/req
      -- CP-element group 209: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1049_Sample/$entry
      -- CP-element group 209: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1049_sample_start_
      -- 
    req_2282_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2282_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(209), ack => WPIPE_Concat_output_pipe_1049_inst_req_0); -- 
    concat_cp_element_group_209: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_209"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_664_elements(189) & concat_CP_664_elements(208);
      gj_concat_cp_element_group_209 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_664_elements(209), clk => clk, reset => reset); --
    end block;
    -- CP-element group 210:  transition  input  output  bypass 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	209 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	211 
    -- CP-element group 210:  members (6) 
      -- CP-element group 210: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1049_Update/$entry
      -- CP-element group 210: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1049_Update/req
      -- CP-element group 210: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1049_Sample/$exit
      -- CP-element group 210: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1049_Sample/ack
      -- CP-element group 210: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1049_update_start_
      -- CP-element group 210: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1049_sample_completed_
      -- 
    ack_2283_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 210_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1049_inst_ack_0, ack => concat_CP_664_elements(210)); -- 
    req_2287_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2287_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(210), ack => WPIPE_Concat_output_pipe_1049_inst_req_1); -- 
    -- CP-element group 211:  transition  input  bypass 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	210 
    -- CP-element group 211: successors 
    -- CP-element group 211: 	212 
    -- CP-element group 211:  members (3) 
      -- CP-element group 211: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1049_Update/$exit
      -- CP-element group 211: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1049_Update/ack
      -- CP-element group 211: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1049_update_completed_
      -- 
    ack_2288_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 211_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1049_inst_ack_1, ack => concat_CP_664_elements(211)); -- 
    -- CP-element group 212:  join  transition  output  bypass 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	187 
    -- CP-element group 212: 	211 
    -- CP-element group 212: successors 
    -- CP-element group 212: 	213 
    -- CP-element group 212:  members (3) 
      -- CP-element group 212: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1052_sample_start_
      -- CP-element group 212: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1052_Sample/$entry
      -- CP-element group 212: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1052_Sample/req
      -- 
    req_2296_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2296_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(212), ack => WPIPE_Concat_output_pipe_1052_inst_req_0); -- 
    concat_cp_element_group_212: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_212"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_664_elements(187) & concat_CP_664_elements(211);
      gj_concat_cp_element_group_212 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_664_elements(212), clk => clk, reset => reset); --
    end block;
    -- CP-element group 213:  transition  input  output  bypass 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	212 
    -- CP-element group 213: successors 
    -- CP-element group 213: 	214 
    -- CP-element group 213:  members (6) 
      -- CP-element group 213: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1052_sample_completed_
      -- CP-element group 213: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1052_update_start_
      -- CP-element group 213: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1052_Sample/$exit
      -- CP-element group 213: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1052_Sample/ack
      -- CP-element group 213: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1052_Update/$entry
      -- CP-element group 213: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1052_Update/req
      -- 
    ack_2297_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1052_inst_ack_0, ack => concat_CP_664_elements(213)); -- 
    req_2301_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2301_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(213), ack => WPIPE_Concat_output_pipe_1052_inst_req_1); -- 
    -- CP-element group 214:  transition  input  bypass 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	213 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	215 
    -- CP-element group 214:  members (3) 
      -- CP-element group 214: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1052_update_completed_
      -- CP-element group 214: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1052_Update/$exit
      -- CP-element group 214: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1052_Update/ack
      -- 
    ack_2302_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 214_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1052_inst_ack_1, ack => concat_CP_664_elements(214)); -- 
    -- CP-element group 215:  join  transition  output  bypass 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	185 
    -- CP-element group 215: 	214 
    -- CP-element group 215: successors 
    -- CP-element group 215: 	216 
    -- CP-element group 215:  members (3) 
      -- CP-element group 215: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1055_Sample/$entry
      -- CP-element group 215: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1055_Sample/req
      -- CP-element group 215: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1055_sample_start_
      -- 
    req_2310_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2310_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(215), ack => WPIPE_Concat_output_pipe_1055_inst_req_0); -- 
    concat_cp_element_group_215: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_215"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_664_elements(185) & concat_CP_664_elements(214);
      gj_concat_cp_element_group_215 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_664_elements(215), clk => clk, reset => reset); --
    end block;
    -- CP-element group 216:  transition  input  output  bypass 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	215 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	217 
    -- CP-element group 216:  members (6) 
      -- CP-element group 216: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1055_update_start_
      -- CP-element group 216: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1055_Sample/$exit
      -- CP-element group 216: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1055_Sample/ack
      -- CP-element group 216: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1055_Update/$entry
      -- CP-element group 216: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1055_sample_completed_
      -- CP-element group 216: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1055_Update/req
      -- 
    ack_2311_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1055_inst_ack_0, ack => concat_CP_664_elements(216)); -- 
    req_2315_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2315_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(216), ack => WPIPE_Concat_output_pipe_1055_inst_req_1); -- 
    -- CP-element group 217:  transition  input  bypass 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	216 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	218 
    -- CP-element group 217:  members (3) 
      -- CP-element group 217: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1055_update_completed_
      -- CP-element group 217: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1055_Update/$exit
      -- CP-element group 217: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1055_Update/ack
      -- 
    ack_2316_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 217_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1055_inst_ack_1, ack => concat_CP_664_elements(217)); -- 
    -- CP-element group 218:  join  transition  output  bypass 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	183 
    -- CP-element group 218: 	217 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	219 
    -- CP-element group 218:  members (3) 
      -- CP-element group 218: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1058_Sample/req
      -- CP-element group 218: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1058_Sample/$entry
      -- CP-element group 218: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1058_sample_start_
      -- 
    req_2324_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2324_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(218), ack => WPIPE_Concat_output_pipe_1058_inst_req_0); -- 
    concat_cp_element_group_218: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_218"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_664_elements(183) & concat_CP_664_elements(217);
      gj_concat_cp_element_group_218 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_664_elements(218), clk => clk, reset => reset); --
    end block;
    -- CP-element group 219:  transition  input  output  bypass 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	218 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	220 
    -- CP-element group 219:  members (6) 
      -- CP-element group 219: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1058_Update/req
      -- CP-element group 219: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1058_Update/$entry
      -- CP-element group 219: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1058_Sample/ack
      -- CP-element group 219: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1058_Sample/$exit
      -- CP-element group 219: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1058_update_start_
      -- CP-element group 219: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1058_sample_completed_
      -- 
    ack_2325_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 219_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1058_inst_ack_0, ack => concat_CP_664_elements(219)); -- 
    req_2329_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2329_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(219), ack => WPIPE_Concat_output_pipe_1058_inst_req_1); -- 
    -- CP-element group 220:  branch  transition  place  input  output  bypass 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	219 
    -- CP-element group 220: successors 
    -- CP-element group 220: 	221 
    -- CP-element group 220: 	222 
    -- CP-element group 220:  members (17) 
      -- CP-element group 220: 	 branch_block_stmt_216/assign_stmt_1067__entry__
      -- CP-element group 220: 	 branch_block_stmt_216/assign_stmt_1067__exit__
      -- CP-element group 220: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060__exit__
      -- CP-element group 220: 	 branch_block_stmt_216/if_stmt_1068__entry__
      -- CP-element group 220: 	 branch_block_stmt_216/R_cmp303381_1069_place
      -- CP-element group 220: 	 branch_block_stmt_216/if_stmt_1068_else_link/$entry
      -- CP-element group 220: 	 branch_block_stmt_216/if_stmt_1068_if_link/$entry
      -- CP-element group 220: 	 branch_block_stmt_216/if_stmt_1068_eval_test/branch_req
      -- CP-element group 220: 	 branch_block_stmt_216/if_stmt_1068_eval_test/$exit
      -- CP-element group 220: 	 branch_block_stmt_216/if_stmt_1068_eval_test/$entry
      -- CP-element group 220: 	 branch_block_stmt_216/if_stmt_1068_dead_link/$entry
      -- CP-element group 220: 	 branch_block_stmt_216/assign_stmt_1067/$exit
      -- CP-element group 220: 	 branch_block_stmt_216/assign_stmt_1067/$entry
      -- CP-element group 220: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1058_Update/ack
      -- CP-element group 220: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1058_Update/$exit
      -- CP-element group 220: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/WPIPE_Concat_output_pipe_1058_update_completed_
      -- CP-element group 220: 	 branch_block_stmt_216/call_stmt_952_to_assign_stmt_1060/$exit
      -- 
    ack_2330_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1058_inst_ack_1, ack => concat_CP_664_elements(220)); -- 
    branch_req_2341_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2341_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(220), ack => if_stmt_1068_branch_req_0); -- 
    -- CP-element group 221:  merge  transition  place  input  bypass 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	220 
    -- CP-element group 221: successors 
    -- CP-element group 221: 	285 
    -- CP-element group 221:  members (18) 
      -- CP-element group 221: 	 branch_block_stmt_216/assign_stmt_1079_to_assign_stmt_1103__entry__
      -- CP-element group 221: 	 branch_block_stmt_216/assign_stmt_1079_to_assign_stmt_1103__exit__
      -- CP-element group 221: 	 branch_block_stmt_216/merge_stmt_1074__exit__
      -- CP-element group 221: 	 branch_block_stmt_216/bbx_xnph_forx_xbody305
      -- CP-element group 221: 	 branch_block_stmt_216/forx_xend224_bbx_xnph
      -- CP-element group 221: 	 branch_block_stmt_216/assign_stmt_1079_to_assign_stmt_1103/$exit
      -- CP-element group 221: 	 branch_block_stmt_216/assign_stmt_1079_to_assign_stmt_1103/$entry
      -- CP-element group 221: 	 branch_block_stmt_216/if_stmt_1068_if_link/if_choice_transition
      -- CP-element group 221: 	 branch_block_stmt_216/if_stmt_1068_if_link/$exit
      -- CP-element group 221: 	 branch_block_stmt_216/forx_xend224_bbx_xnph_PhiReq/$entry
      -- CP-element group 221: 	 branch_block_stmt_216/forx_xend224_bbx_xnph_PhiReq/$exit
      -- CP-element group 221: 	 branch_block_stmt_216/merge_stmt_1074_PhiReqMerge
      -- CP-element group 221: 	 branch_block_stmt_216/merge_stmt_1074_PhiAck/$entry
      -- CP-element group 221: 	 branch_block_stmt_216/merge_stmt_1074_PhiAck/$exit
      -- CP-element group 221: 	 branch_block_stmt_216/merge_stmt_1074_PhiAck/dummy
      -- CP-element group 221: 	 branch_block_stmt_216/bbx_xnph_forx_xbody305_PhiReq/$entry
      -- CP-element group 221: 	 branch_block_stmt_216/bbx_xnph_forx_xbody305_PhiReq/phi_stmt_1106/$entry
      -- CP-element group 221: 	 branch_block_stmt_216/bbx_xnph_forx_xbody305_PhiReq/phi_stmt_1106/phi_stmt_1106_sources/$entry
      -- 
    if_choice_transition_2346_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1068_branch_ack_1, ack => concat_CP_664_elements(221)); -- 
    -- CP-element group 222:  transition  place  input  bypass 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	220 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	291 
    -- CP-element group 222:  members (5) 
      -- CP-element group 222: 	 branch_block_stmt_216/forx_xend224_forx_xend377
      -- CP-element group 222: 	 branch_block_stmt_216/if_stmt_1068_else_link/else_choice_transition
      -- CP-element group 222: 	 branch_block_stmt_216/if_stmt_1068_else_link/$exit
      -- CP-element group 222: 	 branch_block_stmt_216/forx_xend224_forx_xend377_PhiReq/$entry
      -- CP-element group 222: 	 branch_block_stmt_216/forx_xend224_forx_xend377_PhiReq/$exit
      -- 
    else_choice_transition_2350_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 222_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1068_branch_ack_0, ack => concat_CP_664_elements(222)); -- 
    -- CP-element group 223:  transition  input  bypass 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	290 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	268 
    -- CP-element group 223:  members (3) 
      -- CP-element group 223: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/array_obj_ref_1120_final_index_sum_regn_Sample/ack
      -- CP-element group 223: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/array_obj_ref_1120_final_index_sum_regn_Sample/$exit
      -- CP-element group 223: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/array_obj_ref_1120_final_index_sum_regn_sample_complete
      -- 
    ack_2384_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 223_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1120_index_offset_ack_0, ack => concat_CP_664_elements(223)); -- 
    -- CP-element group 224:  transition  input  output  bypass 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	290 
    -- CP-element group 224: successors 
    -- CP-element group 224: 	225 
    -- CP-element group 224:  members (11) 
      -- CP-element group 224: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/addr_of_1121_request/req
      -- CP-element group 224: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/array_obj_ref_1120_final_index_sum_regn_Update/$exit
      -- CP-element group 224: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/array_obj_ref_1120_final_index_sum_regn_Update/ack
      -- CP-element group 224: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/array_obj_ref_1120_base_plus_offset/sum_rename_ack
      -- CP-element group 224: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/array_obj_ref_1120_base_plus_offset/$exit
      -- CP-element group 224: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/addr_of_1121_request/$entry
      -- CP-element group 224: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/array_obj_ref_1120_base_plus_offset/$entry
      -- CP-element group 224: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/array_obj_ref_1120_base_plus_offset/sum_rename_req
      -- CP-element group 224: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/array_obj_ref_1120_offset_calculated
      -- CP-element group 224: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/array_obj_ref_1120_root_address_calculated
      -- CP-element group 224: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/addr_of_1121_sample_start_
      -- 
    ack_2389_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1120_index_offset_ack_1, ack => concat_CP_664_elements(224)); -- 
    req_2398_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2398_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(224), ack => addr_of_1121_final_reg_req_0); -- 
    -- CP-element group 225:  transition  input  bypass 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	224 
    -- CP-element group 225: successors 
    -- CP-element group 225:  members (3) 
      -- CP-element group 225: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/addr_of_1121_request/$exit
      -- CP-element group 225: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/addr_of_1121_request/ack
      -- CP-element group 225: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/addr_of_1121_sample_completed_
      -- 
    ack_2399_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 225_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1121_final_reg_ack_0, ack => concat_CP_664_elements(225)); -- 
    -- CP-element group 226:  join  fork  transition  input  output  bypass 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	290 
    -- CP-element group 226: successors 
    -- CP-element group 226: 	227 
    -- CP-element group 226:  members (24) 
      -- CP-element group 226: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/ptr_deref_1125_base_plus_offset/sum_rename_ack
      -- CP-element group 226: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/ptr_deref_1125_word_addrgen/$exit
      -- CP-element group 226: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/ptr_deref_1125_base_plus_offset/sum_rename_req
      -- CP-element group 226: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/ptr_deref_1125_word_addrgen/$entry
      -- CP-element group 226: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/ptr_deref_1125_Sample/word_access_start/$entry
      -- CP-element group 226: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/ptr_deref_1125_Sample/$entry
      -- CP-element group 226: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/ptr_deref_1125_word_addrgen/root_register_req
      -- CP-element group 226: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/ptr_deref_1125_word_addrgen/root_register_ack
      -- CP-element group 226: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/addr_of_1121_complete/$exit
      -- CP-element group 226: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/addr_of_1121_complete/ack
      -- CP-element group 226: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/ptr_deref_1125_sample_start_
      -- CP-element group 226: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/ptr_deref_1125_Sample/word_access_start/word_0/$entry
      -- CP-element group 226: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/ptr_deref_1125_base_address_calculated
      -- CP-element group 226: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/ptr_deref_1125_word_address_calculated
      -- CP-element group 226: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/ptr_deref_1125_root_address_calculated
      -- CP-element group 226: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/ptr_deref_1125_base_address_resized
      -- CP-element group 226: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/ptr_deref_1125_base_addr_resize/$entry
      -- CP-element group 226: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/ptr_deref_1125_base_addr_resize/$exit
      -- CP-element group 226: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/ptr_deref_1125_base_addr_resize/base_resize_req
      -- CP-element group 226: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/ptr_deref_1125_base_addr_resize/base_resize_ack
      -- CP-element group 226: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/ptr_deref_1125_Sample/word_access_start/word_0/rr
      -- CP-element group 226: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/ptr_deref_1125_base_plus_offset/$exit
      -- CP-element group 226: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/ptr_deref_1125_base_plus_offset/$entry
      -- CP-element group 226: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/addr_of_1121_update_completed_
      -- 
    ack_2404_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 226_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1121_final_reg_ack_1, ack => concat_CP_664_elements(226)); -- 
    rr_2437_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2437_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(226), ack => ptr_deref_1125_load_0_req_0); -- 
    -- CP-element group 227:  transition  input  bypass 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	226 
    -- CP-element group 227: successors 
    -- CP-element group 227:  members (5) 
      -- CP-element group 227: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/ptr_deref_1125_Sample/word_access_start/$exit
      -- CP-element group 227: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/ptr_deref_1125_Sample/$exit
      -- CP-element group 227: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/ptr_deref_1125_Sample/word_access_start/word_0/$exit
      -- CP-element group 227: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/ptr_deref_1125_sample_completed_
      -- CP-element group 227: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/ptr_deref_1125_Sample/word_access_start/word_0/ra
      -- 
    ra_2438_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 227_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1125_load_0_ack_0, ack => concat_CP_664_elements(227)); -- 
    -- CP-element group 228:  fork  transition  input  output  bypass 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	290 
    -- CP-element group 228: successors 
    -- CP-element group 228: 	229 
    -- CP-element group 228: 	231 
    -- CP-element group 228: 	233 
    -- CP-element group 228: 	235 
    -- CP-element group 228: 	237 
    -- CP-element group 228: 	239 
    -- CP-element group 228: 	241 
    -- CP-element group 228: 	243 
    -- CP-element group 228:  members (33) 
      -- CP-element group 228: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1179_Sample/rr
      -- CP-element group 228: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1139_Sample/rr
      -- CP-element group 228: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1169_Sample/rr
      -- CP-element group 228: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1199_Sample/rr
      -- CP-element group 228: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1149_sample_start_
      -- CP-element group 228: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1179_Sample/$entry
      -- CP-element group 228: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1179_sample_start_
      -- CP-element group 228: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1149_Sample/$entry
      -- CP-element group 228: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1149_Sample/rr
      -- CP-element group 228: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/ptr_deref_1125_update_completed_
      -- CP-element group 228: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1189_sample_start_
      -- CP-element group 228: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1159_sample_start_
      -- CP-element group 228: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1169_Sample/$entry
      -- CP-element group 228: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1139_Sample/$entry
      -- CP-element group 228: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1199_Sample/$entry
      -- CP-element group 228: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1139_sample_start_
      -- CP-element group 228: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1129_Sample/rr
      -- CP-element group 228: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1129_Sample/$entry
      -- CP-element group 228: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1169_sample_start_
      -- CP-element group 228: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1129_sample_start_
      -- CP-element group 228: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/ptr_deref_1125_Update/ptr_deref_1125_Merge/merge_ack
      -- CP-element group 228: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1199_sample_start_
      -- CP-element group 228: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/ptr_deref_1125_Update/ptr_deref_1125_Merge/merge_req
      -- CP-element group 228: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/ptr_deref_1125_Update/ptr_deref_1125_Merge/$exit
      -- CP-element group 228: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/ptr_deref_1125_Update/ptr_deref_1125_Merge/$entry
      -- CP-element group 228: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/ptr_deref_1125_Update/word_access_complete/word_0/ca
      -- CP-element group 228: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/ptr_deref_1125_Update/word_access_complete/word_0/$exit
      -- CP-element group 228: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1159_Sample/rr
      -- CP-element group 228: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1189_Sample/rr
      -- CP-element group 228: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/ptr_deref_1125_Update/word_access_complete/$exit
      -- CP-element group 228: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/ptr_deref_1125_Update/$exit
      -- CP-element group 228: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1159_Sample/$entry
      -- CP-element group 228: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1189_Sample/$entry
      -- 
    ca_2449_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 228_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1125_load_0_ack_1, ack => concat_CP_664_elements(228)); -- 
    rr_2462_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2462_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(228), ack => type_cast_1129_inst_req_0); -- 
    rr_2476_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2476_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(228), ack => type_cast_1139_inst_req_0); -- 
    rr_2490_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2490_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(228), ack => type_cast_1149_inst_req_0); -- 
    rr_2504_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2504_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(228), ack => type_cast_1159_inst_req_0); -- 
    rr_2518_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2518_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(228), ack => type_cast_1169_inst_req_0); -- 
    rr_2532_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2532_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(228), ack => type_cast_1179_inst_req_0); -- 
    rr_2546_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2546_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(228), ack => type_cast_1189_inst_req_0); -- 
    rr_2560_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2560_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(228), ack => type_cast_1199_inst_req_0); -- 
    -- CP-element group 229:  transition  input  bypass 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	228 
    -- CP-element group 229: successors 
    -- CP-element group 229:  members (3) 
      -- CP-element group 229: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1129_Sample/ra
      -- CP-element group 229: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1129_Sample/$exit
      -- CP-element group 229: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1129_sample_completed_
      -- 
    ra_2463_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 229_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1129_inst_ack_0, ack => concat_CP_664_elements(229)); -- 
    -- CP-element group 230:  transition  input  bypass 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	290 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	265 
    -- CP-element group 230:  members (3) 
      -- CP-element group 230: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1129_Update/ca
      -- CP-element group 230: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1129_Update/$exit
      -- CP-element group 230: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1129_update_completed_
      -- 
    ca_2468_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 230_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1129_inst_ack_1, ack => concat_CP_664_elements(230)); -- 
    -- CP-element group 231:  transition  input  bypass 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	228 
    -- CP-element group 231: successors 
    -- CP-element group 231:  members (3) 
      -- CP-element group 231: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1139_Sample/$exit
      -- CP-element group 231: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1139_Sample/ra
      -- CP-element group 231: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1139_sample_completed_
      -- 
    ra_2477_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 231_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1139_inst_ack_0, ack => concat_CP_664_elements(231)); -- 
    -- CP-element group 232:  transition  input  bypass 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	290 
    -- CP-element group 232: successors 
    -- CP-element group 232: 	262 
    -- CP-element group 232:  members (3) 
      -- CP-element group 232: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1139_Update/ca
      -- CP-element group 232: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1139_Update/$exit
      -- CP-element group 232: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1139_update_completed_
      -- 
    ca_2482_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 232_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1139_inst_ack_1, ack => concat_CP_664_elements(232)); -- 
    -- CP-element group 233:  transition  input  bypass 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	228 
    -- CP-element group 233: successors 
    -- CP-element group 233:  members (3) 
      -- CP-element group 233: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1149_sample_completed_
      -- CP-element group 233: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1149_Sample/$exit
      -- CP-element group 233: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1149_Sample/ra
      -- 
    ra_2491_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 233_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1149_inst_ack_0, ack => concat_CP_664_elements(233)); -- 
    -- CP-element group 234:  transition  input  bypass 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	290 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	259 
    -- CP-element group 234:  members (3) 
      -- CP-element group 234: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1149_update_completed_
      -- CP-element group 234: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1149_Update/$exit
      -- CP-element group 234: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1149_Update/ca
      -- 
    ca_2496_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 234_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1149_inst_ack_1, ack => concat_CP_664_elements(234)); -- 
    -- CP-element group 235:  transition  input  bypass 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	228 
    -- CP-element group 235: successors 
    -- CP-element group 235:  members (3) 
      -- CP-element group 235: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1159_sample_completed_
      -- CP-element group 235: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1159_Sample/ra
      -- CP-element group 235: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1159_Sample/$exit
      -- 
    ra_2505_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 235_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1159_inst_ack_0, ack => concat_CP_664_elements(235)); -- 
    -- CP-element group 236:  transition  input  bypass 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	290 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	256 
    -- CP-element group 236:  members (3) 
      -- CP-element group 236: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1159_update_completed_
      -- CP-element group 236: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1159_Update/ca
      -- CP-element group 236: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1159_Update/$exit
      -- 
    ca_2510_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 236_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1159_inst_ack_1, ack => concat_CP_664_elements(236)); -- 
    -- CP-element group 237:  transition  input  bypass 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	228 
    -- CP-element group 237: successors 
    -- CP-element group 237:  members (3) 
      -- CP-element group 237: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1169_Sample/$exit
      -- CP-element group 237: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1169_Sample/ra
      -- CP-element group 237: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1169_sample_completed_
      -- 
    ra_2519_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 237_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1169_inst_ack_0, ack => concat_CP_664_elements(237)); -- 
    -- CP-element group 238:  transition  input  bypass 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	290 
    -- CP-element group 238: successors 
    -- CP-element group 238: 	253 
    -- CP-element group 238:  members (3) 
      -- CP-element group 238: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1169_Update/ca
      -- CP-element group 238: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1169_Update/$exit
      -- CP-element group 238: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1169_update_completed_
      -- 
    ca_2524_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 238_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1169_inst_ack_1, ack => concat_CP_664_elements(238)); -- 
    -- CP-element group 239:  transition  input  bypass 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	228 
    -- CP-element group 239: successors 
    -- CP-element group 239:  members (3) 
      -- CP-element group 239: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1179_Sample/$exit
      -- CP-element group 239: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1179_sample_completed_
      -- CP-element group 239: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1179_Sample/ra
      -- 
    ra_2533_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 239_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1179_inst_ack_0, ack => concat_CP_664_elements(239)); -- 
    -- CP-element group 240:  transition  input  bypass 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	290 
    -- CP-element group 240: successors 
    -- CP-element group 240: 	250 
    -- CP-element group 240:  members (3) 
      -- CP-element group 240: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1179_update_completed_
      -- CP-element group 240: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1179_Update/$exit
      -- CP-element group 240: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1179_Update/ca
      -- 
    ca_2538_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 240_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1179_inst_ack_1, ack => concat_CP_664_elements(240)); -- 
    -- CP-element group 241:  transition  input  bypass 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	228 
    -- CP-element group 241: successors 
    -- CP-element group 241:  members (3) 
      -- CP-element group 241: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1189_sample_completed_
      -- CP-element group 241: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1189_Sample/ra
      -- CP-element group 241: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1189_Sample/$exit
      -- 
    ra_2547_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 241_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1189_inst_ack_0, ack => concat_CP_664_elements(241)); -- 
    -- CP-element group 242:  transition  input  bypass 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	290 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	247 
    -- CP-element group 242:  members (3) 
      -- CP-element group 242: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1189_Update/ca
      -- CP-element group 242: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1189_Update/$exit
      -- CP-element group 242: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1189_update_completed_
      -- 
    ca_2552_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 242_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1189_inst_ack_1, ack => concat_CP_664_elements(242)); -- 
    -- CP-element group 243:  transition  input  bypass 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	228 
    -- CP-element group 243: successors 
    -- CP-element group 243:  members (3) 
      -- CP-element group 243: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1199_Sample/ra
      -- CP-element group 243: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1199_Sample/$exit
      -- CP-element group 243: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1199_sample_completed_
      -- 
    ra_2561_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 243_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1199_inst_ack_0, ack => concat_CP_664_elements(243)); -- 
    -- CP-element group 244:  transition  input  output  bypass 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	290 
    -- CP-element group 244: successors 
    -- CP-element group 244: 	245 
    -- CP-element group 244:  members (6) 
      -- CP-element group 244: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1199_Update/$exit
      -- CP-element group 244: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1199_Update/ca
      -- CP-element group 244: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1201_sample_start_
      -- CP-element group 244: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1201_Sample/req
      -- CP-element group 244: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1199_update_completed_
      -- CP-element group 244: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1201_Sample/$entry
      -- 
    ca_2566_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 244_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1199_inst_ack_1, ack => concat_CP_664_elements(244)); -- 
    req_2574_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2574_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(244), ack => WPIPE_Concat_output_pipe_1201_inst_req_0); -- 
    -- CP-element group 245:  transition  input  output  bypass 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	244 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	246 
    -- CP-element group 245:  members (6) 
      -- CP-element group 245: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1201_Update/req
      -- CP-element group 245: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1201_Update/$entry
      -- CP-element group 245: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1201_Sample/ack
      -- CP-element group 245: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1201_Sample/$exit
      -- CP-element group 245: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1201_update_start_
      -- CP-element group 245: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1201_sample_completed_
      -- 
    ack_2575_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 245_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1201_inst_ack_0, ack => concat_CP_664_elements(245)); -- 
    req_2579_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2579_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(245), ack => WPIPE_Concat_output_pipe_1201_inst_req_1); -- 
    -- CP-element group 246:  transition  input  bypass 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	245 
    -- CP-element group 246: successors 
    -- CP-element group 246: 	247 
    -- CP-element group 246:  members (3) 
      -- CP-element group 246: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1201_Update/ack
      -- CP-element group 246: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1201_Update/$exit
      -- CP-element group 246: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1201_update_completed_
      -- 
    ack_2580_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 246_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1201_inst_ack_1, ack => concat_CP_664_elements(246)); -- 
    -- CP-element group 247:  join  transition  output  bypass 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	242 
    -- CP-element group 247: 	246 
    -- CP-element group 247: successors 
    -- CP-element group 247: 	248 
    -- CP-element group 247:  members (3) 
      -- CP-element group 247: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1204_Sample/req
      -- CP-element group 247: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1204_Sample/$entry
      -- CP-element group 247: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1204_sample_start_
      -- 
    req_2588_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2588_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(247), ack => WPIPE_Concat_output_pipe_1204_inst_req_0); -- 
    concat_cp_element_group_247: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_247"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_664_elements(242) & concat_CP_664_elements(246);
      gj_concat_cp_element_group_247 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_664_elements(247), clk => clk, reset => reset); --
    end block;
    -- CP-element group 248:  transition  input  output  bypass 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	247 
    -- CP-element group 248: successors 
    -- CP-element group 248: 	249 
    -- CP-element group 248:  members (6) 
      -- CP-element group 248: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1204_Update/$entry
      -- CP-element group 248: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1204_Update/req
      -- CP-element group 248: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1204_Sample/ack
      -- CP-element group 248: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1204_Sample/$exit
      -- CP-element group 248: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1204_update_start_
      -- CP-element group 248: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1204_sample_completed_
      -- 
    ack_2589_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 248_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1204_inst_ack_0, ack => concat_CP_664_elements(248)); -- 
    req_2593_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2593_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(248), ack => WPIPE_Concat_output_pipe_1204_inst_req_1); -- 
    -- CP-element group 249:  transition  input  bypass 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	248 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	250 
    -- CP-element group 249:  members (3) 
      -- CP-element group 249: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1204_Update/$exit
      -- CP-element group 249: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1204_Update/ack
      -- CP-element group 249: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1204_update_completed_
      -- 
    ack_2594_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 249_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1204_inst_ack_1, ack => concat_CP_664_elements(249)); -- 
    -- CP-element group 250:  join  transition  output  bypass 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	249 
    -- CP-element group 250: 	240 
    -- CP-element group 250: successors 
    -- CP-element group 250: 	251 
    -- CP-element group 250:  members (3) 
      -- CP-element group 250: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1207_sample_start_
      -- CP-element group 250: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1207_Sample/$entry
      -- CP-element group 250: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1207_Sample/req
      -- 
    req_2602_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2602_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(250), ack => WPIPE_Concat_output_pipe_1207_inst_req_0); -- 
    concat_cp_element_group_250: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_250"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_664_elements(249) & concat_CP_664_elements(240);
      gj_concat_cp_element_group_250 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_664_elements(250), clk => clk, reset => reset); --
    end block;
    -- CP-element group 251:  transition  input  output  bypass 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	250 
    -- CP-element group 251: successors 
    -- CP-element group 251: 	252 
    -- CP-element group 251:  members (6) 
      -- CP-element group 251: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1207_Sample/$exit
      -- CP-element group 251: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1207_Sample/ack
      -- CP-element group 251: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1207_update_start_
      -- CP-element group 251: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1207_Update/req
      -- CP-element group 251: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1207_sample_completed_
      -- CP-element group 251: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1207_Update/$entry
      -- 
    ack_2603_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 251_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1207_inst_ack_0, ack => concat_CP_664_elements(251)); -- 
    req_2607_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2607_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(251), ack => WPIPE_Concat_output_pipe_1207_inst_req_1); -- 
    -- CP-element group 252:  transition  input  bypass 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	251 
    -- CP-element group 252: successors 
    -- CP-element group 252: 	253 
    -- CP-element group 252:  members (3) 
      -- CP-element group 252: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1207_update_completed_
      -- CP-element group 252: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1207_Update/$exit
      -- CP-element group 252: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1207_Update/ack
      -- 
    ack_2608_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 252_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1207_inst_ack_1, ack => concat_CP_664_elements(252)); -- 
    -- CP-element group 253:  join  transition  output  bypass 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	252 
    -- CP-element group 253: 	238 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	254 
    -- CP-element group 253:  members (3) 
      -- CP-element group 253: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1210_sample_start_
      -- CP-element group 253: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1210_Sample/$entry
      -- CP-element group 253: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1210_Sample/req
      -- 
    req_2616_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2616_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(253), ack => WPIPE_Concat_output_pipe_1210_inst_req_0); -- 
    concat_cp_element_group_253: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_253"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_664_elements(252) & concat_CP_664_elements(238);
      gj_concat_cp_element_group_253 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_664_elements(253), clk => clk, reset => reset); --
    end block;
    -- CP-element group 254:  transition  input  output  bypass 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	253 
    -- CP-element group 254: successors 
    -- CP-element group 254: 	255 
    -- CP-element group 254:  members (6) 
      -- CP-element group 254: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1210_update_start_
      -- CP-element group 254: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1210_sample_completed_
      -- CP-element group 254: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1210_Sample/$exit
      -- CP-element group 254: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1210_Sample/ack
      -- CP-element group 254: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1210_Update/$entry
      -- CP-element group 254: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1210_Update/req
      -- 
    ack_2617_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 254_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1210_inst_ack_0, ack => concat_CP_664_elements(254)); -- 
    req_2621_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2621_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(254), ack => WPIPE_Concat_output_pipe_1210_inst_req_1); -- 
    -- CP-element group 255:  transition  input  bypass 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	254 
    -- CP-element group 255: successors 
    -- CP-element group 255: 	256 
    -- CP-element group 255:  members (3) 
      -- CP-element group 255: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1210_update_completed_
      -- CP-element group 255: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1210_Update/$exit
      -- CP-element group 255: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1210_Update/ack
      -- 
    ack_2622_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 255_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1210_inst_ack_1, ack => concat_CP_664_elements(255)); -- 
    -- CP-element group 256:  join  transition  output  bypass 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	255 
    -- CP-element group 256: 	236 
    -- CP-element group 256: successors 
    -- CP-element group 256: 	257 
    -- CP-element group 256:  members (3) 
      -- CP-element group 256: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1213_sample_start_
      -- CP-element group 256: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1213_Sample/$entry
      -- CP-element group 256: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1213_Sample/req
      -- 
    req_2630_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2630_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(256), ack => WPIPE_Concat_output_pipe_1213_inst_req_0); -- 
    concat_cp_element_group_256: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_256"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_664_elements(255) & concat_CP_664_elements(236);
      gj_concat_cp_element_group_256 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_664_elements(256), clk => clk, reset => reset); --
    end block;
    -- CP-element group 257:  transition  input  output  bypass 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	256 
    -- CP-element group 257: successors 
    -- CP-element group 257: 	258 
    -- CP-element group 257:  members (6) 
      -- CP-element group 257: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1213_sample_completed_
      -- CP-element group 257: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1213_update_start_
      -- CP-element group 257: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1213_Sample/$exit
      -- CP-element group 257: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1213_Sample/ack
      -- CP-element group 257: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1213_Update/$entry
      -- CP-element group 257: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1213_Update/req
      -- 
    ack_2631_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 257_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1213_inst_ack_0, ack => concat_CP_664_elements(257)); -- 
    req_2635_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2635_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(257), ack => WPIPE_Concat_output_pipe_1213_inst_req_1); -- 
    -- CP-element group 258:  transition  input  bypass 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	257 
    -- CP-element group 258: successors 
    -- CP-element group 258: 	259 
    -- CP-element group 258:  members (3) 
      -- CP-element group 258: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1213_update_completed_
      -- CP-element group 258: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1213_Update/$exit
      -- CP-element group 258: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1213_Update/ack
      -- 
    ack_2636_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 258_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1213_inst_ack_1, ack => concat_CP_664_elements(258)); -- 
    -- CP-element group 259:  join  transition  output  bypass 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	258 
    -- CP-element group 259: 	234 
    -- CP-element group 259: successors 
    -- CP-element group 259: 	260 
    -- CP-element group 259:  members (3) 
      -- CP-element group 259: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1216_sample_start_
      -- CP-element group 259: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1216_Sample/$entry
      -- CP-element group 259: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1216_Sample/req
      -- 
    req_2644_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2644_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(259), ack => WPIPE_Concat_output_pipe_1216_inst_req_0); -- 
    concat_cp_element_group_259: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_259"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_664_elements(258) & concat_CP_664_elements(234);
      gj_concat_cp_element_group_259 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_664_elements(259), clk => clk, reset => reset); --
    end block;
    -- CP-element group 260:  transition  input  output  bypass 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	259 
    -- CP-element group 260: successors 
    -- CP-element group 260: 	261 
    -- CP-element group 260:  members (6) 
      -- CP-element group 260: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1216_sample_completed_
      -- CP-element group 260: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1216_update_start_
      -- CP-element group 260: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1216_Sample/$exit
      -- CP-element group 260: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1216_Sample/ack
      -- CP-element group 260: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1216_Update/$entry
      -- CP-element group 260: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1216_Update/req
      -- 
    ack_2645_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 260_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1216_inst_ack_0, ack => concat_CP_664_elements(260)); -- 
    req_2649_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2649_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(260), ack => WPIPE_Concat_output_pipe_1216_inst_req_1); -- 
    -- CP-element group 261:  transition  input  bypass 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	260 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	262 
    -- CP-element group 261:  members (3) 
      -- CP-element group 261: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1216_update_completed_
      -- CP-element group 261: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1216_Update/$exit
      -- CP-element group 261: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1216_Update/ack
      -- 
    ack_2650_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 261_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1216_inst_ack_1, ack => concat_CP_664_elements(261)); -- 
    -- CP-element group 262:  join  transition  output  bypass 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	261 
    -- CP-element group 262: 	232 
    -- CP-element group 262: successors 
    -- CP-element group 262: 	263 
    -- CP-element group 262:  members (3) 
      -- CP-element group 262: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1219_sample_start_
      -- CP-element group 262: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1219_Sample/$entry
      -- CP-element group 262: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1219_Sample/req
      -- 
    req_2658_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2658_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(262), ack => WPIPE_Concat_output_pipe_1219_inst_req_0); -- 
    concat_cp_element_group_262: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_262"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_664_elements(261) & concat_CP_664_elements(232);
      gj_concat_cp_element_group_262 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_664_elements(262), clk => clk, reset => reset); --
    end block;
    -- CP-element group 263:  transition  input  output  bypass 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	262 
    -- CP-element group 263: successors 
    -- CP-element group 263: 	264 
    -- CP-element group 263:  members (6) 
      -- CP-element group 263: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1219_sample_completed_
      -- CP-element group 263: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1219_update_start_
      -- CP-element group 263: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1219_Sample/$exit
      -- CP-element group 263: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1219_Sample/ack
      -- CP-element group 263: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1219_Update/$entry
      -- CP-element group 263: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1219_Update/req
      -- 
    ack_2659_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 263_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1219_inst_ack_0, ack => concat_CP_664_elements(263)); -- 
    req_2663_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2663_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(263), ack => WPIPE_Concat_output_pipe_1219_inst_req_1); -- 
    -- CP-element group 264:  transition  input  bypass 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	263 
    -- CP-element group 264: successors 
    -- CP-element group 264: 	265 
    -- CP-element group 264:  members (3) 
      -- CP-element group 264: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1219_update_completed_
      -- CP-element group 264: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1219_Update/$exit
      -- CP-element group 264: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1219_Update/ack
      -- 
    ack_2664_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 264_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1219_inst_ack_1, ack => concat_CP_664_elements(264)); -- 
    -- CP-element group 265:  join  transition  output  bypass 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	264 
    -- CP-element group 265: 	230 
    -- CP-element group 265: successors 
    -- CP-element group 265: 	266 
    -- CP-element group 265:  members (3) 
      -- CP-element group 265: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1222_sample_start_
      -- CP-element group 265: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1222_Sample/$entry
      -- CP-element group 265: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1222_Sample/req
      -- 
    req_2672_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2672_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(265), ack => WPIPE_Concat_output_pipe_1222_inst_req_0); -- 
    concat_cp_element_group_265: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_265"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_664_elements(264) & concat_CP_664_elements(230);
      gj_concat_cp_element_group_265 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_664_elements(265), clk => clk, reset => reset); --
    end block;
    -- CP-element group 266:  transition  input  output  bypass 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	265 
    -- CP-element group 266: successors 
    -- CP-element group 266: 	267 
    -- CP-element group 266:  members (6) 
      -- CP-element group 266: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1222_sample_completed_
      -- CP-element group 266: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1222_update_start_
      -- CP-element group 266: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1222_Sample/$exit
      -- CP-element group 266: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1222_Sample/ack
      -- CP-element group 266: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1222_Update/$entry
      -- CP-element group 266: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1222_Update/req
      -- 
    ack_2673_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 266_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1222_inst_ack_0, ack => concat_CP_664_elements(266)); -- 
    req_2677_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2677_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(266), ack => WPIPE_Concat_output_pipe_1222_inst_req_1); -- 
    -- CP-element group 267:  transition  input  bypass 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	266 
    -- CP-element group 267: successors 
    -- CP-element group 267: 	268 
    -- CP-element group 267:  members (3) 
      -- CP-element group 267: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1222_update_completed_
      -- CP-element group 267: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1222_Update/$exit
      -- CP-element group 267: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/WPIPE_Concat_output_pipe_1222_Update/ack
      -- 
    ack_2678_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 267_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Concat_output_pipe_1222_inst_ack_1, ack => concat_CP_664_elements(267)); -- 
    -- CP-element group 268:  branch  join  transition  place  output  bypass 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	267 
    -- CP-element group 268: 	223 
    -- CP-element group 268: successors 
    -- CP-element group 268: 	269 
    -- CP-element group 268: 	270 
    -- CP-element group 268:  members (10) 
      -- CP-element group 268: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235__exit__
      -- CP-element group 268: 	 branch_block_stmt_216/if_stmt_1236__entry__
      -- CP-element group 268: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/$exit
      -- CP-element group 268: 	 branch_block_stmt_216/if_stmt_1236_dead_link/$entry
      -- CP-element group 268: 	 branch_block_stmt_216/if_stmt_1236_eval_test/$entry
      -- CP-element group 268: 	 branch_block_stmt_216/if_stmt_1236_eval_test/$exit
      -- CP-element group 268: 	 branch_block_stmt_216/if_stmt_1236_eval_test/branch_req
      -- CP-element group 268: 	 branch_block_stmt_216/R_exitcond5_1237_place
      -- CP-element group 268: 	 branch_block_stmt_216/if_stmt_1236_if_link/$entry
      -- CP-element group 268: 	 branch_block_stmt_216/if_stmt_1236_else_link/$entry
      -- 
    branch_req_2686_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2686_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(268), ack => if_stmt_1236_branch_req_0); -- 
    concat_cp_element_group_268: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_268"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_664_elements(267) & concat_CP_664_elements(223);
      gj_concat_cp_element_group_268 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_664_elements(268), clk => clk, reset => reset); --
    end block;
    -- CP-element group 269:  merge  transition  place  input  bypass 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: 	268 
    -- CP-element group 269: successors 
    -- CP-element group 269: 	291 
    -- CP-element group 269:  members (13) 
      -- CP-element group 269: 	 branch_block_stmt_216/merge_stmt_1242__exit__
      -- CP-element group 269: 	 branch_block_stmt_216/forx_xend377x_xloopexit_forx_xend377
      -- CP-element group 269: 	 branch_block_stmt_216/if_stmt_1236_if_link/$exit
      -- CP-element group 269: 	 branch_block_stmt_216/if_stmt_1236_if_link/if_choice_transition
      -- CP-element group 269: 	 branch_block_stmt_216/forx_xbody305_forx_xend377x_xloopexit
      -- CP-element group 269: 	 branch_block_stmt_216/forx_xbody305_forx_xend377x_xloopexit_PhiReq/$entry
      -- CP-element group 269: 	 branch_block_stmt_216/forx_xbody305_forx_xend377x_xloopexit_PhiReq/$exit
      -- CP-element group 269: 	 branch_block_stmt_216/merge_stmt_1242_PhiReqMerge
      -- CP-element group 269: 	 branch_block_stmt_216/merge_stmt_1242_PhiAck/$entry
      -- CP-element group 269: 	 branch_block_stmt_216/merge_stmt_1242_PhiAck/$exit
      -- CP-element group 269: 	 branch_block_stmt_216/merge_stmt_1242_PhiAck/dummy
      -- CP-element group 269: 	 branch_block_stmt_216/forx_xend377x_xloopexit_forx_xend377_PhiReq/$entry
      -- CP-element group 269: 	 branch_block_stmt_216/forx_xend377x_xloopexit_forx_xend377_PhiReq/$exit
      -- 
    if_choice_transition_2691_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 269_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1236_branch_ack_1, ack => concat_CP_664_elements(269)); -- 
    -- CP-element group 270:  fork  transition  place  input  output  bypass 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	268 
    -- CP-element group 270: successors 
    -- CP-element group 270: 	286 
    -- CP-element group 270: 	287 
    -- CP-element group 270:  members (12) 
      -- CP-element group 270: 	 branch_block_stmt_216/if_stmt_1236_else_link/$exit
      -- CP-element group 270: 	 branch_block_stmt_216/if_stmt_1236_else_link/else_choice_transition
      -- CP-element group 270: 	 branch_block_stmt_216/forx_xbody305_forx_xbody305
      -- CP-element group 270: 	 branch_block_stmt_216/forx_xbody305_forx_xbody305_PhiReq/$entry
      -- CP-element group 270: 	 branch_block_stmt_216/forx_xbody305_forx_xbody305_PhiReq/phi_stmt_1106/$entry
      -- CP-element group 270: 	 branch_block_stmt_216/forx_xbody305_forx_xbody305_PhiReq/phi_stmt_1106/phi_stmt_1106_sources/$entry
      -- CP-element group 270: 	 branch_block_stmt_216/forx_xbody305_forx_xbody305_PhiReq/phi_stmt_1106/phi_stmt_1106_sources/type_cast_1112/$entry
      -- CP-element group 270: 	 branch_block_stmt_216/forx_xbody305_forx_xbody305_PhiReq/phi_stmt_1106/phi_stmt_1106_sources/type_cast_1112/SplitProtocol/$entry
      -- CP-element group 270: 	 branch_block_stmt_216/forx_xbody305_forx_xbody305_PhiReq/phi_stmt_1106/phi_stmt_1106_sources/type_cast_1112/SplitProtocol/Sample/$entry
      -- CP-element group 270: 	 branch_block_stmt_216/forx_xbody305_forx_xbody305_PhiReq/phi_stmt_1106/phi_stmt_1106_sources/type_cast_1112/SplitProtocol/Sample/rr
      -- CP-element group 270: 	 branch_block_stmt_216/forx_xbody305_forx_xbody305_PhiReq/phi_stmt_1106/phi_stmt_1106_sources/type_cast_1112/SplitProtocol/Update/$entry
      -- CP-element group 270: 	 branch_block_stmt_216/forx_xbody305_forx_xbody305_PhiReq/phi_stmt_1106/phi_stmt_1106_sources/type_cast_1112/SplitProtocol/Update/cr
      -- 
    else_choice_transition_2695_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 270_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1236_branch_ack_0, ack => concat_CP_664_elements(270)); -- 
    rr_2893_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2893_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(270), ack => type_cast_1112_inst_req_0); -- 
    cr_2898_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2898_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(270), ack => type_cast_1112_inst_req_1); -- 
    -- CP-element group 271:  merge  branch  transition  place  output  bypass 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	81 
    -- CP-element group 271: 	126 
    -- CP-element group 271: successors 
    -- CP-element group 271: 	82 
    -- CP-element group 271: 	83 
    -- CP-element group 271:  members (17) 
      -- CP-element group 271: 	 branch_block_stmt_216/assign_stmt_512/$entry
      -- CP-element group 271: 	 branch_block_stmt_216/R_cmp169384_514_place
      -- CP-element group 271: 	 branch_block_stmt_216/if_stmt_513_eval_test/$exit
      -- CP-element group 271: 	 branch_block_stmt_216/assign_stmt_512/$exit
      -- CP-element group 271: 	 branch_block_stmt_216/assign_stmt_512__entry__
      -- CP-element group 271: 	 branch_block_stmt_216/if_stmt_513_else_link/$entry
      -- CP-element group 271: 	 branch_block_stmt_216/if_stmt_513_dead_link/$entry
      -- CP-element group 271: 	 branch_block_stmt_216/if_stmt_513_if_link/$entry
      -- CP-element group 271: 	 branch_block_stmt_216/if_stmt_513_eval_test/$entry
      -- CP-element group 271: 	 branch_block_stmt_216/merge_stmt_506__exit__
      -- CP-element group 271: 	 branch_block_stmt_216/if_stmt_513_eval_test/branch_req
      -- CP-element group 271: 	 branch_block_stmt_216/if_stmt_513__entry__
      -- CP-element group 271: 	 branch_block_stmt_216/assign_stmt_512__exit__
      -- CP-element group 271: 	 branch_block_stmt_216/merge_stmt_506_PhiReqMerge
      -- CP-element group 271: 	 branch_block_stmt_216/merge_stmt_506_PhiAck/$entry
      -- CP-element group 271: 	 branch_block_stmt_216/merge_stmt_506_PhiAck/$exit
      -- CP-element group 271: 	 branch_block_stmt_216/merge_stmt_506_PhiAck/dummy
      -- 
    branch_req_1298_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1298_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(271), ack => if_stmt_513_branch_req_0); -- 
    concat_CP_664_elements(271) <= OrReduce(concat_CP_664_elements(81) & concat_CP_664_elements(126));
    -- CP-element group 272:  transition  output  delay-element  bypass 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	85 
    -- CP-element group 272: successors 
    -- CP-element group 272: 	276 
    -- CP-element group 272:  members (5) 
      -- CP-element group 272: 	 branch_block_stmt_216/bbx_xnph390_forx_xbody_PhiReq/$exit
      -- CP-element group 272: 	 branch_block_stmt_216/bbx_xnph390_forx_xbody_PhiReq/phi_stmt_555/$exit
      -- CP-element group 272: 	 branch_block_stmt_216/bbx_xnph390_forx_xbody_PhiReq/phi_stmt_555/phi_stmt_555_sources/$exit
      -- CP-element group 272: 	 branch_block_stmt_216/bbx_xnph390_forx_xbody_PhiReq/phi_stmt_555/phi_stmt_555_sources/type_cast_559_konst_delay_trans
      -- CP-element group 272: 	 branch_block_stmt_216/bbx_xnph390_forx_xbody_PhiReq/phi_stmt_555/phi_stmt_555_req
      -- 
    phi_stmt_555_req_2743_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_555_req_2743_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(272), ack => phi_stmt_555_req_0); -- 
    -- Element group concat_CP_664_elements(272) is a control-delay.
    cp_element_272_delay: control_delay_element  generic map(name => " 272_delay", delay_value => 1)  port map(req => concat_CP_664_elements(85), ack => concat_CP_664_elements(272), clk => clk, reset =>reset);
    -- CP-element group 273:  transition  input  bypass 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: 	127 
    -- CP-element group 273: successors 
    -- CP-element group 273: 	275 
    -- CP-element group 273:  members (2) 
      -- CP-element group 273: 	 branch_block_stmt_216/forx_xbody_forx_xbody_PhiReq/phi_stmt_555/phi_stmt_555_sources/type_cast_561/SplitProtocol/Sample/$exit
      -- CP-element group 273: 	 branch_block_stmt_216/forx_xbody_forx_xbody_PhiReq/phi_stmt_555/phi_stmt_555_sources/type_cast_561/SplitProtocol/Sample/ra
      -- 
    ra_2763_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 273_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_561_inst_ack_0, ack => concat_CP_664_elements(273)); -- 
    -- CP-element group 274:  transition  input  bypass 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	127 
    -- CP-element group 274: successors 
    -- CP-element group 274: 	275 
    -- CP-element group 274:  members (2) 
      -- CP-element group 274: 	 branch_block_stmt_216/forx_xbody_forx_xbody_PhiReq/phi_stmt_555/phi_stmt_555_sources/type_cast_561/SplitProtocol/Update/$exit
      -- CP-element group 274: 	 branch_block_stmt_216/forx_xbody_forx_xbody_PhiReq/phi_stmt_555/phi_stmt_555_sources/type_cast_561/SplitProtocol/Update/ca
      -- 
    ca_2768_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 274_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_561_inst_ack_1, ack => concat_CP_664_elements(274)); -- 
    -- CP-element group 275:  join  transition  output  bypass 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	273 
    -- CP-element group 275: 	274 
    -- CP-element group 275: successors 
    -- CP-element group 275: 	276 
    -- CP-element group 275:  members (6) 
      -- CP-element group 275: 	 branch_block_stmt_216/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 275: 	 branch_block_stmt_216/forx_xbody_forx_xbody_PhiReq/phi_stmt_555/$exit
      -- CP-element group 275: 	 branch_block_stmt_216/forx_xbody_forx_xbody_PhiReq/phi_stmt_555/phi_stmt_555_sources/$exit
      -- CP-element group 275: 	 branch_block_stmt_216/forx_xbody_forx_xbody_PhiReq/phi_stmt_555/phi_stmt_555_sources/type_cast_561/$exit
      -- CP-element group 275: 	 branch_block_stmt_216/forx_xbody_forx_xbody_PhiReq/phi_stmt_555/phi_stmt_555_sources/type_cast_561/SplitProtocol/$exit
      -- CP-element group 275: 	 branch_block_stmt_216/forx_xbody_forx_xbody_PhiReq/phi_stmt_555/phi_stmt_555_req
      -- 
    phi_stmt_555_req_2769_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_555_req_2769_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(275), ack => phi_stmt_555_req_1); -- 
    concat_cp_element_group_275: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_275"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_664_elements(273) & concat_CP_664_elements(274);
      gj_concat_cp_element_group_275 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_664_elements(275), clk => clk, reset => reset); --
    end block;
    -- CP-element group 276:  merge  transition  place  bypass 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	272 
    -- CP-element group 276: 	275 
    -- CP-element group 276: successors 
    -- CP-element group 276: 	277 
    -- CP-element group 276:  members (2) 
      -- CP-element group 276: 	 branch_block_stmt_216/merge_stmt_554_PhiReqMerge
      -- CP-element group 276: 	 branch_block_stmt_216/merge_stmt_554_PhiAck/$entry
      -- 
    concat_CP_664_elements(276) <= OrReduce(concat_CP_664_elements(272) & concat_CP_664_elements(275));
    -- CP-element group 277:  fork  transition  place  input  output  bypass 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	276 
    -- CP-element group 277: successors 
    -- CP-element group 277: 	86 
    -- CP-element group 277: 	87 
    -- CP-element group 277: 	89 
    -- CP-element group 277: 	90 
    -- CP-element group 277: 	93 
    -- CP-element group 277: 	97 
    -- CP-element group 277: 	101 
    -- CP-element group 277: 	105 
    -- CP-element group 277: 	109 
    -- CP-element group 277: 	113 
    -- CP-element group 277: 	117 
    -- CP-element group 277: 	121 
    -- CP-element group 277: 	124 
    -- CP-element group 277:  members (56) 
      -- CP-element group 277: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/array_obj_ref_569_final_index_sum_regn_update_start
      -- CP-element group 277: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_626_update_start_
      -- CP-element group 277: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_577_Update/cr
      -- CP-element group 277: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_662_update_start_
      -- CP-element group 277: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_680_Update/cr
      -- CP-element group 277: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_577_Update/$entry
      -- CP-element group 277: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/ptr_deref_706_Update/word_access_complete/$entry
      -- CP-element group 277: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_644_Update/$entry
      -- CP-element group 277: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/array_obj_ref_569_final_index_sum_regn_Update/$entry
      -- CP-element group 277: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/array_obj_ref_569_index_scale_2/scale_rename_req
      -- CP-element group 277: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/ptr_deref_706_Update/word_access_complete/word_0/$entry
      -- CP-element group 277: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/array_obj_ref_569_index_resize_2/index_resize_ack
      -- CP-element group 277: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_608_Update/$entry
      -- CP-element group 277: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/array_obj_ref_569_index_resize_2/$exit
      -- CP-element group 277: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/addr_of_570_complete/req
      -- CP-element group 277: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/ptr_deref_706_update_start_
      -- CP-element group 277: 	 branch_block_stmt_216/merge_stmt_554__exit__
      -- CP-element group 277: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719__entry__
      -- CP-element group 277: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/array_obj_ref_569_index_scale_2/$exit
      -- CP-element group 277: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_573_Sample/$entry
      -- CP-element group 277: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_698_Update/$entry
      -- CP-element group 277: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_698_Update/cr
      -- CP-element group 277: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_680_Update/$entry
      -- CP-element group 277: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/array_obj_ref_569_index_resize_2/index_resize_req
      -- CP-element group 277: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_573_Sample/rr
      -- CP-element group 277: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/array_obj_ref_569_index_scale_2/scale_rename_ack
      -- CP-element group 277: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/ptr_deref_706_Update/word_access_complete/word_0/cr
      -- CP-element group 277: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_608_Update/cr
      -- CP-element group 277: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_644_update_start_
      -- CP-element group 277: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/array_obj_ref_569_index_resize_2/$entry
      -- CP-element group 277: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/RPIPE_Concat_input_pipe_573_sample_start_
      -- CP-element group 277: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/array_obj_ref_569_final_index_sum_regn_Sample/$entry
      -- CP-element group 277: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_644_Update/cr
      -- CP-element group 277: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/array_obj_ref_569_final_index_sum_regn_Update/req
      -- CP-element group 277: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_680_update_start_
      -- CP-element group 277: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/array_obj_ref_569_index_scale_2/$entry
      -- CP-element group 277: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_577_update_start_
      -- CP-element group 277: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/array_obj_ref_569_final_index_sum_regn_Sample/req
      -- CP-element group 277: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/ptr_deref_706_Update/$entry
      -- CP-element group 277: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/addr_of_570_complete/$entry
      -- CP-element group 277: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_608_update_start_
      -- CP-element group 277: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/array_obj_ref_569_index_computed_2
      -- CP-element group 277: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/array_obj_ref_569_index_scaled_2
      -- CP-element group 277: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/array_obj_ref_569_index_resized_2
      -- CP-element group 277: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_698_update_start_
      -- CP-element group 277: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_626_Update/cr
      -- CP-element group 277: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/addr_of_570_update_start_
      -- CP-element group 277: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_626_Update/$entry
      -- CP-element group 277: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_590_Update/cr
      -- CP-element group 277: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_662_Update/cr
      -- CP-element group 277: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/$entry
      -- CP-element group 277: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_590_Update/$entry
      -- CP-element group 277: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_590_update_start_
      -- CP-element group 277: 	 branch_block_stmt_216/assign_stmt_571_to_assign_stmt_719/type_cast_662_Update/$entry
      -- CP-element group 277: 	 branch_block_stmt_216/merge_stmt_554_PhiAck/$exit
      -- CP-element group 277: 	 branch_block_stmt_216/merge_stmt_554_PhiAck/phi_stmt_555_ack
      -- 
    phi_stmt_555_ack_2774_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 277_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_555_ack_0, ack => concat_CP_664_elements(277)); -- 
    cr_1402_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1402_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(277), ack => type_cast_577_inst_req_1); -- 
    cr_1570_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1570_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(277), ack => type_cast_680_inst_req_1); -- 
    req_1374_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1374_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(277), ack => addr_of_570_final_reg_req_1); -- 
    cr_1598_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1598_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(277), ack => type_cast_698_inst_req_1); -- 
    rr_1383_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1383_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(277), ack => RPIPE_Concat_input_pipe_573_inst_req_0); -- 
    cr_1648_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1648_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(277), ack => ptr_deref_706_store_0_req_1); -- 
    cr_1458_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1458_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(277), ack => type_cast_608_inst_req_1); -- 
    cr_1514_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1514_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(277), ack => type_cast_644_inst_req_1); -- 
    req_1359_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1359_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(277), ack => array_obj_ref_569_index_offset_req_1); -- 
    req_1354_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1354_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(277), ack => array_obj_ref_569_index_offset_req_0); -- 
    cr_1486_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1486_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(277), ack => type_cast_626_inst_req_1); -- 
    cr_1430_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1430_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(277), ack => type_cast_590_inst_req_1); -- 
    cr_1542_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1542_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(277), ack => type_cast_662_inst_req_1); -- 
    -- CP-element group 278:  transition  output  delay-element  bypass 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	129 
    -- CP-element group 278: successors 
    -- CP-element group 278: 	282 
    -- CP-element group 278:  members (5) 
      -- CP-element group 278: 	 branch_block_stmt_216/bbx_xnph386_forx_xbody171_PhiReq/$exit
      -- CP-element group 278: 	 branch_block_stmt_216/bbx_xnph386_forx_xbody171_PhiReq/phi_stmt_762/$exit
      -- CP-element group 278: 	 branch_block_stmt_216/bbx_xnph386_forx_xbody171_PhiReq/phi_stmt_762/phi_stmt_762_sources/$exit
      -- CP-element group 278: 	 branch_block_stmt_216/bbx_xnph386_forx_xbody171_PhiReq/phi_stmt_762/phi_stmt_762_sources/type_cast_766_konst_delay_trans
      -- CP-element group 278: 	 branch_block_stmt_216/bbx_xnph386_forx_xbody171_PhiReq/phi_stmt_762/phi_stmt_762_req
      -- 
    phi_stmt_762_req_2797_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_762_req_2797_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(278), ack => phi_stmt_762_req_0); -- 
    -- Element group concat_CP_664_elements(278) is a control-delay.
    cp_element_278_delay: control_delay_element  generic map(name => " 278_delay", delay_value => 1)  port map(req => concat_CP_664_elements(129), ack => concat_CP_664_elements(278), clk => clk, reset =>reset);
    -- CP-element group 279:  transition  input  bypass 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	171 
    -- CP-element group 279: successors 
    -- CP-element group 279: 	281 
    -- CP-element group 279:  members (2) 
      -- CP-element group 279: 	 branch_block_stmt_216/forx_xbody171_forx_xbody171_PhiReq/phi_stmt_762/phi_stmt_762_sources/type_cast_768/SplitProtocol/Sample/$exit
      -- CP-element group 279: 	 branch_block_stmt_216/forx_xbody171_forx_xbody171_PhiReq/phi_stmt_762/phi_stmt_762_sources/type_cast_768/SplitProtocol/Sample/ra
      -- 
    ra_2817_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 279_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_768_inst_ack_0, ack => concat_CP_664_elements(279)); -- 
    -- CP-element group 280:  transition  input  bypass 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	171 
    -- CP-element group 280: successors 
    -- CP-element group 280: 	281 
    -- CP-element group 280:  members (2) 
      -- CP-element group 280: 	 branch_block_stmt_216/forx_xbody171_forx_xbody171_PhiReq/phi_stmt_762/phi_stmt_762_sources/type_cast_768/SplitProtocol/Update/$exit
      -- CP-element group 280: 	 branch_block_stmt_216/forx_xbody171_forx_xbody171_PhiReq/phi_stmt_762/phi_stmt_762_sources/type_cast_768/SplitProtocol/Update/ca
      -- 
    ca_2822_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 280_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_768_inst_ack_1, ack => concat_CP_664_elements(280)); -- 
    -- CP-element group 281:  join  transition  output  bypass 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	279 
    -- CP-element group 281: 	280 
    -- CP-element group 281: successors 
    -- CP-element group 281: 	282 
    -- CP-element group 281:  members (6) 
      -- CP-element group 281: 	 branch_block_stmt_216/forx_xbody171_forx_xbody171_PhiReq/$exit
      -- CP-element group 281: 	 branch_block_stmt_216/forx_xbody171_forx_xbody171_PhiReq/phi_stmt_762/$exit
      -- CP-element group 281: 	 branch_block_stmt_216/forx_xbody171_forx_xbody171_PhiReq/phi_stmt_762/phi_stmt_762_sources/$exit
      -- CP-element group 281: 	 branch_block_stmt_216/forx_xbody171_forx_xbody171_PhiReq/phi_stmt_762/phi_stmt_762_sources/type_cast_768/$exit
      -- CP-element group 281: 	 branch_block_stmt_216/forx_xbody171_forx_xbody171_PhiReq/phi_stmt_762/phi_stmt_762_sources/type_cast_768/SplitProtocol/$exit
      -- CP-element group 281: 	 branch_block_stmt_216/forx_xbody171_forx_xbody171_PhiReq/phi_stmt_762/phi_stmt_762_req
      -- 
    phi_stmt_762_req_2823_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_762_req_2823_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(281), ack => phi_stmt_762_req_1); -- 
    concat_cp_element_group_281: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_281"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_664_elements(279) & concat_CP_664_elements(280);
      gj_concat_cp_element_group_281 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_664_elements(281), clk => clk, reset => reset); --
    end block;
    -- CP-element group 282:  merge  transition  place  bypass 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	278 
    -- CP-element group 282: 	281 
    -- CP-element group 282: successors 
    -- CP-element group 282: 	283 
    -- CP-element group 282:  members (2) 
      -- CP-element group 282: 	 branch_block_stmt_216/merge_stmt_761_PhiReqMerge
      -- CP-element group 282: 	 branch_block_stmt_216/merge_stmt_761_PhiAck/$entry
      -- 
    concat_CP_664_elements(282) <= OrReduce(concat_CP_664_elements(278) & concat_CP_664_elements(281));
    -- CP-element group 283:  fork  transition  place  input  output  bypass 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: 	282 
    -- CP-element group 283: successors 
    -- CP-element group 283: 	130 
    -- CP-element group 283: 	131 
    -- CP-element group 283: 	133 
    -- CP-element group 283: 	134 
    -- CP-element group 283: 	137 
    -- CP-element group 283: 	141 
    -- CP-element group 283: 	145 
    -- CP-element group 283: 	149 
    -- CP-element group 283: 	153 
    -- CP-element group 283: 	157 
    -- CP-element group 283: 	161 
    -- CP-element group 283: 	165 
    -- CP-element group 283: 	168 
    -- CP-element group 283:  members (56) 
      -- CP-element group 283: 	 branch_block_stmt_216/merge_stmt_761__exit__
      -- CP-element group 283: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926__entry__
      -- CP-element group 283: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/$entry
      -- CP-element group 283: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/addr_of_777_update_start_
      -- CP-element group 283: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/array_obj_ref_776_index_resized_2
      -- CP-element group 283: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/array_obj_ref_776_index_scaled_2
      -- CP-element group 283: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/array_obj_ref_776_index_computed_2
      -- CP-element group 283: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/array_obj_ref_776_index_resize_2/$entry
      -- CP-element group 283: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/array_obj_ref_776_index_resize_2/$exit
      -- CP-element group 283: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/array_obj_ref_776_index_resize_2/index_resize_req
      -- CP-element group 283: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/array_obj_ref_776_index_resize_2/index_resize_ack
      -- CP-element group 283: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/array_obj_ref_776_index_scale_2/$entry
      -- CP-element group 283: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/array_obj_ref_776_index_scale_2/$exit
      -- CP-element group 283: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/array_obj_ref_776_index_scale_2/scale_rename_req
      -- CP-element group 283: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/array_obj_ref_776_index_scale_2/scale_rename_ack
      -- CP-element group 283: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/array_obj_ref_776_final_index_sum_regn_update_start
      -- CP-element group 283: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/array_obj_ref_776_final_index_sum_regn_Sample/$entry
      -- CP-element group 283: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/array_obj_ref_776_final_index_sum_regn_Sample/req
      -- CP-element group 283: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/array_obj_ref_776_final_index_sum_regn_Update/$entry
      -- CP-element group 283: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/array_obj_ref_776_final_index_sum_regn_Update/req
      -- CP-element group 283: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/addr_of_777_complete/$entry
      -- CP-element group 283: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/addr_of_777_complete/req
      -- CP-element group 283: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_780_sample_start_
      -- CP-element group 283: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_780_Sample/$entry
      -- CP-element group 283: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/RPIPE_Concat_input_pipe_780_Sample/rr
      -- CP-element group 283: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_784_update_start_
      -- CP-element group 283: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_784_Update/$entry
      -- CP-element group 283: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_784_Update/cr
      -- CP-element group 283: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_797_update_start_
      -- CP-element group 283: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_797_Update/$entry
      -- CP-element group 283: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_797_Update/cr
      -- CP-element group 283: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_815_update_start_
      -- CP-element group 283: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_815_Update/$entry
      -- CP-element group 283: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_815_Update/cr
      -- CP-element group 283: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_833_update_start_
      -- CP-element group 283: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_833_Update/$entry
      -- CP-element group 283: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_833_Update/cr
      -- CP-element group 283: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_851_update_start_
      -- CP-element group 283: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_851_Update/$entry
      -- CP-element group 283: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_851_Update/cr
      -- CP-element group 283: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_869_update_start_
      -- CP-element group 283: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_869_Update/$entry
      -- CP-element group 283: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_869_Update/cr
      -- CP-element group 283: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_887_update_start_
      -- CP-element group 283: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_887_Update/$entry
      -- CP-element group 283: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_887_Update/cr
      -- CP-element group 283: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_905_update_start_
      -- CP-element group 283: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_905_Update/$entry
      -- CP-element group 283: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/type_cast_905_Update/cr
      -- CP-element group 283: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_update_start_
      -- CP-element group 283: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_Update/$entry
      -- CP-element group 283: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_Update/word_access_complete/$entry
      -- CP-element group 283: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_Update/word_access_complete/word_0/$entry
      -- CP-element group 283: 	 branch_block_stmt_216/assign_stmt_778_to_assign_stmt_926/ptr_deref_913_Update/word_access_complete/word_0/cr
      -- CP-element group 283: 	 branch_block_stmt_216/merge_stmt_761_PhiAck/$exit
      -- CP-element group 283: 	 branch_block_stmt_216/merge_stmt_761_PhiAck/phi_stmt_762_ack
      -- 
    phi_stmt_762_ack_2828_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 283_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_762_ack_0, ack => concat_CP_664_elements(283)); -- 
    req_1713_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1713_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(283), ack => array_obj_ref_776_index_offset_req_0); -- 
    req_1718_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1718_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(283), ack => array_obj_ref_776_index_offset_req_1); -- 
    req_1733_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1733_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(283), ack => addr_of_777_final_reg_req_1); -- 
    rr_1742_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1742_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(283), ack => RPIPE_Concat_input_pipe_780_inst_req_0); -- 
    cr_1761_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1761_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(283), ack => type_cast_784_inst_req_1); -- 
    cr_1789_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1789_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(283), ack => type_cast_797_inst_req_1); -- 
    cr_1817_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1817_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(283), ack => type_cast_815_inst_req_1); -- 
    cr_1845_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1845_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(283), ack => type_cast_833_inst_req_1); -- 
    cr_1873_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1873_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(283), ack => type_cast_851_inst_req_1); -- 
    cr_1901_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1901_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(283), ack => type_cast_869_inst_req_1); -- 
    cr_1929_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1929_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(283), ack => type_cast_887_inst_req_1); -- 
    cr_1957_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1957_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(283), ack => type_cast_905_inst_req_1); -- 
    cr_2007_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2007_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(283), ack => ptr_deref_913_store_0_req_1); -- 
    -- CP-element group 284:  merge  fork  transition  place  output  bypass 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	83 
    -- CP-element group 284: 	170 
    -- CP-element group 284: successors 
    -- CP-element group 284: 	172 
    -- CP-element group 284: 	173 
    -- CP-element group 284: 	175 
    -- CP-element group 284:  members (16) 
      -- CP-element group 284: 	 branch_block_stmt_216/call_stmt_938_to_assign_stmt_944__entry__
      -- CP-element group 284: 	 branch_block_stmt_216/merge_stmt_935__exit__
      -- CP-element group 284: 	 branch_block_stmt_216/call_stmt_938_to_assign_stmt_944/$entry
      -- CP-element group 284: 	 branch_block_stmt_216/call_stmt_938_to_assign_stmt_944/call_stmt_938_sample_start_
      -- CP-element group 284: 	 branch_block_stmt_216/call_stmt_938_to_assign_stmt_944/call_stmt_938_update_start_
      -- CP-element group 284: 	 branch_block_stmt_216/call_stmt_938_to_assign_stmt_944/call_stmt_938_Sample/$entry
      -- CP-element group 284: 	 branch_block_stmt_216/call_stmt_938_to_assign_stmt_944/call_stmt_938_Sample/crr
      -- CP-element group 284: 	 branch_block_stmt_216/call_stmt_938_to_assign_stmt_944/call_stmt_938_Update/$entry
      -- CP-element group 284: 	 branch_block_stmt_216/call_stmt_938_to_assign_stmt_944/call_stmt_938_Update/ccr
      -- CP-element group 284: 	 branch_block_stmt_216/call_stmt_938_to_assign_stmt_944/type_cast_943_update_start_
      -- CP-element group 284: 	 branch_block_stmt_216/call_stmt_938_to_assign_stmt_944/type_cast_943_Update/$entry
      -- CP-element group 284: 	 branch_block_stmt_216/call_stmt_938_to_assign_stmt_944/type_cast_943_Update/cr
      -- CP-element group 284: 	 branch_block_stmt_216/merge_stmt_935_PhiReqMerge
      -- CP-element group 284: 	 branch_block_stmt_216/merge_stmt_935_PhiAck/$entry
      -- CP-element group 284: 	 branch_block_stmt_216/merge_stmt_935_PhiAck/$exit
      -- CP-element group 284: 	 branch_block_stmt_216/merge_stmt_935_PhiAck/dummy
      -- 
    crr_2038_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2038_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(284), ack => call_stmt_938_call_req_0); -- 
    ccr_2043_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2043_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(284), ack => call_stmt_938_call_req_1); -- 
    cr_2057_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2057_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(284), ack => type_cast_943_inst_req_1); -- 
    concat_CP_664_elements(284) <= OrReduce(concat_CP_664_elements(83) & concat_CP_664_elements(170));
    -- CP-element group 285:  transition  output  delay-element  bypass 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: 	221 
    -- CP-element group 285: successors 
    -- CP-element group 285: 	289 
    -- CP-element group 285:  members (5) 
      -- CP-element group 285: 	 branch_block_stmt_216/bbx_xnph_forx_xbody305_PhiReq/$exit
      -- CP-element group 285: 	 branch_block_stmt_216/bbx_xnph_forx_xbody305_PhiReq/phi_stmt_1106/$exit
      -- CP-element group 285: 	 branch_block_stmt_216/bbx_xnph_forx_xbody305_PhiReq/phi_stmt_1106/phi_stmt_1106_sources/$exit
      -- CP-element group 285: 	 branch_block_stmt_216/bbx_xnph_forx_xbody305_PhiReq/phi_stmt_1106/phi_stmt_1106_sources/type_cast_1110_konst_delay_trans
      -- CP-element group 285: 	 branch_block_stmt_216/bbx_xnph_forx_xbody305_PhiReq/phi_stmt_1106/phi_stmt_1106_req
      -- 
    phi_stmt_1106_req_2874_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1106_req_2874_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(285), ack => phi_stmt_1106_req_0); -- 
    -- Element group concat_CP_664_elements(285) is a control-delay.
    cp_element_285_delay: control_delay_element  generic map(name => " 285_delay", delay_value => 1)  port map(req => concat_CP_664_elements(221), ack => concat_CP_664_elements(285), clk => clk, reset =>reset);
    -- CP-element group 286:  transition  input  bypass 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	270 
    -- CP-element group 286: successors 
    -- CP-element group 286: 	288 
    -- CP-element group 286:  members (2) 
      -- CP-element group 286: 	 branch_block_stmt_216/forx_xbody305_forx_xbody305_PhiReq/phi_stmt_1106/phi_stmt_1106_sources/type_cast_1112/SplitProtocol/Sample/$exit
      -- CP-element group 286: 	 branch_block_stmt_216/forx_xbody305_forx_xbody305_PhiReq/phi_stmt_1106/phi_stmt_1106_sources/type_cast_1112/SplitProtocol/Sample/ra
      -- 
    ra_2894_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 286_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1112_inst_ack_0, ack => concat_CP_664_elements(286)); -- 
    -- CP-element group 287:  transition  input  bypass 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	270 
    -- CP-element group 287: successors 
    -- CP-element group 287: 	288 
    -- CP-element group 287:  members (2) 
      -- CP-element group 287: 	 branch_block_stmt_216/forx_xbody305_forx_xbody305_PhiReq/phi_stmt_1106/phi_stmt_1106_sources/type_cast_1112/SplitProtocol/Update/$exit
      -- CP-element group 287: 	 branch_block_stmt_216/forx_xbody305_forx_xbody305_PhiReq/phi_stmt_1106/phi_stmt_1106_sources/type_cast_1112/SplitProtocol/Update/ca
      -- 
    ca_2899_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 287_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1112_inst_ack_1, ack => concat_CP_664_elements(287)); -- 
    -- CP-element group 288:  join  transition  output  bypass 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	286 
    -- CP-element group 288: 	287 
    -- CP-element group 288: successors 
    -- CP-element group 288: 	289 
    -- CP-element group 288:  members (6) 
      -- CP-element group 288: 	 branch_block_stmt_216/forx_xbody305_forx_xbody305_PhiReq/$exit
      -- CP-element group 288: 	 branch_block_stmt_216/forx_xbody305_forx_xbody305_PhiReq/phi_stmt_1106/$exit
      -- CP-element group 288: 	 branch_block_stmt_216/forx_xbody305_forx_xbody305_PhiReq/phi_stmt_1106/phi_stmt_1106_sources/$exit
      -- CP-element group 288: 	 branch_block_stmt_216/forx_xbody305_forx_xbody305_PhiReq/phi_stmt_1106/phi_stmt_1106_sources/type_cast_1112/$exit
      -- CP-element group 288: 	 branch_block_stmt_216/forx_xbody305_forx_xbody305_PhiReq/phi_stmt_1106/phi_stmt_1106_sources/type_cast_1112/SplitProtocol/$exit
      -- CP-element group 288: 	 branch_block_stmt_216/forx_xbody305_forx_xbody305_PhiReq/phi_stmt_1106/phi_stmt_1106_req
      -- 
    phi_stmt_1106_req_2900_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1106_req_2900_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(288), ack => phi_stmt_1106_req_1); -- 
    concat_cp_element_group_288: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "concat_cp_element_group_288"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_CP_664_elements(286) & concat_CP_664_elements(287);
      gj_concat_cp_element_group_288 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_CP_664_elements(288), clk => clk, reset => reset); --
    end block;
    -- CP-element group 289:  merge  transition  place  bypass 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: 	285 
    -- CP-element group 289: 	288 
    -- CP-element group 289: successors 
    -- CP-element group 289: 	290 
    -- CP-element group 289:  members (2) 
      -- CP-element group 289: 	 branch_block_stmt_216/merge_stmt_1105_PhiReqMerge
      -- CP-element group 289: 	 branch_block_stmt_216/merge_stmt_1105_PhiAck/$entry
      -- 
    concat_CP_664_elements(289) <= OrReduce(concat_CP_664_elements(285) & concat_CP_664_elements(288));
    -- CP-element group 290:  fork  transition  place  input  output  bypass 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: 	289 
    -- CP-element group 290: successors 
    -- CP-element group 290: 	223 
    -- CP-element group 290: 	224 
    -- CP-element group 290: 	226 
    -- CP-element group 290: 	228 
    -- CP-element group 290: 	230 
    -- CP-element group 290: 	232 
    -- CP-element group 290: 	234 
    -- CP-element group 290: 	236 
    -- CP-element group 290: 	238 
    -- CP-element group 290: 	240 
    -- CP-element group 290: 	242 
    -- CP-element group 290: 	244 
    -- CP-element group 290:  members (53) 
      -- CP-element group 290: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235__entry__
      -- CP-element group 290: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/array_obj_ref_1120_final_index_sum_regn_Sample/req
      -- CP-element group 290: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/addr_of_1121_complete/$entry
      -- CP-element group 290: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/array_obj_ref_1120_final_index_sum_regn_update_start
      -- CP-element group 290: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/array_obj_ref_1120_final_index_sum_regn_Sample/$entry
      -- CP-element group 290: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1169_Update/$entry
      -- CP-element group 290: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1139_Update/cr
      -- CP-element group 290: 	 branch_block_stmt_216/merge_stmt_1105__exit__
      -- CP-element group 290: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1139_Update/$entry
      -- CP-element group 290: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/array_obj_ref_1120_final_index_sum_regn_Update/$entry
      -- CP-element group 290: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1179_update_start_
      -- CP-element group 290: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1169_Update/cr
      -- CP-element group 290: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1149_update_start_
      -- CP-element group 290: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/array_obj_ref_1120_final_index_sum_regn_Update/req
      -- CP-element group 290: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1199_Update/$entry
      -- CP-element group 290: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1179_Update/$entry
      -- CP-element group 290: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/addr_of_1121_complete/req
      -- CP-element group 290: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1179_Update/cr
      -- CP-element group 290: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/ptr_deref_1125_update_start_
      -- CP-element group 290: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1149_Update/$entry
      -- CP-element group 290: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1149_Update/cr
      -- CP-element group 290: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1199_Update/cr
      -- CP-element group 290: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1159_update_start_
      -- CP-element group 290: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/array_obj_ref_1120_index_scale_2/scale_rename_ack
      -- CP-element group 290: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/array_obj_ref_1120_index_scale_2/scale_rename_req
      -- CP-element group 290: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/array_obj_ref_1120_index_scale_2/$exit
      -- CP-element group 290: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/array_obj_ref_1120_index_scale_2/$entry
      -- CP-element group 290: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/array_obj_ref_1120_index_resize_2/index_resize_ack
      -- CP-element group 290: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/array_obj_ref_1120_index_resize_2/index_resize_req
      -- CP-element group 290: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/array_obj_ref_1120_index_resize_2/$exit
      -- CP-element group 290: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/array_obj_ref_1120_index_resize_2/$entry
      -- CP-element group 290: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1139_update_start_
      -- CP-element group 290: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/array_obj_ref_1120_index_computed_2
      -- CP-element group 290: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/array_obj_ref_1120_index_scaled_2
      -- CP-element group 290: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/array_obj_ref_1120_index_resized_2
      -- CP-element group 290: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/addr_of_1121_update_start_
      -- CP-element group 290: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1129_Update/cr
      -- CP-element group 290: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1129_Update/$entry
      -- CP-element group 290: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1169_update_start_
      -- CP-element group 290: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/$entry
      -- CP-element group 290: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1199_update_start_
      -- CP-element group 290: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1129_update_start_
      -- CP-element group 290: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1159_Update/cr
      -- CP-element group 290: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1159_Update/$entry
      -- CP-element group 290: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1189_Update/cr
      -- CP-element group 290: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1189_Update/$entry
      -- CP-element group 290: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/ptr_deref_1125_Update/word_access_complete/word_0/cr
      -- CP-element group 290: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/ptr_deref_1125_Update/word_access_complete/word_0/$entry
      -- CP-element group 290: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/ptr_deref_1125_Update/word_access_complete/$entry
      -- CP-element group 290: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/type_cast_1189_update_start_
      -- CP-element group 290: 	 branch_block_stmt_216/assign_stmt_1122_to_assign_stmt_1235/ptr_deref_1125_Update/$entry
      -- CP-element group 290: 	 branch_block_stmt_216/merge_stmt_1105_PhiAck/$exit
      -- CP-element group 290: 	 branch_block_stmt_216/merge_stmt_1105_PhiAck/phi_stmt_1106_ack
      -- 
    phi_stmt_1106_ack_2905_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 290_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1106_ack_0, ack => concat_CP_664_elements(290)); -- 
    req_2383_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2383_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(290), ack => array_obj_ref_1120_index_offset_req_0); -- 
    cr_2481_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2481_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(290), ack => type_cast_1139_inst_req_1); -- 
    cr_2523_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2523_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(290), ack => type_cast_1169_inst_req_1); -- 
    req_2388_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2388_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(290), ack => array_obj_ref_1120_index_offset_req_1); -- 
    req_2403_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2403_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(290), ack => addr_of_1121_final_reg_req_1); -- 
    cr_2537_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2537_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(290), ack => type_cast_1179_inst_req_1); -- 
    cr_2495_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2495_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(290), ack => type_cast_1149_inst_req_1); -- 
    cr_2565_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2565_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(290), ack => type_cast_1199_inst_req_1); -- 
    cr_2467_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2467_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(290), ack => type_cast_1129_inst_req_1); -- 
    cr_2509_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2509_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(290), ack => type_cast_1159_inst_req_1); -- 
    cr_2551_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2551_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(290), ack => type_cast_1189_inst_req_1); -- 
    cr_2448_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2448_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_CP_664_elements(290), ack => ptr_deref_1125_load_0_req_1); -- 
    -- CP-element group 291:  merge  transition  place  bypass 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	269 
    -- CP-element group 291: 	222 
    -- CP-element group 291: successors 
    -- CP-element group 291:  members (16) 
      -- CP-element group 291: 	 branch_block_stmt_216/$exit
      -- CP-element group 291: 	 branch_block_stmt_216/branch_block_stmt_216__exit__
      -- CP-element group 291: 	 $exit
      -- CP-element group 291: 	 branch_block_stmt_216/merge_stmt_1244__exit__
      -- CP-element group 291: 	 branch_block_stmt_216/return__
      -- CP-element group 291: 	 branch_block_stmt_216/merge_stmt_1246__exit__
      -- CP-element group 291: 	 branch_block_stmt_216/merge_stmt_1244_PhiReqMerge
      -- CP-element group 291: 	 branch_block_stmt_216/merge_stmt_1244_PhiAck/$entry
      -- CP-element group 291: 	 branch_block_stmt_216/merge_stmt_1244_PhiAck/$exit
      -- CP-element group 291: 	 branch_block_stmt_216/merge_stmt_1244_PhiAck/dummy
      -- CP-element group 291: 	 branch_block_stmt_216/return___PhiReq/$entry
      -- CP-element group 291: 	 branch_block_stmt_216/return___PhiReq/$exit
      -- CP-element group 291: 	 branch_block_stmt_216/merge_stmt_1246_PhiReqMerge
      -- CP-element group 291: 	 branch_block_stmt_216/merge_stmt_1246_PhiAck/$entry
      -- CP-element group 291: 	 branch_block_stmt_216/merge_stmt_1246_PhiAck/$exit
      -- CP-element group 291: 	 branch_block_stmt_216/merge_stmt_1246_PhiAck/dummy
      -- 
    concat_CP_664_elements(291) <= OrReduce(concat_CP_664_elements(269) & concat_CP_664_elements(222));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_ix_x0389_568_resized : std_logic_vector(15 downto 0);
    signal R_ix_x0389_568_scaled : std_logic_vector(15 downto 0);
    signal R_ix_x1385_775_resized : std_logic_vector(15 downto 0);
    signal R_ix_x1385_775_scaled : std_logic_vector(15 downto 0);
    signal R_ix_x2382_1119_resized : std_logic_vector(15 downto 0);
    signal R_ix_x2382_1119_scaled : std_logic_vector(15 downto 0);
    signal add125_596 : std_logic_vector(63 downto 0);
    signal add12_266 : std_logic_vector(31 downto 0);
    signal add131_614 : std_logic_vector(63 downto 0);
    signal add137_632 : std_logic_vector(63 downto 0);
    signal add143_650 : std_logic_vector(63 downto 0);
    signal add149_668 : std_logic_vector(63 downto 0);
    signal add155_686 : std_logic_vector(63 downto 0);
    signal add161_704 : std_logic_vector(63 downto 0);
    signal add181_803 : std_logic_vector(63 downto 0);
    signal add187_821 : std_logic_vector(63 downto 0);
    signal add193_839 : std_logic_vector(63 downto 0);
    signal add199_857 : std_logic_vector(63 downto 0);
    signal add205_875 : std_logic_vector(63 downto 0);
    signal add211_893 : std_logic_vector(63 downto 0);
    signal add217_911 : std_logic_vector(63 downto 0);
    signal add21_291 : std_logic_vector(15 downto 0);
    signal add30_316 : std_logic_vector(31 downto 0);
    signal add39_341 : std_logic_vector(31 downto 0);
    signal add48_366 : std_logic_vector(15 downto 0);
    signal add57_391 : std_logic_vector(31 downto 0);
    signal add66_416 : std_logic_vector(31 downto 0);
    signal add75_441 : std_logic_vector(31 downto 0);
    signal add_241 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1120_constant_part_of_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_1120_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_1120_offset_scale_factor_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1120_offset_scale_factor_1 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1120_offset_scale_factor_2 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1120_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_1120_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_569_constant_part_of_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_569_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_569_offset_scale_factor_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_569_offset_scale_factor_1 : std_logic_vector(15 downto 0);
    signal array_obj_ref_569_offset_scale_factor_2 : std_logic_vector(15 downto 0);
    signal array_obj_ref_569_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_569_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_776_constant_part_of_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_776_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_776_offset_scale_factor_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_776_offset_scale_factor_1 : std_logic_vector(15 downto 0);
    signal array_obj_ref_776_offset_scale_factor_2 : std_logic_vector(15 downto 0);
    signal array_obj_ref_776_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_776_root_address : std_logic_vector(15 downto 0);
    signal arrayidx220_778 : std_logic_vector(31 downto 0);
    signal arrayidx309_1122 : std_logic_vector(31 downto 0);
    signal arrayidx_571 : std_logic_vector(31 downto 0);
    signal call10_257 : std_logic_vector(7 downto 0);
    signal call118_574 : std_logic_vector(7 downto 0);
    signal call122_587 : std_logic_vector(7 downto 0);
    signal call128_605 : std_logic_vector(7 downto 0);
    signal call134_623 : std_logic_vector(7 downto 0);
    signal call140_641 : std_logic_vector(7 downto 0);
    signal call146_659 : std_logic_vector(7 downto 0);
    signal call14_269 : std_logic_vector(7 downto 0);
    signal call152_677 : std_logic_vector(7 downto 0);
    signal call158_695 : std_logic_vector(7 downto 0);
    signal call174_781 : std_logic_vector(7 downto 0);
    signal call178_794 : std_logic_vector(7 downto 0);
    signal call184_812 : std_logic_vector(7 downto 0);
    signal call190_830 : std_logic_vector(7 downto 0);
    signal call196_848 : std_logic_vector(7 downto 0);
    signal call19_282 : std_logic_vector(7 downto 0);
    signal call202_866 : std_logic_vector(7 downto 0);
    signal call208_884 : std_logic_vector(7 downto 0);
    signal call214_902 : std_logic_vector(7 downto 0);
    signal call226_938 : std_logic_vector(63 downto 0);
    signal call232_952 : std_logic_vector(63 downto 0);
    signal call23_294 : std_logic_vector(7 downto 0);
    signal call28_307 : std_logic_vector(7 downto 0);
    signal call2_232 : std_logic_vector(7 downto 0);
    signal call32_319 : std_logic_vector(7 downto 0);
    signal call37_332 : std_logic_vector(7 downto 0);
    signal call41_344 : std_logic_vector(7 downto 0);
    signal call46_357 : std_logic_vector(7 downto 0);
    signal call50_369 : std_logic_vector(7 downto 0);
    signal call55_382 : std_logic_vector(7 downto 0);
    signal call59_394 : std_logic_vector(7 downto 0);
    signal call5_244 : std_logic_vector(7 downto 0);
    signal call64_407 : std_logic_vector(7 downto 0);
    signal call68_419 : std_logic_vector(7 downto 0);
    signal call73_432 : std_logic_vector(7 downto 0);
    signal call_219 : std_logic_vector(7 downto 0);
    signal cmp169384_512 : std_logic_vector(0 downto 0);
    signal cmp303381_1067 : std_logic_vector(0 downto 0);
    signal cmp388_497 : std_logic_vector(0 downto 0);
    signal conv119_578 : std_logic_vector(63 downto 0);
    signal conv11_261 : std_logic_vector(31 downto 0);
    signal conv124_591 : std_logic_vector(63 downto 0);
    signal conv130_609 : std_logic_vector(63 downto 0);
    signal conv136_627 : std_logic_vector(63 downto 0);
    signal conv142_645 : std_logic_vector(63 downto 0);
    signal conv148_663 : std_logic_vector(63 downto 0);
    signal conv154_681 : std_logic_vector(63 downto 0);
    signal conv160_699 : std_logic_vector(63 downto 0);
    signal conv175_785 : std_logic_vector(63 downto 0);
    signal conv17_273 : std_logic_vector(15 downto 0);
    signal conv180_798 : std_logic_vector(63 downto 0);
    signal conv186_816 : std_logic_vector(63 downto 0);
    signal conv192_834 : std_logic_vector(63 downto 0);
    signal conv198_852 : std_logic_vector(63 downto 0);
    signal conv1_223 : std_logic_vector(31 downto 0);
    signal conv204_870 : std_logic_vector(63 downto 0);
    signal conv20_286 : std_logic_vector(15 downto 0);
    signal conv210_888 : std_logic_vector(63 downto 0);
    signal conv216_906 : std_logic_vector(63 downto 0);
    signal conv227_944 : std_logic_vector(63 downto 0);
    signal conv233_957 : std_logic_vector(63 downto 0);
    signal conv239_966 : std_logic_vector(7 downto 0);
    signal conv245_976 : std_logic_vector(7 downto 0);
    signal conv251_986 : std_logic_vector(7 downto 0);
    signal conv257_996 : std_logic_vector(7 downto 0);
    signal conv263_1006 : std_logic_vector(7 downto 0);
    signal conv269_1016 : std_logic_vector(7 downto 0);
    signal conv26_298 : std_logic_vector(31 downto 0);
    signal conv275_1026 : std_logic_vector(7 downto 0);
    signal conv281_1036 : std_logic_vector(7 downto 0);
    signal conv29_311 : std_logic_vector(31 downto 0);
    signal conv314_1130 : std_logic_vector(7 downto 0);
    signal conv320_1140 : std_logic_vector(7 downto 0);
    signal conv326_1150 : std_logic_vector(7 downto 0);
    signal conv332_1160 : std_logic_vector(7 downto 0);
    signal conv338_1170 : std_logic_vector(7 downto 0);
    signal conv344_1180 : std_logic_vector(7 downto 0);
    signal conv350_1190 : std_logic_vector(7 downto 0);
    signal conv356_1200 : std_logic_vector(7 downto 0);
    signal conv35_323 : std_logic_vector(31 downto 0);
    signal conv38_336 : std_logic_vector(31 downto 0);
    signal conv3_236 : std_logic_vector(31 downto 0);
    signal conv44_348 : std_logic_vector(15 downto 0);
    signal conv47_361 : std_logic_vector(15 downto 0);
    signal conv53_373 : std_logic_vector(31 downto 0);
    signal conv56_386 : std_logic_vector(31 downto 0);
    signal conv62_398 : std_logic_vector(31 downto 0);
    signal conv65_411 : std_logic_vector(31 downto 0);
    signal conv71_423 : std_logic_vector(31 downto 0);
    signal conv74_436 : std_logic_vector(31 downto 0);
    signal conv84_445 : std_logic_vector(31 downto 0);
    signal conv8_248 : std_logic_vector(31 downto 0);
    signal conv93_459 : std_logic_vector(31 downto 0);
    signal exitcond17_719 : std_logic_vector(0 downto 0);
    signal exitcond5_1235 : std_logic_vector(0 downto 0);
    signal exitcond_926 : std_logic_vector(0 downto 0);
    signal inc223_921 : std_logic_vector(31 downto 0);
    signal inc376_1230 : std_logic_vector(31 downto 0);
    signal inc_714 : std_logic_vector(31 downto 0);
    signal ix_x0389_555 : std_logic_vector(31 downto 0);
    signal ix_x1385_762 : std_logic_vector(31 downto 0);
    signal ix_x2382_1106 : std_logic_vector(31 downto 0);
    signal mul100_474 : std_logic_vector(31 downto 0);
    signal mul103_479 : std_logic_vector(31 downto 0);
    signal mul85_455 : std_logic_vector(31 downto 0);
    signal mul91_464 : std_logic_vector(31 downto 0);
    signal mul94_469 : std_logic_vector(31 downto 0);
    signal mul_450 : std_logic_vector(31 downto 0);
    signal ptr_deref_1125_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1125_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1125_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1125_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1125_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_706_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_706_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_706_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_706_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_706_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_706_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_913_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_913_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_913_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_913_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_913_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_913_word_offset_0 : std_logic_vector(15 downto 0);
    signal shl121_584 : std_logic_vector(63 downto 0);
    signal shl127_602 : std_logic_vector(63 downto 0);
    signal shl133_620 : std_logic_vector(63 downto 0);
    signal shl139_638 : std_logic_vector(63 downto 0);
    signal shl145_656 : std_logic_vector(63 downto 0);
    signal shl151_674 : std_logic_vector(63 downto 0);
    signal shl157_692 : std_logic_vector(63 downto 0);
    signal shl177_791 : std_logic_vector(63 downto 0);
    signal shl183_809 : std_logic_vector(63 downto 0);
    signal shl189_827 : std_logic_vector(63 downto 0);
    signal shl18_279 : std_logic_vector(15 downto 0);
    signal shl195_845 : std_logic_vector(63 downto 0);
    signal shl201_863 : std_logic_vector(63 downto 0);
    signal shl207_881 : std_logic_vector(63 downto 0);
    signal shl213_899 : std_logic_vector(63 downto 0);
    signal shl27_304 : std_logic_vector(31 downto 0);
    signal shl36_329 : std_logic_vector(31 downto 0);
    signal shl45_354 : std_logic_vector(15 downto 0);
    signal shl54_379 : std_logic_vector(31 downto 0);
    signal shl63_404 : std_logic_vector(31 downto 0);
    signal shl72_429 : std_logic_vector(31 downto 0);
    signal shl9_254 : std_logic_vector(31 downto 0);
    signal shl_229 : std_logic_vector(31 downto 0);
    signal shr111379_491 : std_logic_vector(15 downto 0);
    signal shr242_972 : std_logic_vector(63 downto 0);
    signal shr248_982 : std_logic_vector(63 downto 0);
    signal shr254_992 : std_logic_vector(63 downto 0);
    signal shr260_1002 : std_logic_vector(63 downto 0);
    signal shr266_1012 : std_logic_vector(63 downto 0);
    signal shr272_1022 : std_logic_vector(63 downto 0);
    signal shr278_1032 : std_logic_vector(63 downto 0);
    signal shr317_1136 : std_logic_vector(63 downto 0);
    signal shr323_1146 : std_logic_vector(63 downto 0);
    signal shr329_1156 : std_logic_vector(63 downto 0);
    signal shr335_1166 : std_logic_vector(63 downto 0);
    signal shr341_1176 : std_logic_vector(63 downto 0);
    signal shr347_1186 : std_logic_vector(63 downto 0);
    signal shr353_1196 : std_logic_vector(63 downto 0);
    signal shr378_485 : std_logic_vector(15 downto 0);
    signal sub_962 : std_logic_vector(63 downto 0);
    signal tmp10_752 : std_logic_vector(0 downto 0);
    signal tmp11_524 : std_logic_vector(31 downto 0);
    signal tmp12_528 : std_logic_vector(31 downto 0);
    signal tmp13_533 : std_logic_vector(31 downto 0);
    signal tmp14_539 : std_logic_vector(31 downto 0);
    signal tmp15_545 : std_logic_vector(0 downto 0);
    signal tmp1_1084 : std_logic_vector(31 downto 0);
    signal tmp2_1090 : std_logic_vector(31 downto 0);
    signal tmp310_1126 : std_logic_vector(63 downto 0);
    signal tmp3_1096 : std_logic_vector(0 downto 0);
    signal tmp6_731 : std_logic_vector(31 downto 0);
    signal tmp7_735 : std_logic_vector(31 downto 0);
    signal tmp8_740 : std_logic_vector(31 downto 0);
    signal tmp9_746 : std_logic_vector(31 downto 0);
    signal tmp_1079 : std_logic_vector(31 downto 0);
    signal type_cast_1000_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1010_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1020_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1030_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1065_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1088_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1094_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1101_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1110_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1112_wire : std_logic_vector(31 downto 0);
    signal type_cast_1134_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1144_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1154_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1164_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1174_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1184_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1194_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1228_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_227_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_252_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_277_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_302_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_327_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_352_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_377_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_402_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_427_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_483_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_489_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_495_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_510_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_537_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_543_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_550_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_559_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_561_wire : std_logic_vector(31 downto 0);
    signal type_cast_582_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_600_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_618_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_636_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_654_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_672_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_690_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_712_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_744_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_750_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_757_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_766_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_768_wire : std_logic_vector(31 downto 0);
    signal type_cast_789_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_807_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_825_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_843_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_861_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_879_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_897_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_919_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_942_wire : std_logic_vector(63 downto 0);
    signal type_cast_955_wire : std_logic_vector(63 downto 0);
    signal type_cast_970_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_980_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_990_wire_constant : std_logic_vector(63 downto 0);
    signal umax16_552 : std_logic_vector(31 downto 0);
    signal umax4_1103 : std_logic_vector(31 downto 0);
    signal umax_759 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    array_obj_ref_1120_constant_part_of_offset <= "1000000000000000";
    array_obj_ref_1120_offset_scale_factor_0 <= "0100000000000000";
    array_obj_ref_1120_offset_scale_factor_1 <= "0100000000000000";
    array_obj_ref_1120_offset_scale_factor_2 <= "0000000000000001";
    array_obj_ref_1120_resized_base_address <= "0000000000000000";
    array_obj_ref_569_constant_part_of_offset <= "0000000000000000";
    array_obj_ref_569_offset_scale_factor_0 <= "0100000000000000";
    array_obj_ref_569_offset_scale_factor_1 <= "0100000000000000";
    array_obj_ref_569_offset_scale_factor_2 <= "0000000000000001";
    array_obj_ref_569_resized_base_address <= "0000000000000000";
    array_obj_ref_776_constant_part_of_offset <= "0100000000000000";
    array_obj_ref_776_offset_scale_factor_0 <= "0100000000000000";
    array_obj_ref_776_offset_scale_factor_1 <= "0100000000000000";
    array_obj_ref_776_offset_scale_factor_2 <= "0000000000000001";
    array_obj_ref_776_resized_base_address <= "0000000000000000";
    ptr_deref_1125_word_offset_0 <= "0000000000000000";
    ptr_deref_706_word_offset_0 <= "0000000000000000";
    ptr_deref_913_word_offset_0 <= "0000000000000000";
    type_cast_1000_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1010_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1020_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1030_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1065_wire_constant <= "00000000000000000000000000000111";
    type_cast_1088_wire_constant <= "00000000000000000000000000000011";
    type_cast_1094_wire_constant <= "00000000000000000000000000000001";
    type_cast_1101_wire_constant <= "00000000000000000000000000000001";
    type_cast_1110_wire_constant <= "00000000000000000000000000000000";
    type_cast_1134_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1144_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1154_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1164_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1174_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1184_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1194_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1228_wire_constant <= "00000000000000000000000000000001";
    type_cast_227_wire_constant <= "00000000000000000000000000001000";
    type_cast_252_wire_constant <= "00000000000000000000000000001000";
    type_cast_277_wire_constant <= "0000000000001000";
    type_cast_302_wire_constant <= "00000000000000000000000000001000";
    type_cast_327_wire_constant <= "00000000000000000000000000001000";
    type_cast_352_wire_constant <= "0000000000001000";
    type_cast_377_wire_constant <= "00000000000000000000000000001000";
    type_cast_402_wire_constant <= "00000000000000000000000000001000";
    type_cast_427_wire_constant <= "00000000000000000000000000001000";
    type_cast_483_wire_constant <= "0000000000000011";
    type_cast_489_wire_constant <= "0000000000000011";
    type_cast_495_wire_constant <= "00000000000000000000000000000111";
    type_cast_510_wire_constant <= "00000000000000000000000000000111";
    type_cast_537_wire_constant <= "00000000000000000000000000000011";
    type_cast_543_wire_constant <= "00000000000000000000000000000001";
    type_cast_550_wire_constant <= "00000000000000000000000000000001";
    type_cast_559_wire_constant <= "00000000000000000000000000000000";
    type_cast_582_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_600_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_618_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_636_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_654_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_672_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_690_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_712_wire_constant <= "00000000000000000000000000000001";
    type_cast_744_wire_constant <= "00000000000000000000000000000011";
    type_cast_750_wire_constant <= "00000000000000000000000000000001";
    type_cast_757_wire_constant <= "00000000000000000000000000000001";
    type_cast_766_wire_constant <= "00000000000000000000000000000000";
    type_cast_789_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_807_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_825_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_843_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_861_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_879_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_897_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_919_wire_constant <= "00000000000000000000000000000001";
    type_cast_970_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_980_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_990_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    phi_stmt_1106: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1110_wire_constant & type_cast_1112_wire;
      req <= phi_stmt_1106_req_0 & phi_stmt_1106_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1106",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1106_ack_0,
          idata => idata,
          odata => ix_x2382_1106,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1106
    phi_stmt_555: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_559_wire_constant & type_cast_561_wire;
      req <= phi_stmt_555_req_0 & phi_stmt_555_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_555",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_555_ack_0,
          idata => idata,
          odata => ix_x0389_555,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_555
    phi_stmt_762: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_766_wire_constant & type_cast_768_wire;
      req <= phi_stmt_762_req_0 & phi_stmt_762_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_762",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_762_ack_0,
          idata => idata,
          odata => ix_x1385_762,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_762
    -- flow-through select operator MUX_1102_inst
    umax4_1103 <= tmp2_1090 when (tmp3_1096(0) /=  '0') else type_cast_1101_wire_constant;
    -- flow-through select operator MUX_551_inst
    umax16_552 <= tmp14_539 when (tmp15_545(0) /=  '0') else type_cast_550_wire_constant;
    -- flow-through select operator MUX_758_inst
    umax_759 <= tmp9_746 when (tmp10_752(0) /=  '0') else type_cast_757_wire_constant;
    addr_of_1121_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1121_final_reg_req_0;
      addr_of_1121_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1121_final_reg_req_1;
      addr_of_1121_final_reg_ack_1<= rack(0);
      addr_of_1121_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1121_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1120_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx309_1122,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_570_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_570_final_reg_req_0;
      addr_of_570_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_570_final_reg_req_1;
      addr_of_570_final_reg_ack_1<= rack(0);
      addr_of_570_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_570_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_569_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_571,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_777_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_777_final_reg_req_0;
      addr_of_777_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_777_final_reg_req_1;
      addr_of_777_final_reg_ack_1<= rack(0);
      addr_of_777_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_777_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_776_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx220_778,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1005_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1005_inst_req_0;
      type_cast_1005_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1005_inst_req_1;
      type_cast_1005_inst_ack_1<= rack(0);
      type_cast_1005_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1005_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr260_1002,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv263_1006,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1015_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1015_inst_req_0;
      type_cast_1015_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1015_inst_req_1;
      type_cast_1015_inst_ack_1<= rack(0);
      type_cast_1015_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1015_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr266_1012,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv269_1016,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1025_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1025_inst_req_0;
      type_cast_1025_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1025_inst_req_1;
      type_cast_1025_inst_ack_1<= rack(0);
      type_cast_1025_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1025_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr272_1022,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv275_1026,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1035_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1035_inst_req_0;
      type_cast_1035_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1035_inst_req_1;
      type_cast_1035_inst_ack_1<= rack(0);
      type_cast_1035_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1035_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr278_1032,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv281_1036,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1112_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1112_inst_req_0;
      type_cast_1112_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1112_inst_req_1;
      type_cast_1112_inst_ack_1<= rack(0);
      type_cast_1112_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1112_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc376_1230,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1112_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1129_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1129_inst_req_0;
      type_cast_1129_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1129_inst_req_1;
      type_cast_1129_inst_ack_1<= rack(0);
      type_cast_1129_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1129_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp310_1126,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv314_1130,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1139_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1139_inst_req_0;
      type_cast_1139_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1139_inst_req_1;
      type_cast_1139_inst_ack_1<= rack(0);
      type_cast_1139_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1139_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr317_1136,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv320_1140,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1149_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1149_inst_req_0;
      type_cast_1149_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1149_inst_req_1;
      type_cast_1149_inst_ack_1<= rack(0);
      type_cast_1149_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1149_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr323_1146,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv326_1150,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1159_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1159_inst_req_0;
      type_cast_1159_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1159_inst_req_1;
      type_cast_1159_inst_ack_1<= rack(0);
      type_cast_1159_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1159_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr329_1156,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv332_1160,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1169_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1169_inst_req_0;
      type_cast_1169_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1169_inst_req_1;
      type_cast_1169_inst_ack_1<= rack(0);
      type_cast_1169_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1169_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr335_1166,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv338_1170,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1179_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1179_inst_req_0;
      type_cast_1179_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1179_inst_req_1;
      type_cast_1179_inst_ack_1<= rack(0);
      type_cast_1179_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1179_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr341_1176,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv344_1180,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1189_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1189_inst_req_0;
      type_cast_1189_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1189_inst_req_1;
      type_cast_1189_inst_ack_1<= rack(0);
      type_cast_1189_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1189_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr347_1186,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv350_1190,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1199_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1199_inst_req_0;
      type_cast_1199_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1199_inst_req_1;
      type_cast_1199_inst_ack_1<= rack(0);
      type_cast_1199_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1199_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr353_1196,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv356_1200,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_222_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_222_inst_req_0;
      type_cast_222_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_222_inst_req_1;
      type_cast_222_inst_ack_1<= rack(0);
      type_cast_222_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_222_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_219,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1_223,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_235_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_235_inst_req_0;
      type_cast_235_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_235_inst_req_1;
      type_cast_235_inst_ack_1<= rack(0);
      type_cast_235_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_235_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_232,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv3_236,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_247_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_247_inst_req_0;
      type_cast_247_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_247_inst_req_1;
      type_cast_247_inst_ack_1<= rack(0);
      type_cast_247_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_247_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call5_244,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv8_248,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_260_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_260_inst_req_0;
      type_cast_260_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_260_inst_req_1;
      type_cast_260_inst_ack_1<= rack(0);
      type_cast_260_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_260_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call10_257,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv11_261,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_272_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_272_inst_req_0;
      type_cast_272_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_272_inst_req_1;
      type_cast_272_inst_ack_1<= rack(0);
      type_cast_272_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_272_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call14_269,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_273,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_285_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_285_inst_req_0;
      type_cast_285_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_285_inst_req_1;
      type_cast_285_inst_ack_1<= rack(0);
      type_cast_285_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_285_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call19_282,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv20_286,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_297_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_297_inst_req_0;
      type_cast_297_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_297_inst_req_1;
      type_cast_297_inst_ack_1<= rack(0);
      type_cast_297_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_297_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call23_294,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv26_298,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_310_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_310_inst_req_0;
      type_cast_310_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_310_inst_req_1;
      type_cast_310_inst_ack_1<= rack(0);
      type_cast_310_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_310_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call28_307,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv29_311,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_322_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_322_inst_req_0;
      type_cast_322_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_322_inst_req_1;
      type_cast_322_inst_ack_1<= rack(0);
      type_cast_322_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_322_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call32_319,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv35_323,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_335_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_335_inst_req_0;
      type_cast_335_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_335_inst_req_1;
      type_cast_335_inst_ack_1<= rack(0);
      type_cast_335_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_335_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call37_332,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv38_336,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_347_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_347_inst_req_0;
      type_cast_347_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_347_inst_req_1;
      type_cast_347_inst_ack_1<= rack(0);
      type_cast_347_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_347_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call41_344,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv44_348,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_360_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_360_inst_req_0;
      type_cast_360_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_360_inst_req_1;
      type_cast_360_inst_ack_1<= rack(0);
      type_cast_360_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_360_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call46_357,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv47_361,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_372_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_372_inst_req_0;
      type_cast_372_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_372_inst_req_1;
      type_cast_372_inst_ack_1<= rack(0);
      type_cast_372_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_372_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call50_369,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv53_373,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_385_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_385_inst_req_0;
      type_cast_385_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_385_inst_req_1;
      type_cast_385_inst_ack_1<= rack(0);
      type_cast_385_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_385_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call55_382,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv56_386,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_397_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_397_inst_req_0;
      type_cast_397_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_397_inst_req_1;
      type_cast_397_inst_ack_1<= rack(0);
      type_cast_397_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_397_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call59_394,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv62_398,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_410_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_410_inst_req_0;
      type_cast_410_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_410_inst_req_1;
      type_cast_410_inst_ack_1<= rack(0);
      type_cast_410_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_410_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call64_407,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv65_411,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_422_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_422_inst_req_0;
      type_cast_422_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_422_inst_req_1;
      type_cast_422_inst_ack_1<= rack(0);
      type_cast_422_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_422_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call68_419,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv71_423,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_435_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_435_inst_req_0;
      type_cast_435_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_435_inst_req_1;
      type_cast_435_inst_ack_1<= rack(0);
      type_cast_435_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_435_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call73_432,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv74_436,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_444_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_444_inst_req_0;
      type_cast_444_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_444_inst_req_1;
      type_cast_444_inst_ack_1<= rack(0);
      type_cast_444_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_444_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add21_291,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv84_445,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_458_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_458_inst_req_0;
      type_cast_458_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_458_inst_req_1;
      type_cast_458_inst_ack_1<= rack(0);
      type_cast_458_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_458_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add48_366,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv93_459,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_527_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_527_inst_req_0;
      type_cast_527_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_527_inst_req_1;
      type_cast_527_inst_ack_1<= rack(0);
      type_cast_527_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_527_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add21_291,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp12_528,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_561_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_561_inst_req_0;
      type_cast_561_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_561_inst_req_1;
      type_cast_561_inst_ack_1<= rack(0);
      type_cast_561_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_561_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc_714,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_561_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_577_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_577_inst_req_0;
      type_cast_577_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_577_inst_req_1;
      type_cast_577_inst_ack_1<= rack(0);
      type_cast_577_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_577_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call118_574,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv119_578,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_590_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_590_inst_req_0;
      type_cast_590_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_590_inst_req_1;
      type_cast_590_inst_ack_1<= rack(0);
      type_cast_590_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_590_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call122_587,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv124_591,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_608_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_608_inst_req_0;
      type_cast_608_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_608_inst_req_1;
      type_cast_608_inst_ack_1<= rack(0);
      type_cast_608_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_608_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call128_605,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv130_609,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_626_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_626_inst_req_0;
      type_cast_626_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_626_inst_req_1;
      type_cast_626_inst_ack_1<= rack(0);
      type_cast_626_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_626_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call134_623,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv136_627,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_644_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_644_inst_req_0;
      type_cast_644_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_644_inst_req_1;
      type_cast_644_inst_ack_1<= rack(0);
      type_cast_644_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_644_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call140_641,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv142_645,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_662_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_662_inst_req_0;
      type_cast_662_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_662_inst_req_1;
      type_cast_662_inst_ack_1<= rack(0);
      type_cast_662_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_662_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call146_659,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv148_663,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_680_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_680_inst_req_0;
      type_cast_680_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_680_inst_req_1;
      type_cast_680_inst_ack_1<= rack(0);
      type_cast_680_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_680_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call152_677,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv154_681,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_698_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_698_inst_req_0;
      type_cast_698_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_698_inst_req_1;
      type_cast_698_inst_ack_1<= rack(0);
      type_cast_698_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_698_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call158_695,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv160_699,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_734_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_734_inst_req_0;
      type_cast_734_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_734_inst_req_1;
      type_cast_734_inst_ack_1<= rack(0);
      type_cast_734_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_734_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add48_366,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp7_735,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_768_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_768_inst_req_0;
      type_cast_768_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_768_inst_req_1;
      type_cast_768_inst_ack_1<= rack(0);
      type_cast_768_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_768_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc223_921,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_768_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_784_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_784_inst_req_0;
      type_cast_784_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_784_inst_req_1;
      type_cast_784_inst_ack_1<= rack(0);
      type_cast_784_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_784_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call174_781,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv175_785,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_797_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_797_inst_req_0;
      type_cast_797_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_797_inst_req_1;
      type_cast_797_inst_ack_1<= rack(0);
      type_cast_797_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_797_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call178_794,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv180_798,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_815_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_815_inst_req_0;
      type_cast_815_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_815_inst_req_1;
      type_cast_815_inst_ack_1<= rack(0);
      type_cast_815_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_815_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call184_812,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv186_816,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_833_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_833_inst_req_0;
      type_cast_833_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_833_inst_req_1;
      type_cast_833_inst_ack_1<= rack(0);
      type_cast_833_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_833_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call190_830,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv192_834,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_851_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_851_inst_req_0;
      type_cast_851_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_851_inst_req_1;
      type_cast_851_inst_ack_1<= rack(0);
      type_cast_851_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_851_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call196_848,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv198_852,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_869_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_869_inst_req_0;
      type_cast_869_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_869_inst_req_1;
      type_cast_869_inst_ack_1<= rack(0);
      type_cast_869_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_869_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call202_866,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv204_870,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_887_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_887_inst_req_0;
      type_cast_887_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_887_inst_req_1;
      type_cast_887_inst_ack_1<= rack(0);
      type_cast_887_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_887_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call208_884,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv210_888,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_905_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_905_inst_req_0;
      type_cast_905_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_905_inst_req_1;
      type_cast_905_inst_ack_1<= rack(0);
      type_cast_905_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_905_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call214_902,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv216_906,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_943_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_943_inst_req_0;
      type_cast_943_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_943_inst_req_1;
      type_cast_943_inst_ack_1<= rack(0);
      type_cast_943_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_943_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_942_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv227_944,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_956_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_956_inst_req_0;
      type_cast_956_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_956_inst_req_1;
      type_cast_956_inst_ack_1<= rack(0);
      type_cast_956_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_956_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_955_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv233_957,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_965_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_965_inst_req_0;
      type_cast_965_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_965_inst_req_1;
      type_cast_965_inst_ack_1<= rack(0);
      type_cast_965_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_965_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub_962,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv239_966,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_975_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_975_inst_req_0;
      type_cast_975_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_975_inst_req_1;
      type_cast_975_inst_ack_1<= rack(0);
      type_cast_975_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_975_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr242_972,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv245_976,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_985_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_985_inst_req_0;
      type_cast_985_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_985_inst_req_1;
      type_cast_985_inst_ack_1<= rack(0);
      type_cast_985_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_985_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr248_982,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv251_986,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_995_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_995_inst_req_0;
      type_cast_995_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_995_inst_req_1;
      type_cast_995_inst_ack_1<= rack(0);
      type_cast_995_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_995_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr254_992,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv257_996,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1120_index_2_rename
    process(R_ix_x2382_1119_resized) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_ix_x2382_1119_resized;
      ov(15 downto 0) := iv;
      R_ix_x2382_1119_scaled <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1120_index_2_resize
    process(ix_x2382_1106) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ix_x2382_1106;
      ov := iv(15 downto 0);
      R_ix_x2382_1119_resized <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1120_root_address_inst
    process(array_obj_ref_1120_final_offset) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1120_final_offset;
      ov(15 downto 0) := iv;
      array_obj_ref_1120_root_address <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_569_index_2_rename
    process(R_ix_x0389_568_resized) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_ix_x0389_568_resized;
      ov(15 downto 0) := iv;
      R_ix_x0389_568_scaled <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_569_index_2_resize
    process(ix_x0389_555) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ix_x0389_555;
      ov := iv(15 downto 0);
      R_ix_x0389_568_resized <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_569_root_address_inst
    process(array_obj_ref_569_final_offset) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_569_final_offset;
      ov(15 downto 0) := iv;
      array_obj_ref_569_root_address <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_776_index_2_rename
    process(R_ix_x1385_775_resized) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_ix_x1385_775_resized;
      ov(15 downto 0) := iv;
      R_ix_x1385_775_scaled <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_776_index_2_resize
    process(ix_x1385_762) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ix_x1385_762;
      ov := iv(15 downto 0);
      R_ix_x1385_775_resized <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_776_root_address_inst
    process(array_obj_ref_776_final_offset) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_776_final_offset;
      ov(15 downto 0) := iv;
      array_obj_ref_776_root_address <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1125_addr_0
    process(ptr_deref_1125_root_address) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1125_root_address;
      ov(15 downto 0) := iv;
      ptr_deref_1125_word_address_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1125_base_resize
    process(arrayidx309_1122) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx309_1122;
      ov := iv(15 downto 0);
      ptr_deref_1125_resized_base_address <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1125_gather_scatter
    process(ptr_deref_1125_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1125_data_0;
      ov(63 downto 0) := iv;
      tmp310_1126 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1125_root_address_inst
    process(ptr_deref_1125_resized_base_address) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1125_resized_base_address;
      ov(15 downto 0) := iv;
      ptr_deref_1125_root_address <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_706_addr_0
    process(ptr_deref_706_root_address) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_706_root_address;
      ov(15 downto 0) := iv;
      ptr_deref_706_word_address_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_706_base_resize
    process(arrayidx_571) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_571;
      ov := iv(15 downto 0);
      ptr_deref_706_resized_base_address <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_706_gather_scatter
    process(add161_704) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add161_704;
      ov(63 downto 0) := iv;
      ptr_deref_706_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_706_root_address_inst
    process(ptr_deref_706_resized_base_address) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_706_resized_base_address;
      ov(15 downto 0) := iv;
      ptr_deref_706_root_address <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_913_addr_0
    process(ptr_deref_913_root_address) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_913_root_address;
      ov(15 downto 0) := iv;
      ptr_deref_913_word_address_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_913_base_resize
    process(arrayidx220_778) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx220_778;
      ov := iv(15 downto 0);
      ptr_deref_913_resized_base_address <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_913_gather_scatter
    process(add217_911) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add217_911;
      ov(63 downto 0) := iv;
      ptr_deref_913_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_913_root_address_inst
    process(ptr_deref_913_resized_base_address) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_913_resized_base_address;
      ov(15 downto 0) := iv;
      ptr_deref_913_root_address <= ov(15 downto 0);
      --
    end process;
    if_stmt_1068_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp303381_1067;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1068_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1068_branch_req_0,
          ack0 => if_stmt_1068_branch_ack_0,
          ack1 => if_stmt_1068_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1236_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond5_1235;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1236_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1236_branch_req_0,
          ack0 => if_stmt_1236_branch_ack_0,
          ack1 => if_stmt_1236_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_498_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp388_497;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_498_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_498_branch_req_0,
          ack0 => if_stmt_498_branch_ack_0,
          ack1 => if_stmt_498_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_513_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp169384_512;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_513_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_513_branch_req_0,
          ack0 => if_stmt_513_branch_ack_0,
          ack1 => if_stmt_513_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_720_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond17_719;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_720_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_720_branch_req_0,
          ack0 => if_stmt_720_branch_ack_0,
          ack1 => if_stmt_720_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_927_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond_926;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_927_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_927_branch_req_0,
          ack0 => if_stmt_927_branch_ack_0,
          ack1 => if_stmt_927_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u32_u32_1229_inst
    process(ix_x2382_1106) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(ix_x2382_1106, type_cast_1228_wire_constant, tmp_var);
      inc376_1230 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_713_inst
    process(ix_x0389_555) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(ix_x0389_555, type_cast_712_wire_constant, tmp_var);
      inc_714 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_920_inst
    process(ix_x1385_762) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(ix_x1385_762, type_cast_919_wire_constant, tmp_var);
      inc223_921 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1234_inst
    process(inc376_1230, umax4_1103) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc376_1230, umax4_1103, tmp_var);
      exitcond5_1235 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_718_inst
    process(inc_714, umax16_552) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc_714, umax16_552, tmp_var);
      exitcond17_719 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_925_inst
    process(inc223_921, umax_759) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc223_921, umax_759, tmp_var);
      exitcond_926 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_484_inst
    process(add21_291) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add21_291, type_cast_483_wire_constant, tmp_var);
      shr378_485 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_490_inst
    process(add48_366) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add48_366, type_cast_489_wire_constant, tmp_var);
      shr111379_491 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1089_inst
    process(tmp1_1084) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp1_1084, type_cast_1088_wire_constant, tmp_var);
      tmp2_1090 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_538_inst
    process(tmp13_533) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp13_533, type_cast_537_wire_constant, tmp_var);
      tmp14_539 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_745_inst
    process(tmp8_740) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp8_740, type_cast_744_wire_constant, tmp_var);
      tmp9_746 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1001_inst
    process(sub_962) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_962, type_cast_1000_wire_constant, tmp_var);
      shr260_1002 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1011_inst
    process(sub_962) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_962, type_cast_1010_wire_constant, tmp_var);
      shr266_1012 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1021_inst
    process(sub_962) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_962, type_cast_1020_wire_constant, tmp_var);
      shr272_1022 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1031_inst
    process(sub_962) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_962, type_cast_1030_wire_constant, tmp_var);
      shr278_1032 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1135_inst
    process(tmp310_1126) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp310_1126, type_cast_1134_wire_constant, tmp_var);
      shr317_1136 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1145_inst
    process(tmp310_1126) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp310_1126, type_cast_1144_wire_constant, tmp_var);
      shr323_1146 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1155_inst
    process(tmp310_1126) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp310_1126, type_cast_1154_wire_constant, tmp_var);
      shr329_1156 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1165_inst
    process(tmp310_1126) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp310_1126, type_cast_1164_wire_constant, tmp_var);
      shr335_1166 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1175_inst
    process(tmp310_1126) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp310_1126, type_cast_1174_wire_constant, tmp_var);
      shr341_1176 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1185_inst
    process(tmp310_1126) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp310_1126, type_cast_1184_wire_constant, tmp_var);
      shr347_1186 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1195_inst
    process(tmp310_1126) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp310_1126, type_cast_1194_wire_constant, tmp_var);
      shr353_1196 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_971_inst
    process(sub_962) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_962, type_cast_970_wire_constant, tmp_var);
      shr242_972 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_981_inst
    process(sub_962) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_962, type_cast_980_wire_constant, tmp_var);
      shr248_982 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_991_inst
    process(sub_962) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_962, type_cast_990_wire_constant, tmp_var);
      shr254_992 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1078_inst
    process(add66_416, add57_391) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add66_416, add57_391, tmp_var);
      tmp_1079 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1083_inst
    process(tmp_1079, add75_441) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp_1079, add75_441, tmp_var);
      tmp1_1084 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_449_inst
    process(add12_266, add_241) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add12_266, add_241, tmp_var);
      mul_450 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_454_inst
    process(mul_450, conv84_445) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_450, conv84_445, tmp_var);
      mul85_455 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_463_inst
    process(add39_341, add30_316) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add39_341, add30_316, tmp_var);
      mul91_464 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_468_inst
    process(mul91_464, conv93_459) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul91_464, conv93_459, tmp_var);
      mul94_469 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_473_inst
    process(add66_416, add57_391) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add66_416, add57_391, tmp_var);
      mul100_474 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_478_inst
    process(mul100_474, add75_441) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul100_474, add75_441, tmp_var);
      mul103_479 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_523_inst
    process(add12_266, add_241) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add12_266, add_241, tmp_var);
      tmp11_524 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_532_inst
    process(tmp11_524, tmp12_528) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp11_524, tmp12_528, tmp_var);
      tmp13_533 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_730_inst
    process(add39_341, add30_316) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add39_341, add30_316, tmp_var);
      tmp6_731 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_739_inst
    process(tmp6_731, tmp7_735) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp6_731, tmp7_735, tmp_var);
      tmp8_740 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_290_inst
    process(shl18_279, conv20_286) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl18_279, conv20_286, tmp_var);
      add21_291 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_365_inst
    process(shl45_354, conv47_361) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl45_354, conv47_361, tmp_var);
      add48_366 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_240_inst
    process(shl_229, conv3_236) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_229, conv3_236, tmp_var);
      add_241 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_265_inst
    process(shl9_254, conv11_261) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl9_254, conv11_261, tmp_var);
      add12_266 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_315_inst
    process(shl27_304, conv29_311) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl27_304, conv29_311, tmp_var);
      add30_316 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_340_inst
    process(shl36_329, conv38_336) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl36_329, conv38_336, tmp_var);
      add39_341 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_390_inst
    process(shl54_379, conv56_386) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl54_379, conv56_386, tmp_var);
      add57_391 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_415_inst
    process(shl63_404, conv65_411) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl63_404, conv65_411, tmp_var);
      add66_416 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_440_inst
    process(shl72_429, conv74_436) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl72_429, conv74_436, tmp_var);
      add75_441 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_595_inst
    process(shl121_584, conv124_591) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl121_584, conv124_591, tmp_var);
      add125_596 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_613_inst
    process(shl127_602, conv130_609) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl127_602, conv130_609, tmp_var);
      add131_614 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_631_inst
    process(shl133_620, conv136_627) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl133_620, conv136_627, tmp_var);
      add137_632 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_649_inst
    process(shl139_638, conv142_645) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl139_638, conv142_645, tmp_var);
      add143_650 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_667_inst
    process(shl145_656, conv148_663) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl145_656, conv148_663, tmp_var);
      add149_668 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_685_inst
    process(shl151_674, conv154_681) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl151_674, conv154_681, tmp_var);
      add155_686 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_703_inst
    process(shl157_692, conv160_699) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl157_692, conv160_699, tmp_var);
      add161_704 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_802_inst
    process(shl177_791, conv180_798) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl177_791, conv180_798, tmp_var);
      add181_803 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_820_inst
    process(shl183_809, conv186_816) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl183_809, conv186_816, tmp_var);
      add187_821 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_838_inst
    process(shl189_827, conv192_834) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl189_827, conv192_834, tmp_var);
      add193_839 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_856_inst
    process(shl195_845, conv198_852) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl195_845, conv198_852, tmp_var);
      add199_857 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_874_inst
    process(shl201_863, conv204_870) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl201_863, conv204_870, tmp_var);
      add205_875 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_892_inst
    process(shl207_881, conv210_888) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl207_881, conv210_888, tmp_var);
      add211_893 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_910_inst
    process(shl213_899, conv216_906) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl213_899, conv216_906, tmp_var);
      add217_911 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_278_inst
    process(conv17_273) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv17_273, type_cast_277_wire_constant, tmp_var);
      shl18_279 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_353_inst
    process(conv44_348) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv44_348, type_cast_352_wire_constant, tmp_var);
      shl45_354 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_228_inst
    process(conv1_223) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv1_223, type_cast_227_wire_constant, tmp_var);
      shl_229 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_253_inst
    process(conv8_248) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv8_248, type_cast_252_wire_constant, tmp_var);
      shl9_254 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_303_inst
    process(conv26_298) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv26_298, type_cast_302_wire_constant, tmp_var);
      shl27_304 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_328_inst
    process(conv35_323) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv35_323, type_cast_327_wire_constant, tmp_var);
      shl36_329 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_378_inst
    process(conv53_373) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv53_373, type_cast_377_wire_constant, tmp_var);
      shl54_379 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_403_inst
    process(conv62_398) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv62_398, type_cast_402_wire_constant, tmp_var);
      shl63_404 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_428_inst
    process(conv71_423) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv71_423, type_cast_427_wire_constant, tmp_var);
      shl72_429 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_583_inst
    process(conv119_578) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv119_578, type_cast_582_wire_constant, tmp_var);
      shl121_584 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_601_inst
    process(add125_596) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add125_596, type_cast_600_wire_constant, tmp_var);
      shl127_602 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_619_inst
    process(add131_614) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add131_614, type_cast_618_wire_constant, tmp_var);
      shl133_620 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_637_inst
    process(add137_632) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add137_632, type_cast_636_wire_constant, tmp_var);
      shl139_638 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_655_inst
    process(add143_650) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add143_650, type_cast_654_wire_constant, tmp_var);
      shl145_656 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_673_inst
    process(add149_668) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add149_668, type_cast_672_wire_constant, tmp_var);
      shl151_674 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_691_inst
    process(add155_686) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add155_686, type_cast_690_wire_constant, tmp_var);
      shl157_692 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_790_inst
    process(conv175_785) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv175_785, type_cast_789_wire_constant, tmp_var);
      shl177_791 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_808_inst
    process(add181_803) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add181_803, type_cast_807_wire_constant, tmp_var);
      shl183_809 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_826_inst
    process(add187_821) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add187_821, type_cast_825_wire_constant, tmp_var);
      shl189_827 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_844_inst
    process(add193_839) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add193_839, type_cast_843_wire_constant, tmp_var);
      shl195_845 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_862_inst
    process(add199_857) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add199_857, type_cast_861_wire_constant, tmp_var);
      shl201_863 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_880_inst
    process(add205_875) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add205_875, type_cast_879_wire_constant, tmp_var);
      shl207_881 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_898_inst
    process(add211_893) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add211_893, type_cast_897_wire_constant, tmp_var);
      shl213_899 <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_961_inst
    process(conv233_957, conv227_944) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv233_957, conv227_944, tmp_var);
      sub_962 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1066_inst
    process(mul103_479) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul103_479, type_cast_1065_wire_constant, tmp_var);
      cmp303381_1067 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1095_inst
    process(tmp2_1090) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp2_1090, type_cast_1094_wire_constant, tmp_var);
      tmp3_1096 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_496_inst
    process(mul85_455) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul85_455, type_cast_495_wire_constant, tmp_var);
      cmp388_497 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_511_inst
    process(mul94_469) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul94_469, type_cast_510_wire_constant, tmp_var);
      cmp169384_512 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_544_inst
    process(tmp14_539) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp14_539, type_cast_543_wire_constant, tmp_var);
      tmp15_545 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_751_inst
    process(tmp9_746) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp9_746, type_cast_750_wire_constant, tmp_var);
      tmp10_752 <= tmp_var; --
    end process;
    -- shared split operator group (90) : array_obj_ref_1120_index_offset 
    ApIntAdd_group_90: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_ix_x2382_1119_scaled;
      array_obj_ref_1120_final_offset <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1120_index_offset_req_0;
      array_obj_ref_1120_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1120_index_offset_req_1;
      array_obj_ref_1120_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_90_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_90_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_90",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "1000000000000000",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 90
    -- shared split operator group (91) : array_obj_ref_569_index_offset 
    ApIntAdd_group_91: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_ix_x0389_568_scaled;
      array_obj_ref_569_final_offset <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_569_index_offset_req_0;
      array_obj_ref_569_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_569_index_offset_req_1;
      array_obj_ref_569_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_91_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_91_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_91",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 91
    -- shared split operator group (92) : array_obj_ref_776_index_offset 
    ApIntAdd_group_92: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_ix_x1385_775_scaled;
      array_obj_ref_776_final_offset <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_776_index_offset_req_0;
      array_obj_ref_776_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_776_index_offset_req_1;
      array_obj_ref_776_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_92_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_92_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_92",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0100000000000000",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 92
    -- unary operator type_cast_942_inst
    process(call226_938) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call226_938, tmp_var);
      type_cast_942_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_955_inst
    process(call232_952) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call232_952, tmp_var);
      type_cast_955_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : ptr_deref_1125_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1125_load_0_req_0;
      ptr_deref_1125_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1125_load_0_req_1;
      ptr_deref_1125_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1125_word_address_0;
      ptr_deref_1125_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 16,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(15 downto 0),
          mtag => memory_space_0_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_706_store_0 ptr_deref_913_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(31 downto 0);
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_706_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_913_store_0_req_0;
      ptr_deref_706_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_913_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_706_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_913_store_0_req_1;
      ptr_deref_706_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_913_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup0_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_706_word_address_0 & ptr_deref_913_word_address_0;
      data_in <= ptr_deref_706_data_0 & ptr_deref_913_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 16,
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(15 downto 0),
          mdata => memory_space_0_sr_data(63 downto 0),
          mtag => memory_space_0_sr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Concat_input_pipe_268_inst RPIPE_Concat_input_pipe_431_inst RPIPE_Concat_input_pipe_381_inst RPIPE_Concat_input_pipe_406_inst RPIPE_Concat_input_pipe_243_inst RPIPE_Concat_input_pipe_218_inst RPIPE_Concat_input_pipe_256_inst RPIPE_Concat_input_pipe_343_inst RPIPE_Concat_input_pipe_393_inst RPIPE_Concat_input_pipe_231_inst RPIPE_Concat_input_pipe_306_inst RPIPE_Concat_input_pipe_331_inst RPIPE_Concat_input_pipe_418_inst RPIPE_Concat_input_pipe_368_inst RPIPE_Concat_input_pipe_293_inst RPIPE_Concat_input_pipe_356_inst RPIPE_Concat_input_pipe_281_inst RPIPE_Concat_input_pipe_318_inst RPIPE_Concat_input_pipe_573_inst RPIPE_Concat_input_pipe_604_inst RPIPE_Concat_input_pipe_586_inst RPIPE_Concat_input_pipe_622_inst RPIPE_Concat_input_pipe_640_inst RPIPE_Concat_input_pipe_658_inst RPIPE_Concat_input_pipe_676_inst RPIPE_Concat_input_pipe_694_inst RPIPE_Concat_input_pipe_780_inst RPIPE_Concat_input_pipe_793_inst RPIPE_Concat_input_pipe_811_inst RPIPE_Concat_input_pipe_829_inst RPIPE_Concat_input_pipe_847_inst RPIPE_Concat_input_pipe_865_inst RPIPE_Concat_input_pipe_883_inst RPIPE_Concat_input_pipe_901_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(271 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 33 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 33 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 33 downto 0);
      signal guard_vector : std_logic_vector( 33 downto 0);
      constant outBUFs : IntegerArray(33 downto 0) := (33 => 1, 32 => 1, 31 => 1, 30 => 1, 29 => 1, 28 => 1, 27 => 1, 26 => 1, 25 => 1, 24 => 1, 23 => 1, 22 => 1, 21 => 1, 20 => 1, 19 => 1, 18 => 1, 17 => 1, 16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(33 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false, 17 => false, 18 => false, 19 => false, 20 => false, 21 => false, 22 => false, 23 => false, 24 => false, 25 => false, 26 => false, 27 => false, 28 => false, 29 => false, 30 => false, 31 => false, 32 => false, 33 => false);
      constant guardBuffering: IntegerArray(33 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2, 17 => 2, 18 => 2, 19 => 2, 20 => 2, 21 => 2, 22 => 2, 23 => 2, 24 => 2, 25 => 2, 26 => 2, 27 => 2, 28 => 2, 29 => 2, 30 => 2, 31 => 2, 32 => 2, 33 => 2);
      -- 
    begin -- 
      reqL_unguarded(33) <= RPIPE_Concat_input_pipe_268_inst_req_0;
      reqL_unguarded(32) <= RPIPE_Concat_input_pipe_431_inst_req_0;
      reqL_unguarded(31) <= RPIPE_Concat_input_pipe_381_inst_req_0;
      reqL_unguarded(30) <= RPIPE_Concat_input_pipe_406_inst_req_0;
      reqL_unguarded(29) <= RPIPE_Concat_input_pipe_243_inst_req_0;
      reqL_unguarded(28) <= RPIPE_Concat_input_pipe_218_inst_req_0;
      reqL_unguarded(27) <= RPIPE_Concat_input_pipe_256_inst_req_0;
      reqL_unguarded(26) <= RPIPE_Concat_input_pipe_343_inst_req_0;
      reqL_unguarded(25) <= RPIPE_Concat_input_pipe_393_inst_req_0;
      reqL_unguarded(24) <= RPIPE_Concat_input_pipe_231_inst_req_0;
      reqL_unguarded(23) <= RPIPE_Concat_input_pipe_306_inst_req_0;
      reqL_unguarded(22) <= RPIPE_Concat_input_pipe_331_inst_req_0;
      reqL_unguarded(21) <= RPIPE_Concat_input_pipe_418_inst_req_0;
      reqL_unguarded(20) <= RPIPE_Concat_input_pipe_368_inst_req_0;
      reqL_unguarded(19) <= RPIPE_Concat_input_pipe_293_inst_req_0;
      reqL_unguarded(18) <= RPIPE_Concat_input_pipe_356_inst_req_0;
      reqL_unguarded(17) <= RPIPE_Concat_input_pipe_281_inst_req_0;
      reqL_unguarded(16) <= RPIPE_Concat_input_pipe_318_inst_req_0;
      reqL_unguarded(15) <= RPIPE_Concat_input_pipe_573_inst_req_0;
      reqL_unguarded(14) <= RPIPE_Concat_input_pipe_604_inst_req_0;
      reqL_unguarded(13) <= RPIPE_Concat_input_pipe_586_inst_req_0;
      reqL_unguarded(12) <= RPIPE_Concat_input_pipe_622_inst_req_0;
      reqL_unguarded(11) <= RPIPE_Concat_input_pipe_640_inst_req_0;
      reqL_unguarded(10) <= RPIPE_Concat_input_pipe_658_inst_req_0;
      reqL_unguarded(9) <= RPIPE_Concat_input_pipe_676_inst_req_0;
      reqL_unguarded(8) <= RPIPE_Concat_input_pipe_694_inst_req_0;
      reqL_unguarded(7) <= RPIPE_Concat_input_pipe_780_inst_req_0;
      reqL_unguarded(6) <= RPIPE_Concat_input_pipe_793_inst_req_0;
      reqL_unguarded(5) <= RPIPE_Concat_input_pipe_811_inst_req_0;
      reqL_unguarded(4) <= RPIPE_Concat_input_pipe_829_inst_req_0;
      reqL_unguarded(3) <= RPIPE_Concat_input_pipe_847_inst_req_0;
      reqL_unguarded(2) <= RPIPE_Concat_input_pipe_865_inst_req_0;
      reqL_unguarded(1) <= RPIPE_Concat_input_pipe_883_inst_req_0;
      reqL_unguarded(0) <= RPIPE_Concat_input_pipe_901_inst_req_0;
      RPIPE_Concat_input_pipe_268_inst_ack_0 <= ackL_unguarded(33);
      RPIPE_Concat_input_pipe_431_inst_ack_0 <= ackL_unguarded(32);
      RPIPE_Concat_input_pipe_381_inst_ack_0 <= ackL_unguarded(31);
      RPIPE_Concat_input_pipe_406_inst_ack_0 <= ackL_unguarded(30);
      RPIPE_Concat_input_pipe_243_inst_ack_0 <= ackL_unguarded(29);
      RPIPE_Concat_input_pipe_218_inst_ack_0 <= ackL_unguarded(28);
      RPIPE_Concat_input_pipe_256_inst_ack_0 <= ackL_unguarded(27);
      RPIPE_Concat_input_pipe_343_inst_ack_0 <= ackL_unguarded(26);
      RPIPE_Concat_input_pipe_393_inst_ack_0 <= ackL_unguarded(25);
      RPIPE_Concat_input_pipe_231_inst_ack_0 <= ackL_unguarded(24);
      RPIPE_Concat_input_pipe_306_inst_ack_0 <= ackL_unguarded(23);
      RPIPE_Concat_input_pipe_331_inst_ack_0 <= ackL_unguarded(22);
      RPIPE_Concat_input_pipe_418_inst_ack_0 <= ackL_unguarded(21);
      RPIPE_Concat_input_pipe_368_inst_ack_0 <= ackL_unguarded(20);
      RPIPE_Concat_input_pipe_293_inst_ack_0 <= ackL_unguarded(19);
      RPIPE_Concat_input_pipe_356_inst_ack_0 <= ackL_unguarded(18);
      RPIPE_Concat_input_pipe_281_inst_ack_0 <= ackL_unguarded(17);
      RPIPE_Concat_input_pipe_318_inst_ack_0 <= ackL_unguarded(16);
      RPIPE_Concat_input_pipe_573_inst_ack_0 <= ackL_unguarded(15);
      RPIPE_Concat_input_pipe_604_inst_ack_0 <= ackL_unguarded(14);
      RPIPE_Concat_input_pipe_586_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_Concat_input_pipe_622_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_Concat_input_pipe_640_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_Concat_input_pipe_658_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_Concat_input_pipe_676_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_Concat_input_pipe_694_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_Concat_input_pipe_780_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_Concat_input_pipe_793_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_Concat_input_pipe_811_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_Concat_input_pipe_829_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_Concat_input_pipe_847_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_Concat_input_pipe_865_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_Concat_input_pipe_883_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_Concat_input_pipe_901_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(33) <= RPIPE_Concat_input_pipe_268_inst_req_1;
      reqR_unguarded(32) <= RPIPE_Concat_input_pipe_431_inst_req_1;
      reqR_unguarded(31) <= RPIPE_Concat_input_pipe_381_inst_req_1;
      reqR_unguarded(30) <= RPIPE_Concat_input_pipe_406_inst_req_1;
      reqR_unguarded(29) <= RPIPE_Concat_input_pipe_243_inst_req_1;
      reqR_unguarded(28) <= RPIPE_Concat_input_pipe_218_inst_req_1;
      reqR_unguarded(27) <= RPIPE_Concat_input_pipe_256_inst_req_1;
      reqR_unguarded(26) <= RPIPE_Concat_input_pipe_343_inst_req_1;
      reqR_unguarded(25) <= RPIPE_Concat_input_pipe_393_inst_req_1;
      reqR_unguarded(24) <= RPIPE_Concat_input_pipe_231_inst_req_1;
      reqR_unguarded(23) <= RPIPE_Concat_input_pipe_306_inst_req_1;
      reqR_unguarded(22) <= RPIPE_Concat_input_pipe_331_inst_req_1;
      reqR_unguarded(21) <= RPIPE_Concat_input_pipe_418_inst_req_1;
      reqR_unguarded(20) <= RPIPE_Concat_input_pipe_368_inst_req_1;
      reqR_unguarded(19) <= RPIPE_Concat_input_pipe_293_inst_req_1;
      reqR_unguarded(18) <= RPIPE_Concat_input_pipe_356_inst_req_1;
      reqR_unguarded(17) <= RPIPE_Concat_input_pipe_281_inst_req_1;
      reqR_unguarded(16) <= RPIPE_Concat_input_pipe_318_inst_req_1;
      reqR_unguarded(15) <= RPIPE_Concat_input_pipe_573_inst_req_1;
      reqR_unguarded(14) <= RPIPE_Concat_input_pipe_604_inst_req_1;
      reqR_unguarded(13) <= RPIPE_Concat_input_pipe_586_inst_req_1;
      reqR_unguarded(12) <= RPIPE_Concat_input_pipe_622_inst_req_1;
      reqR_unguarded(11) <= RPIPE_Concat_input_pipe_640_inst_req_1;
      reqR_unguarded(10) <= RPIPE_Concat_input_pipe_658_inst_req_1;
      reqR_unguarded(9) <= RPIPE_Concat_input_pipe_676_inst_req_1;
      reqR_unguarded(8) <= RPIPE_Concat_input_pipe_694_inst_req_1;
      reqR_unguarded(7) <= RPIPE_Concat_input_pipe_780_inst_req_1;
      reqR_unguarded(6) <= RPIPE_Concat_input_pipe_793_inst_req_1;
      reqR_unguarded(5) <= RPIPE_Concat_input_pipe_811_inst_req_1;
      reqR_unguarded(4) <= RPIPE_Concat_input_pipe_829_inst_req_1;
      reqR_unguarded(3) <= RPIPE_Concat_input_pipe_847_inst_req_1;
      reqR_unguarded(2) <= RPIPE_Concat_input_pipe_865_inst_req_1;
      reqR_unguarded(1) <= RPIPE_Concat_input_pipe_883_inst_req_1;
      reqR_unguarded(0) <= RPIPE_Concat_input_pipe_901_inst_req_1;
      RPIPE_Concat_input_pipe_268_inst_ack_1 <= ackR_unguarded(33);
      RPIPE_Concat_input_pipe_431_inst_ack_1 <= ackR_unguarded(32);
      RPIPE_Concat_input_pipe_381_inst_ack_1 <= ackR_unguarded(31);
      RPIPE_Concat_input_pipe_406_inst_ack_1 <= ackR_unguarded(30);
      RPIPE_Concat_input_pipe_243_inst_ack_1 <= ackR_unguarded(29);
      RPIPE_Concat_input_pipe_218_inst_ack_1 <= ackR_unguarded(28);
      RPIPE_Concat_input_pipe_256_inst_ack_1 <= ackR_unguarded(27);
      RPIPE_Concat_input_pipe_343_inst_ack_1 <= ackR_unguarded(26);
      RPIPE_Concat_input_pipe_393_inst_ack_1 <= ackR_unguarded(25);
      RPIPE_Concat_input_pipe_231_inst_ack_1 <= ackR_unguarded(24);
      RPIPE_Concat_input_pipe_306_inst_ack_1 <= ackR_unguarded(23);
      RPIPE_Concat_input_pipe_331_inst_ack_1 <= ackR_unguarded(22);
      RPIPE_Concat_input_pipe_418_inst_ack_1 <= ackR_unguarded(21);
      RPIPE_Concat_input_pipe_368_inst_ack_1 <= ackR_unguarded(20);
      RPIPE_Concat_input_pipe_293_inst_ack_1 <= ackR_unguarded(19);
      RPIPE_Concat_input_pipe_356_inst_ack_1 <= ackR_unguarded(18);
      RPIPE_Concat_input_pipe_281_inst_ack_1 <= ackR_unguarded(17);
      RPIPE_Concat_input_pipe_318_inst_ack_1 <= ackR_unguarded(16);
      RPIPE_Concat_input_pipe_573_inst_ack_1 <= ackR_unguarded(15);
      RPIPE_Concat_input_pipe_604_inst_ack_1 <= ackR_unguarded(14);
      RPIPE_Concat_input_pipe_586_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_Concat_input_pipe_622_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_Concat_input_pipe_640_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_Concat_input_pipe_658_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_Concat_input_pipe_676_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_Concat_input_pipe_694_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_Concat_input_pipe_780_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_Concat_input_pipe_793_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_Concat_input_pipe_811_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_Concat_input_pipe_829_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_Concat_input_pipe_847_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_Concat_input_pipe_865_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_Concat_input_pipe_883_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_Concat_input_pipe_901_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      guard_vector(18)  <=  '1';
      guard_vector(19)  <=  '1';
      guard_vector(20)  <=  '1';
      guard_vector(21)  <=  '1';
      guard_vector(22)  <=  '1';
      guard_vector(23)  <=  '1';
      guard_vector(24)  <=  '1';
      guard_vector(25)  <=  '1';
      guard_vector(26)  <=  '1';
      guard_vector(27)  <=  '1';
      guard_vector(28)  <=  '1';
      guard_vector(29)  <=  '1';
      guard_vector(30)  <=  '1';
      guard_vector(31)  <=  '1';
      guard_vector(32)  <=  '1';
      guard_vector(33)  <=  '1';
      call14_269 <= data_out(271 downto 264);
      call73_432 <= data_out(263 downto 256);
      call55_382 <= data_out(255 downto 248);
      call64_407 <= data_out(247 downto 240);
      call5_244 <= data_out(239 downto 232);
      call_219 <= data_out(231 downto 224);
      call10_257 <= data_out(223 downto 216);
      call41_344 <= data_out(215 downto 208);
      call59_394 <= data_out(207 downto 200);
      call2_232 <= data_out(199 downto 192);
      call28_307 <= data_out(191 downto 184);
      call37_332 <= data_out(183 downto 176);
      call68_419 <= data_out(175 downto 168);
      call50_369 <= data_out(167 downto 160);
      call23_294 <= data_out(159 downto 152);
      call46_357 <= data_out(151 downto 144);
      call19_282 <= data_out(143 downto 136);
      call32_319 <= data_out(135 downto 128);
      call118_574 <= data_out(127 downto 120);
      call128_605 <= data_out(119 downto 112);
      call122_587 <= data_out(111 downto 104);
      call134_623 <= data_out(103 downto 96);
      call140_641 <= data_out(95 downto 88);
      call146_659 <= data_out(87 downto 80);
      call152_677 <= data_out(79 downto 72);
      call158_695 <= data_out(71 downto 64);
      call174_781 <= data_out(63 downto 56);
      call178_794 <= data_out(55 downto 48);
      call184_812 <= data_out(47 downto 40);
      call190_830 <= data_out(39 downto 32);
      call196_848 <= data_out(31 downto 24);
      call202_866 <= data_out(23 downto 16);
      call208_884 <= data_out(15 downto 8);
      call214_902 <= data_out(7 downto 0);
      Concat_input_pipe_read_0_gI: SplitGuardInterface generic map(name => "Concat_input_pipe_read_0_gI", nreqs => 34, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Concat_input_pipe_read_0: InputPortRevised -- 
        generic map ( name => "Concat_input_pipe_read_0", data_width => 8,  num_reqs => 34,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Concat_input_pipe_pipe_read_req(0),
          oack => Concat_input_pipe_pipe_read_ack(0),
          odata => Concat_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Concat_output_pipe_1037_inst WPIPE_Concat_output_pipe_1040_inst WPIPE_Concat_output_pipe_1043_inst WPIPE_Concat_output_pipe_1046_inst WPIPE_Concat_output_pipe_1049_inst WPIPE_Concat_output_pipe_1052_inst WPIPE_Concat_output_pipe_1055_inst WPIPE_Concat_output_pipe_1058_inst WPIPE_Concat_output_pipe_1201_inst WPIPE_Concat_output_pipe_1204_inst WPIPE_Concat_output_pipe_1207_inst WPIPE_Concat_output_pipe_1210_inst WPIPE_Concat_output_pipe_1213_inst WPIPE_Concat_output_pipe_1216_inst WPIPE_Concat_output_pipe_1219_inst WPIPE_Concat_output_pipe_1222_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal sample_req, sample_ack : BooleanArray( 15 downto 0);
      signal update_req, update_ack : BooleanArray( 15 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 15 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 15 downto 0);
      signal guard_vector : std_logic_vector( 15 downto 0);
      constant inBUFs : IntegerArray(15 downto 0) := (15 => 0, 14 => 0, 13 => 0, 12 => 0, 11 => 0, 10 => 0, 9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(15 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false);
      constant guardBuffering: IntegerArray(15 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2);
      -- 
    begin -- 
      sample_req_unguarded(15) <= WPIPE_Concat_output_pipe_1037_inst_req_0;
      sample_req_unguarded(14) <= WPIPE_Concat_output_pipe_1040_inst_req_0;
      sample_req_unguarded(13) <= WPIPE_Concat_output_pipe_1043_inst_req_0;
      sample_req_unguarded(12) <= WPIPE_Concat_output_pipe_1046_inst_req_0;
      sample_req_unguarded(11) <= WPIPE_Concat_output_pipe_1049_inst_req_0;
      sample_req_unguarded(10) <= WPIPE_Concat_output_pipe_1052_inst_req_0;
      sample_req_unguarded(9) <= WPIPE_Concat_output_pipe_1055_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_Concat_output_pipe_1058_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_Concat_output_pipe_1201_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_Concat_output_pipe_1204_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_Concat_output_pipe_1207_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_Concat_output_pipe_1210_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_Concat_output_pipe_1213_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_Concat_output_pipe_1216_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_Concat_output_pipe_1219_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_Concat_output_pipe_1222_inst_req_0;
      WPIPE_Concat_output_pipe_1037_inst_ack_0 <= sample_ack_unguarded(15);
      WPIPE_Concat_output_pipe_1040_inst_ack_0 <= sample_ack_unguarded(14);
      WPIPE_Concat_output_pipe_1043_inst_ack_0 <= sample_ack_unguarded(13);
      WPIPE_Concat_output_pipe_1046_inst_ack_0 <= sample_ack_unguarded(12);
      WPIPE_Concat_output_pipe_1049_inst_ack_0 <= sample_ack_unguarded(11);
      WPIPE_Concat_output_pipe_1052_inst_ack_0 <= sample_ack_unguarded(10);
      WPIPE_Concat_output_pipe_1055_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_Concat_output_pipe_1058_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_Concat_output_pipe_1201_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_Concat_output_pipe_1204_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_Concat_output_pipe_1207_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_Concat_output_pipe_1210_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_Concat_output_pipe_1213_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_Concat_output_pipe_1216_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_Concat_output_pipe_1219_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_Concat_output_pipe_1222_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(15) <= WPIPE_Concat_output_pipe_1037_inst_req_1;
      update_req_unguarded(14) <= WPIPE_Concat_output_pipe_1040_inst_req_1;
      update_req_unguarded(13) <= WPIPE_Concat_output_pipe_1043_inst_req_1;
      update_req_unguarded(12) <= WPIPE_Concat_output_pipe_1046_inst_req_1;
      update_req_unguarded(11) <= WPIPE_Concat_output_pipe_1049_inst_req_1;
      update_req_unguarded(10) <= WPIPE_Concat_output_pipe_1052_inst_req_1;
      update_req_unguarded(9) <= WPIPE_Concat_output_pipe_1055_inst_req_1;
      update_req_unguarded(8) <= WPIPE_Concat_output_pipe_1058_inst_req_1;
      update_req_unguarded(7) <= WPIPE_Concat_output_pipe_1201_inst_req_1;
      update_req_unguarded(6) <= WPIPE_Concat_output_pipe_1204_inst_req_1;
      update_req_unguarded(5) <= WPIPE_Concat_output_pipe_1207_inst_req_1;
      update_req_unguarded(4) <= WPIPE_Concat_output_pipe_1210_inst_req_1;
      update_req_unguarded(3) <= WPIPE_Concat_output_pipe_1213_inst_req_1;
      update_req_unguarded(2) <= WPIPE_Concat_output_pipe_1216_inst_req_1;
      update_req_unguarded(1) <= WPIPE_Concat_output_pipe_1219_inst_req_1;
      update_req_unguarded(0) <= WPIPE_Concat_output_pipe_1222_inst_req_1;
      WPIPE_Concat_output_pipe_1037_inst_ack_1 <= update_ack_unguarded(15);
      WPIPE_Concat_output_pipe_1040_inst_ack_1 <= update_ack_unguarded(14);
      WPIPE_Concat_output_pipe_1043_inst_ack_1 <= update_ack_unguarded(13);
      WPIPE_Concat_output_pipe_1046_inst_ack_1 <= update_ack_unguarded(12);
      WPIPE_Concat_output_pipe_1049_inst_ack_1 <= update_ack_unguarded(11);
      WPIPE_Concat_output_pipe_1052_inst_ack_1 <= update_ack_unguarded(10);
      WPIPE_Concat_output_pipe_1055_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_Concat_output_pipe_1058_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_Concat_output_pipe_1201_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_Concat_output_pipe_1204_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_Concat_output_pipe_1207_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_Concat_output_pipe_1210_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_Concat_output_pipe_1213_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_Concat_output_pipe_1216_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_Concat_output_pipe_1219_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_Concat_output_pipe_1222_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      data_in <= conv281_1036 & conv275_1026 & conv269_1016 & conv263_1006 & conv257_996 & conv251_986 & conv245_976 & conv239_966 & conv356_1200 & conv350_1190 & conv344_1180 & conv338_1170 & conv332_1160 & conv326_1150 & conv320_1140 & conv314_1130;
      Concat_output_pipe_write_0_gI: SplitGuardInterface generic map(name => "Concat_output_pipe_write_0_gI", nreqs => 16, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Concat_output_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "Concat_output_pipe", data_width => 8, num_reqs => 16, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Concat_output_pipe_pipe_write_req(0),
          oack => Concat_output_pipe_pipe_write_ack(0),
          odata => Concat_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared call operator group (0) : call_stmt_938_call call_stmt_952_call 
    timer_call_group_0: Block -- 
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_938_call_req_0;
      reqL_unguarded(0) <= call_stmt_952_call_req_0;
      call_stmt_938_call_ack_0 <= ackL_unguarded(1);
      call_stmt_952_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_938_call_req_1;
      reqR_unguarded(0) <= call_stmt_952_call_req_1;
      call_stmt_938_call_ack_1 <= ackR_unguarded(1);
      call_stmt_952_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      timer_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      timer_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      timer_call_group_0_gI: SplitGuardInterface generic map(name => "timer_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      call226_938 <= data_out(127 downto 64);
      call232_952 <= data_out(63 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 2,
        nreqs => 2,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => timer_call_reqs(0),
          ackR => timer_call_acks(0),
          tagR => timer_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => timer_return_acks(0), -- cross-over
          ackL => timer_return_reqs(0), -- cross-over
          dataL => timer_return_data(63 downto 0),
          tagL => timer_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_949_call 
    concat_core_call_group_1: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_949_call_req_0;
      call_stmt_949_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_949_call_req_1;
      call_stmt_949_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      concat_core_call_group_1_gI: SplitGuardInterface generic map(name => "concat_core_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= shr378_485 & shr111379_491 & mul103_479;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 64,
        owidth => 64,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => concat_core_call_reqs(0),
          ackR => concat_core_call_acks(0),
          dataR => concat_core_call_data(63 downto 0),
          tagR => concat_core_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => concat_core_return_acks(0), -- cross-over
          ackL => concat_core_return_reqs(0), -- cross-over
          tagL => concat_core_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- 
  end Block; -- data_path
  -- 
end concat_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity concat_core is -- 
  generic (tag_length : integer); 
  port ( -- 
    input1_count : in  std_logic_vector(15 downto 0);
    input2_count : in  std_logic_vector(15 downto 0);
    output_size : in  std_logic_vector(31 downto 0);
    readModule1_call_reqs : out  std_logic_vector(0 downto 0);
    readModule1_call_acks : in   std_logic_vector(0 downto 0);
    readModule1_call_data : out  std_logic_vector(39 downto 0);
    readModule1_call_tag  :  out  std_logic_vector(1 downto 0);
    readModule1_return_reqs : out  std_logic_vector(0 downto 0);
    readModule1_return_acks : in   std_logic_vector(0 downto 0);
    readModule1_return_data : in   std_logic_vector(63 downto 0);
    readModule1_return_tag :  in   std_logic_vector(1 downto 0);
    writeModule1_call_reqs : out  std_logic_vector(0 downto 0);
    writeModule1_call_acks : in   std_logic_vector(0 downto 0);
    writeModule1_call_data : out  std_logic_vector(103 downto 0);
    writeModule1_call_tag  :  out  std_logic_vector(0 downto 0);
    writeModule1_return_reqs : out  std_logic_vector(0 downto 0);
    writeModule1_return_acks : in   std_logic_vector(0 downto 0);
    writeModule1_return_data : in   std_logic_vector(0 downto 0);
    writeModule1_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity concat_core;
architecture concat_core_arch of concat_core is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal input1_count_buffer :  std_logic_vector(15 downto 0);
  signal input1_count_update_enable: Boolean;
  signal input2_count_buffer :  std_logic_vector(15 downto 0);
  signal input2_count_update_enable: Boolean;
  signal output_size_buffer :  std_logic_vector(31 downto 0);
  signal output_size_update_enable: Boolean;
  -- output port buffer signals
  signal concat_core_CP_345_start: Boolean;
  signal concat_core_CP_345_symbol: Boolean;
  -- volatile/operator module components. 
  component readModule1 is -- 
    generic (tag_length : integer); 
    port ( -- 
      index : in  std_logic_vector(7 downto 0);
      address : in  std_logic_vector(31 downto 0);
      data : out  std_logic_vector(63 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(15 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component writeModule1 is -- 
    generic (tag_length : integer); 
    port ( -- 
      index : in  std_logic_vector(7 downto 0);
      address : in  std_logic_vector(31 downto 0);
      data : in  std_logic_vector(63 downto 0);
      done : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(15 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_135_call_req_1 : boolean;
  signal call_stmt_135_call_ack_1 : boolean;
  signal W_cmp_143_delayed_15_0_142_inst_ack_0 : boolean;
  signal SUB_u32_u32_201_inst_req_0 : boolean;
  signal call_stmt_135_call_ack_0 : boolean;
  signal W_cmp_143_delayed_15_0_142_inst_req_0 : boolean;
  signal call_stmt_135_call_req_0 : boolean;
  signal W_add_out_149_delayed_15_0_151_inst_ack_1 : boolean;
  signal W_add_out_149_delayed_15_0_151_inst_req_1 : boolean;
  signal call_stmt_158_call_ack_1 : boolean;
  signal next_add_out_197_111_buf_req_0 : boolean;
  signal next_add_out_197_111_buf_ack_0 : boolean;
  signal next_add_out_197_111_buf_req_1 : boolean;
  signal next_add_out_197_111_buf_ack_1 : boolean;
  signal next_count_inp1_176_123_buf_ack_1 : boolean;
  signal W_add_out_149_delayed_15_0_151_inst_ack_0 : boolean;
  signal call_stmt_158_call_req_1 : boolean;
  signal SUB_u16_u16_162_inst_ack_1 : boolean;
  signal SUB_u16_u16_162_inst_req_1 : boolean;
  signal next_count_inp1_176_123_buf_req_1 : boolean;
  signal W_add_out_149_delayed_15_0_151_inst_req_0 : boolean;
  signal next_count_inp1_176_123_buf_ack_0 : boolean;
  signal do_while_stmt_106_branch_ack_1 : boolean;
  signal call_stmt_158_call_ack_0 : boolean;
  signal call_stmt_158_call_req_0 : boolean;
  signal W_cmp_143_delayed_15_0_142_inst_ack_1 : boolean;
  signal next_count_inp1_176_123_buf_req_0 : boolean;
  signal do_while_stmt_106_branch_ack_0 : boolean;
  signal W_cmp_143_delayed_15_0_142_inst_req_1 : boolean;
  signal do_while_stmt_106_branch_req_0 : boolean;
  signal phi_stmt_108_req_1 : boolean;
  signal phi_stmt_108_req_0 : boolean;
  signal phi_stmt_108_ack_0 : boolean;
  signal SUB_u16_u16_162_inst_ack_0 : boolean;
  signal phi_stmt_112_req_1 : boolean;
  signal phi_stmt_112_req_0 : boolean;
  signal phi_stmt_112_ack_0 : boolean;
  signal call_stmt_141_call_ack_1 : boolean;
  signal SUB_u16_u16_162_inst_req_0 : boolean;
  signal next_add_inp1_184_115_buf_req_0 : boolean;
  signal next_add_inp1_184_115_buf_ack_0 : boolean;
  signal next_add_inp1_184_115_buf_req_1 : boolean;
  signal next_add_inp1_184_115_buf_ack_1 : boolean;
  signal call_stmt_141_call_req_1 : boolean;
  signal phi_stmt_116_req_1 : boolean;
  signal SUB_u32_u32_201_inst_ack_1 : boolean;
  signal phi_stmt_116_req_0 : boolean;
  signal SUB_u32_u32_201_inst_req_1 : boolean;
  signal phi_stmt_116_ack_0 : boolean;
  signal SUB_u32_u32_201_inst_ack_0 : boolean;
  signal call_stmt_141_call_ack_0 : boolean;
  signal call_stmt_141_call_req_0 : boolean;
  signal next_add_inp2_192_119_buf_req_0 : boolean;
  signal next_add_inp2_192_119_buf_ack_0 : boolean;
  signal next_add_inp2_192_119_buf_req_1 : boolean;
  signal next_add_inp2_192_119_buf_ack_1 : boolean;
  signal phi_stmt_120_req_1 : boolean;
  signal phi_stmt_120_req_0 : boolean;
  signal phi_stmt_120_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "concat_core_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 64) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(15 downto 0) <= input1_count;
  input1_count_buffer <= in_buffer_data_out(15 downto 0);
  in_buffer_data_in(31 downto 16) <= input2_count;
  input2_count_buffer <= in_buffer_data_out(31 downto 16);
  in_buffer_data_in(63 downto 32) <= output_size;
  output_size_buffer <= in_buffer_data_out(63 downto 32);
  in_buffer_data_in(tag_length + 63 downto 64) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 63 downto 64);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  concat_core_CP_345_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "concat_core_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= concat_core_CP_345_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= concat_core_CP_345_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= concat_core_CP_345_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  concat_core_CP_345: Block -- control-path 
    signal concat_core_CP_345_elements: BooleanArray(121 downto 0);
    -- 
  begin -- 
    concat_core_CP_345_elements(0) <= concat_core_CP_345_start;
    concat_core_CP_345_symbol <= concat_core_CP_345_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_69/$entry
      -- CP-element group 0: 	 branch_block_stmt_69/branch_block_stmt_69__entry__
      -- CP-element group 0: 	 branch_block_stmt_69/assign_stmt_72_to_assign_stmt_105__entry__
      -- CP-element group 0: 	 branch_block_stmt_69/assign_stmt_72_to_assign_stmt_105__exit__
      -- CP-element group 0: 	 branch_block_stmt_69/do_while_stmt_106__entry__
      -- CP-element group 0: 	 branch_block_stmt_69/assign_stmt_72_to_assign_stmt_105/$entry
      -- CP-element group 0: 	 branch_block_stmt_69/assign_stmt_72_to_assign_stmt_105/$exit
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	121 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_69/$exit
      -- CP-element group 1: 	 branch_block_stmt_69/branch_block_stmt_69__exit__
      -- CP-element group 1: 	 branch_block_stmt_69/do_while_stmt_106__exit__
      -- 
    concat_core_CP_345_elements(1) <= concat_core_CP_345_elements(121);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_69/do_while_stmt_106/$entry
      -- CP-element group 2: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106__entry__
      -- 
    concat_core_CP_345_elements(2) <= concat_core_CP_345_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	121 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106__exit__
      -- 
    -- Element group concat_core_CP_345_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_69/do_while_stmt_106/loop_back
      -- 
    -- Element group concat_core_CP_345_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	119 
    -- CP-element group 5: 	120 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_69/do_while_stmt_106/loop_taken/$entry
      -- CP-element group 5: 	 branch_block_stmt_69/do_while_stmt_106/condition_done
      -- CP-element group 5: 	 branch_block_stmt_69/do_while_stmt_106/loop_exit/$entry
      -- 
    concat_core_CP_345_elements(5) <= concat_core_CP_345_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	118 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_69/do_while_stmt_106/loop_body_done
      -- 
    concat_core_CP_345_elements(6) <= concat_core_CP_345_elements(118);
    -- CP-element group 7:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	19 
    -- CP-element group 7: 	38 
    -- CP-element group 7: 	57 
    -- CP-element group 7: 	76 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/back_edge_to_loop_body
      -- 
    concat_core_CP_345_elements(7) <= concat_core_CP_345_elements(4);
    -- CP-element group 8:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	21 
    -- CP-element group 8: 	59 
    -- CP-element group 8: 	40 
    -- CP-element group 8: 	78 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/first_time_through_loop_body
      -- 
    concat_core_CP_345_elements(8) <= concat_core_CP_345_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	33 
    -- CP-element group 9: 	32 
    -- CP-element group 9: 	52 
    -- CP-element group 9: 	51 
    -- CP-element group 9: 	109 
    -- CP-element group 9: 	113 
    -- CP-element group 9: 	117 
    -- CP-element group 9: 	70 
    -- CP-element group 9: 	71 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/loop_body_start
      -- 
    -- Element group concat_core_CP_345_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	14 
    -- CP-element group 10: 	112 
    -- CP-element group 10: 	116 
    -- CP-element group 10: 	117 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/condition_evaluated
      -- 
    condition_evaluated_374_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_374_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_core_CP_345_elements(10), ack => do_while_stmt_106_branch_req_0); -- 
    concat_core_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 15);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 31) := "concat_core_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= concat_core_CP_345_elements(14) & concat_core_CP_345_elements(112) & concat_core_CP_345_elements(116) & concat_core_CP_345_elements(117);
      gj_concat_core_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_core_CP_345_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	15 
    -- CP-element group 11: 	32 
    -- CP-element group 11: 	51 
    -- CP-element group 11: 	70 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	34 
    -- CP-element group 11: 	53 
    -- CP-element group 11: 	72 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/phi_stmt_108_sample_start__ps
      -- 
    concat_core_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 31) := "concat_core_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= concat_core_CP_345_elements(15) & concat_core_CP_345_elements(32) & concat_core_CP_345_elements(51) & concat_core_CP_345_elements(70) & concat_core_CP_345_elements(14);
      gj_concat_core_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_core_CP_345_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	17 
    -- CP-element group 12: 	54 
    -- CP-element group 12: 	35 
    -- CP-element group 12: 	73 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	110 
    -- CP-element group 12: 	118 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	15 
    -- CP-element group 12: 	32 
    -- CP-element group 12: 	51 
    -- CP-element group 12: 	70 
    -- CP-element group 12:  members (5) 
      -- CP-element group 12: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/phi_stmt_108_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/phi_stmt_112_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/phi_stmt_116_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/phi_stmt_120_sample_completed_
      -- 
    concat_core_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 15);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 31) := "concat_core_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= concat_core_CP_345_elements(17) & concat_core_CP_345_elements(54) & concat_core_CP_345_elements(35) & concat_core_CP_345_elements(73);
      gj_concat_core_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_core_CP_345_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	16 
    -- CP-element group 13: 	33 
    -- CP-element group 13: 	52 
    -- CP-element group 13: 	71 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	36 
    -- CP-element group 13: 	55 
    -- CP-element group 13: 	74 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/phi_stmt_108_update_start__ps
      -- 
    concat_core_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 15);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 31) := "concat_core_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= concat_core_CP_345_elements(16) & concat_core_CP_345_elements(33) & concat_core_CP_345_elements(52) & concat_core_CP_345_elements(71);
      gj_concat_core_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_core_CP_345_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	18 
    -- CP-element group 14: 	56 
    -- CP-element group 14: 	37 
    -- CP-element group 14: 	75 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/aggregated_phi_update_ack
      -- 
    concat_core_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 15);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 31) := "concat_core_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= concat_core_CP_345_elements(18) & concat_core_CP_345_elements(56) & concat_core_CP_345_elements(37) & concat_core_CP_345_elements(75);
      gj_concat_core_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_core_CP_345_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/phi_stmt_108_sample_start_
      -- 
    concat_core_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "concat_core_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_core_CP_345_elements(9) & concat_core_CP_345_elements(12);
      gj_concat_core_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_core_CP_345_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	103 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/phi_stmt_108_update_start_
      -- 
    concat_core_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "concat_core_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_core_CP_345_elements(9) & concat_core_CP_345_elements(103);
      gj_concat_core_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_core_CP_345_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	12 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/phi_stmt_108_sample_completed__ps
      -- 
    -- Element group concat_core_CP_345_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	14 
    -- CP-element group 18: 	101 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/phi_stmt_108_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/phi_stmt_108_update_completed__ps
      -- 
    -- Element group concat_core_CP_345_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	7 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/phi_stmt_108_loopback_trigger
      -- 
    concat_core_CP_345_elements(19) <= concat_core_CP_345_elements(7);
    -- CP-element group 20:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/phi_stmt_108_loopback_sample_req
      -- CP-element group 20: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/phi_stmt_108_loopback_sample_req_ps
      -- 
    phi_stmt_108_loopback_sample_req_389_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_108_loopback_sample_req_389_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_core_CP_345_elements(20), ack => phi_stmt_108_req_1); -- 
    -- Element group concat_core_CP_345_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	8 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/phi_stmt_108_entry_trigger
      -- 
    concat_core_CP_345_elements(21) <= concat_core_CP_345_elements(8);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/phi_stmt_108_entry_sample_req
      -- CP-element group 22: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/phi_stmt_108_entry_sample_req_ps
      -- 
    phi_stmt_108_entry_sample_req_392_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_108_entry_sample_req_392_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_core_CP_345_elements(22), ack => phi_stmt_108_req_0); -- 
    -- Element group concat_core_CP_345_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/phi_stmt_108_phi_mux_ack
      -- CP-element group 23: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/phi_stmt_108_phi_mux_ack_ps
      -- 
    phi_stmt_108_phi_mux_ack_395_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_108_ack_0, ack => concat_core_CP_345_elements(23)); -- 
    -- CP-element group 24:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (4) 
      -- CP-element group 24: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_add_out_init_110_sample_start__ps
      -- CP-element group 24: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_add_out_init_110_sample_completed__ps
      -- CP-element group 24: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_add_out_init_110_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_add_out_init_110_sample_completed_
      -- 
    -- Element group concat_core_CP_345_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_add_out_init_110_update_start_
      -- CP-element group 25: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_add_out_init_110_update_start__ps
      -- 
    -- Element group concat_core_CP_345_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_add_out_init_110_update_completed__ps
      -- 
    concat_core_CP_345_elements(26) <= concat_core_CP_345_elements(27);
    -- CP-element group 27:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	26 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_add_out_init_110_update_completed_
      -- 
    -- Element group concat_core_CP_345_elements(27) is a control-delay.
    cp_element_27_delay: control_delay_element  generic map(name => " 27_delay", delay_value => 1)  port map(req => concat_core_CP_345_elements(25), ack => concat_core_CP_345_elements(27), clk => clk, reset =>reset);
    -- CP-element group 28:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_next_add_out_111_sample_start__ps
      -- CP-element group 28: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_next_add_out_111_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_next_add_out_111_Sample/$entry
      -- CP-element group 28: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_next_add_out_111_Sample/req
      -- 
    req_416_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_416_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_core_CP_345_elements(28), ack => next_add_out_197_111_buf_req_0); -- 
    -- Element group concat_core_CP_345_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_next_add_out_111_update_start__ps
      -- CP-element group 29: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_next_add_out_111_update_start_
      -- CP-element group 29: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_next_add_out_111_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_next_add_out_111_Update/req
      -- 
    req_421_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_421_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_core_CP_345_elements(29), ack => next_add_out_197_111_buf_req_1); -- 
    -- Element group concat_core_CP_345_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_next_add_out_111_sample_completed__ps
      -- CP-element group 30: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_next_add_out_111_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_next_add_out_111_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_next_add_out_111_Sample/ack
      -- 
    ack_417_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_add_out_197_111_buf_ack_0, ack => concat_core_CP_345_elements(30)); -- 
    -- CP-element group 31:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_next_add_out_111_update_completed__ps
      -- CP-element group 31: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_next_add_out_111_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_next_add_out_111_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_next_add_out_111_Update/ack
      -- 
    ack_422_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_add_out_197_111_buf_ack_1, ack => concat_core_CP_345_elements(31)); -- 
    -- CP-element group 32:  join  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	9 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	12 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	11 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/phi_stmt_112_sample_start_
      -- 
    concat_core_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "concat_core_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_core_CP_345_elements(9) & concat_core_CP_345_elements(12);
      gj_concat_core_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_core_CP_345_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  join  transition  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	9 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	91 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	13 
    -- CP-element group 33:  members (1) 
      -- CP-element group 33: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/phi_stmt_112_update_start_
      -- 
    concat_core_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "concat_core_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_core_CP_345_elements(9) & concat_core_CP_345_elements(91);
      gj_concat_core_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_core_CP_345_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	11 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (1) 
      -- CP-element group 34: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/phi_stmt_112_sample_start__ps
      -- 
    concat_core_CP_345_elements(34) <= concat_core_CP_345_elements(11);
    -- CP-element group 35:  join  transition  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	12 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/phi_stmt_112_sample_completed__ps
      -- 
    -- Element group concat_core_CP_345_elements(35) is bound as output of CP function.
    -- CP-element group 36:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	13 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/phi_stmt_112_update_start__ps
      -- 
    concat_core_CP_345_elements(36) <= concat_core_CP_345_elements(13);
    -- CP-element group 37:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	14 
    -- CP-element group 37: 	89 
    -- CP-element group 37:  members (2) 
      -- CP-element group 37: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/phi_stmt_112_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/phi_stmt_112_update_completed__ps
      -- 
    -- Element group concat_core_CP_345_elements(37) is bound as output of CP function.
    -- CP-element group 38:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	7 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/phi_stmt_112_loopback_trigger
      -- 
    concat_core_CP_345_elements(38) <= concat_core_CP_345_elements(7);
    -- CP-element group 39:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (2) 
      -- CP-element group 39: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/phi_stmt_112_loopback_sample_req
      -- CP-element group 39: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/phi_stmt_112_loopback_sample_req_ps
      -- 
    phi_stmt_112_loopback_sample_req_433_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_112_loopback_sample_req_433_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_core_CP_345_elements(39), ack => phi_stmt_112_req_1); -- 
    -- Element group concat_core_CP_345_elements(39) is bound as output of CP function.
    -- CP-element group 40:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	8 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/phi_stmt_112_entry_trigger
      -- 
    concat_core_CP_345_elements(40) <= concat_core_CP_345_elements(8);
    -- CP-element group 41:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (2) 
      -- CP-element group 41: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/phi_stmt_112_entry_sample_req
      -- CP-element group 41: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/phi_stmt_112_entry_sample_req_ps
      -- 
    phi_stmt_112_entry_sample_req_436_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_112_entry_sample_req_436_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_core_CP_345_elements(41), ack => phi_stmt_112_req_0); -- 
    -- Element group concat_core_CP_345_elements(41) is bound as output of CP function.
    -- CP-element group 42:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (2) 
      -- CP-element group 42: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/phi_stmt_112_phi_mux_ack
      -- CP-element group 42: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/phi_stmt_112_phi_mux_ack_ps
      -- 
    phi_stmt_112_phi_mux_ack_439_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_112_ack_0, ack => concat_core_CP_345_elements(42)); -- 
    -- CP-element group 43:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (4) 
      -- CP-element group 43: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_add_inp1_init_114_sample_start__ps
      -- CP-element group 43: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_add_inp1_init_114_sample_completed__ps
      -- CP-element group 43: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_add_inp1_init_114_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_add_inp1_init_114_sample_completed_
      -- 
    -- Element group concat_core_CP_345_elements(43) is bound as output of CP function.
    -- CP-element group 44:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	46 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_add_inp1_init_114_update_start__ps
      -- CP-element group 44: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_add_inp1_init_114_update_start_
      -- 
    -- Element group concat_core_CP_345_elements(44) is bound as output of CP function.
    -- CP-element group 45:  join  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	46 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_add_inp1_init_114_update_completed__ps
      -- 
    concat_core_CP_345_elements(45) <= concat_core_CP_345_elements(46);
    -- CP-element group 46:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	44 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	45 
    -- CP-element group 46:  members (1) 
      -- CP-element group 46: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_add_inp1_init_114_update_completed_
      -- 
    -- Element group concat_core_CP_345_elements(46) is a control-delay.
    cp_element_46_delay: control_delay_element  generic map(name => " 46_delay", delay_value => 1)  port map(req => concat_core_CP_345_elements(44), ack => concat_core_CP_345_elements(46), clk => clk, reset =>reset);
    -- CP-element group 47:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	49 
    -- CP-element group 47:  members (4) 
      -- CP-element group 47: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_next_add_inp1_115_sample_start__ps
      -- CP-element group 47: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_next_add_inp1_115_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_next_add_inp1_115_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_next_add_inp1_115_Sample/req
      -- 
    req_460_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_460_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_core_CP_345_elements(47), ack => next_add_inp1_184_115_buf_req_0); -- 
    -- Element group concat_core_CP_345_elements(47) is bound as output of CP function.
    -- CP-element group 48:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	50 
    -- CP-element group 48:  members (4) 
      -- CP-element group 48: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_next_add_inp1_115_update_start__ps
      -- CP-element group 48: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_next_add_inp1_115_update_start_
      -- CP-element group 48: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_next_add_inp1_115_Update/$entry
      -- CP-element group 48: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_next_add_inp1_115_Update/req
      -- 
    req_465_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_465_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_core_CP_345_elements(48), ack => next_add_inp1_184_115_buf_req_1); -- 
    -- Element group concat_core_CP_345_elements(48) is bound as output of CP function.
    -- CP-element group 49:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	47 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (4) 
      -- CP-element group 49: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_next_add_inp1_115_sample_completed__ps
      -- CP-element group 49: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_next_add_inp1_115_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_next_add_inp1_115_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_next_add_inp1_115_Sample/ack
      -- 
    ack_461_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_add_inp1_184_115_buf_ack_0, ack => concat_core_CP_345_elements(49)); -- 
    -- CP-element group 50:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	48 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (4) 
      -- CP-element group 50: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_next_add_inp1_115_update_completed__ps
      -- CP-element group 50: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_next_add_inp1_115_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_next_add_inp1_115_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_next_add_inp1_115_Update/ack
      -- 
    ack_466_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_add_inp1_184_115_buf_ack_1, ack => concat_core_CP_345_elements(50)); -- 
    -- CP-element group 51:  join  transition  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	9 
    -- CP-element group 51: marked-predecessors 
    -- CP-element group 51: 	12 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	11 
    -- CP-element group 51:  members (1) 
      -- CP-element group 51: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/phi_stmt_116_sample_start_
      -- 
    concat_core_cp_element_group_51: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "concat_core_cp_element_group_51"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_core_CP_345_elements(9) & concat_core_CP_345_elements(12);
      gj_concat_core_cp_element_group_51 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_core_CP_345_elements(51), clk => clk, reset => reset); --
    end block;
    -- CP-element group 52:  join  transition  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	9 
    -- CP-element group 52: marked-predecessors 
    -- CP-element group 52: 	95 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	13 
    -- CP-element group 52:  members (1) 
      -- CP-element group 52: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/phi_stmt_116_update_start_
      -- 
    concat_core_cp_element_group_52: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "concat_core_cp_element_group_52"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_core_CP_345_elements(9) & concat_core_CP_345_elements(95);
      gj_concat_core_cp_element_group_52 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_core_CP_345_elements(52), clk => clk, reset => reset); --
    end block;
    -- CP-element group 53:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	11 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (1) 
      -- CP-element group 53: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/phi_stmt_116_sample_start__ps
      -- 
    concat_core_CP_345_elements(53) <= concat_core_CP_345_elements(11);
    -- CP-element group 54:  join  transition  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	12 
    -- CP-element group 54:  members (1) 
      -- CP-element group 54: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/phi_stmt_116_sample_completed__ps
      -- 
    -- Element group concat_core_CP_345_elements(54) is bound as output of CP function.
    -- CP-element group 55:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	13 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (1) 
      -- CP-element group 55: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/phi_stmt_116_update_start__ps
      -- 
    concat_core_CP_345_elements(55) <= concat_core_CP_345_elements(13);
    -- CP-element group 56:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	14 
    -- CP-element group 56: 	93 
    -- CP-element group 56:  members (2) 
      -- CP-element group 56: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/phi_stmt_116_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/phi_stmt_116_update_completed__ps
      -- 
    -- Element group concat_core_CP_345_elements(56) is bound as output of CP function.
    -- CP-element group 57:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	7 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (1) 
      -- CP-element group 57: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/phi_stmt_116_loopback_trigger
      -- 
    concat_core_CP_345_elements(57) <= concat_core_CP_345_elements(7);
    -- CP-element group 58:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (2) 
      -- CP-element group 58: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/phi_stmt_116_loopback_sample_req
      -- CP-element group 58: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/phi_stmt_116_loopback_sample_req_ps
      -- 
    phi_stmt_116_loopback_sample_req_477_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_116_loopback_sample_req_477_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_core_CP_345_elements(58), ack => phi_stmt_116_req_1); -- 
    -- Element group concat_core_CP_345_elements(58) is bound as output of CP function.
    -- CP-element group 59:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	8 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/phi_stmt_116_entry_trigger
      -- 
    concat_core_CP_345_elements(59) <= concat_core_CP_345_elements(8);
    -- CP-element group 60:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: successors 
    -- CP-element group 60:  members (2) 
      -- CP-element group 60: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/phi_stmt_116_entry_sample_req
      -- CP-element group 60: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/phi_stmt_116_entry_sample_req_ps
      -- 
    phi_stmt_116_entry_sample_req_480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_116_entry_sample_req_480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_core_CP_345_elements(60), ack => phi_stmt_116_req_0); -- 
    -- Element group concat_core_CP_345_elements(60) is bound as output of CP function.
    -- CP-element group 61:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (2) 
      -- CP-element group 61: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/phi_stmt_116_phi_mux_ack
      -- CP-element group 61: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/phi_stmt_116_phi_mux_ack_ps
      -- 
    phi_stmt_116_phi_mux_ack_483_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_116_ack_0, ack => concat_core_CP_345_elements(61)); -- 
    -- CP-element group 62:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (4) 
      -- CP-element group 62: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_add_inp2_init_118_sample_start__ps
      -- CP-element group 62: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_add_inp2_init_118_sample_completed__ps
      -- CP-element group 62: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_add_inp2_init_118_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_add_inp2_init_118_sample_completed_
      -- 
    -- Element group concat_core_CP_345_elements(62) is bound as output of CP function.
    -- CP-element group 63:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	65 
    -- CP-element group 63:  members (2) 
      -- CP-element group 63: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_add_inp2_init_118_update_start__ps
      -- CP-element group 63: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_add_inp2_init_118_update_start_
      -- 
    -- Element group concat_core_CP_345_elements(63) is bound as output of CP function.
    -- CP-element group 64:  join  transition  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	65 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (1) 
      -- CP-element group 64: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_add_inp2_init_118_update_completed__ps
      -- 
    concat_core_CP_345_elements(64) <= concat_core_CP_345_elements(65);
    -- CP-element group 65:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	64 
    -- CP-element group 65:  members (1) 
      -- CP-element group 65: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_add_inp2_init_118_update_completed_
      -- 
    -- Element group concat_core_CP_345_elements(65) is a control-delay.
    cp_element_65_delay: control_delay_element  generic map(name => " 65_delay", delay_value => 1)  port map(req => concat_core_CP_345_elements(63), ack => concat_core_CP_345_elements(65), clk => clk, reset =>reset);
    -- CP-element group 66:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	68 
    -- CP-element group 66:  members (4) 
      -- CP-element group 66: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_next_add_inp2_119_sample_start__ps
      -- CP-element group 66: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_next_add_inp2_119_sample_start_
      -- CP-element group 66: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_next_add_inp2_119_Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_next_add_inp2_119_Sample/req
      -- 
    req_504_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_504_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_core_CP_345_elements(66), ack => next_add_inp2_192_119_buf_req_0); -- 
    -- Element group concat_core_CP_345_elements(66) is bound as output of CP function.
    -- CP-element group 67:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67:  members (4) 
      -- CP-element group 67: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_next_add_inp2_119_update_start__ps
      -- CP-element group 67: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_next_add_inp2_119_update_start_
      -- CP-element group 67: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_next_add_inp2_119_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_next_add_inp2_119_Update/req
      -- 
    req_509_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_509_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_core_CP_345_elements(67), ack => next_add_inp2_192_119_buf_req_1); -- 
    -- Element group concat_core_CP_345_elements(67) is bound as output of CP function.
    -- CP-element group 68:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (4) 
      -- CP-element group 68: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_next_add_inp2_119_sample_completed__ps
      -- CP-element group 68: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_next_add_inp2_119_sample_completed_
      -- CP-element group 68: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_next_add_inp2_119_Sample/$exit
      -- CP-element group 68: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_next_add_inp2_119_Sample/ack
      -- 
    ack_505_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_add_inp2_192_119_buf_ack_0, ack => concat_core_CP_345_elements(68)); -- 
    -- CP-element group 69:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	67 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (4) 
      -- CP-element group 69: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_next_add_inp2_119_update_completed__ps
      -- CP-element group 69: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_next_add_inp2_119_update_completed_
      -- CP-element group 69: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_next_add_inp2_119_Update/$exit
      -- CP-element group 69: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_next_add_inp2_119_Update/ack
      -- 
    ack_510_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_add_inp2_192_119_buf_ack_1, ack => concat_core_CP_345_elements(69)); -- 
    -- CP-element group 70:  join  transition  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	9 
    -- CP-element group 70: marked-predecessors 
    -- CP-element group 70: 	12 
    -- CP-element group 70: 	112 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	11 
    -- CP-element group 70:  members (1) 
      -- CP-element group 70: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/phi_stmt_120_sample_start_
      -- 
    concat_core_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
      constant joinName: string(1 to 31) := "concat_core_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_core_CP_345_elements(9) & concat_core_CP_345_elements(12) & concat_core_CP_345_elements(112);
      gj_concat_core_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_core_CP_345_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  join  transition  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	9 
    -- CP-element group 71: marked-predecessors 
    -- CP-element group 71: 	95 
    -- CP-element group 71: 	99 
    -- CP-element group 71: 	91 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	13 
    -- CP-element group 71:  members (1) 
      -- CP-element group 71: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/phi_stmt_120_update_start_
      -- 
    concat_core_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 31) := "concat_core_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= concat_core_CP_345_elements(9) & concat_core_CP_345_elements(95) & concat_core_CP_345_elements(99) & concat_core_CP_345_elements(91);
      gj_concat_core_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_core_CP_345_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	11 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/phi_stmt_120_sample_start__ps
      -- 
    concat_core_CP_345_elements(72) <= concat_core_CP_345_elements(11);
    -- CP-element group 73:  join  transition  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	12 
    -- CP-element group 73:  members (1) 
      -- CP-element group 73: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/phi_stmt_120_sample_completed__ps
      -- 
    -- Element group concat_core_CP_345_elements(73) is bound as output of CP function.
    -- CP-element group 74:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	13 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (1) 
      -- CP-element group 74: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/phi_stmt_120_update_start__ps
      -- 
    concat_core_CP_345_elements(74) <= concat_core_CP_345_elements(13);
    -- CP-element group 75:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	14 
    -- CP-element group 75: 	93 
    -- CP-element group 75: 	97 
    -- CP-element group 75: 	89 
    -- CP-element group 75:  members (2) 
      -- CP-element group 75: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/phi_stmt_120_update_completed_
      -- CP-element group 75: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/phi_stmt_120_update_completed__ps
      -- 
    -- Element group concat_core_CP_345_elements(75) is bound as output of CP function.
    -- CP-element group 76:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	7 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (1) 
      -- CP-element group 76: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/phi_stmt_120_loopback_trigger
      -- 
    concat_core_CP_345_elements(76) <= concat_core_CP_345_elements(7);
    -- CP-element group 77:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: successors 
    -- CP-element group 77:  members (2) 
      -- CP-element group 77: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/phi_stmt_120_loopback_sample_req
      -- CP-element group 77: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/phi_stmt_120_loopback_sample_req_ps
      -- 
    phi_stmt_120_loopback_sample_req_521_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_120_loopback_sample_req_521_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_core_CP_345_elements(77), ack => phi_stmt_120_req_1); -- 
    -- Element group concat_core_CP_345_elements(77) is bound as output of CP function.
    -- CP-element group 78:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	8 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/phi_stmt_120_entry_trigger
      -- 
    concat_core_CP_345_elements(78) <= concat_core_CP_345_elements(8);
    -- CP-element group 79:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/phi_stmt_120_entry_sample_req
      -- CP-element group 79: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/phi_stmt_120_entry_sample_req_ps
      -- 
    phi_stmt_120_entry_sample_req_524_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_120_entry_sample_req_524_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_core_CP_345_elements(79), ack => phi_stmt_120_req_0); -- 
    -- Element group concat_core_CP_345_elements(79) is bound as output of CP function.
    -- CP-element group 80:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (2) 
      -- CP-element group 80: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/phi_stmt_120_phi_mux_ack_ps
      -- CP-element group 80: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/phi_stmt_120_phi_mux_ack
      -- 
    phi_stmt_120_phi_mux_ack_527_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_120_ack_0, ack => concat_core_CP_345_elements(80)); -- 
    -- CP-element group 81:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: successors 
    -- CP-element group 81:  members (4) 
      -- CP-element group 81: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_count_inp1_init_122_sample_start_
      -- CP-element group 81: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_count_inp1_init_122_sample_completed__ps
      -- CP-element group 81: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_count_inp1_init_122_sample_start__ps
      -- CP-element group 81: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_count_inp1_init_122_sample_completed_
      -- 
    -- Element group concat_core_CP_345_elements(81) is bound as output of CP function.
    -- CP-element group 82:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	84 
    -- CP-element group 82:  members (2) 
      -- CP-element group 82: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_count_inp1_init_122_update_start__ps
      -- CP-element group 82: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_count_inp1_init_122_update_start_
      -- 
    -- Element group concat_core_CP_345_elements(82) is bound as output of CP function.
    -- CP-element group 83:  join  transition  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	84 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (1) 
      -- CP-element group 83: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_count_inp1_init_122_update_completed__ps
      -- 
    concat_core_CP_345_elements(83) <= concat_core_CP_345_elements(84);
    -- CP-element group 84:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	83 
    -- CP-element group 84:  members (1) 
      -- CP-element group 84: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_count_inp1_init_122_update_completed_
      -- 
    -- Element group concat_core_CP_345_elements(84) is a control-delay.
    cp_element_84_delay: control_delay_element  generic map(name => " 84_delay", delay_value => 1)  port map(req => concat_core_CP_345_elements(82), ack => concat_core_CP_345_elements(84), clk => clk, reset =>reset);
    -- CP-element group 85:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (4) 
      -- CP-element group 85: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_next_count_inp1_123_sample_start__ps
      -- CP-element group 85: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_next_count_inp1_123_Sample/req
      -- CP-element group 85: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_next_count_inp1_123_Sample/$entry
      -- CP-element group 85: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_next_count_inp1_123_sample_start_
      -- 
    req_548_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_548_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_core_CP_345_elements(85), ack => next_count_inp1_176_123_buf_req_0); -- 
    -- Element group concat_core_CP_345_elements(85) is bound as output of CP function.
    -- CP-element group 86:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	88 
    -- CP-element group 86:  members (4) 
      -- CP-element group 86: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_next_count_inp1_123_update_start__ps
      -- CP-element group 86: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_next_count_inp1_123_Update/req
      -- CP-element group 86: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_next_count_inp1_123_Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_next_count_inp1_123_update_start_
      -- 
    req_553_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_553_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_core_CP_345_elements(86), ack => next_count_inp1_176_123_buf_req_1); -- 
    -- Element group concat_core_CP_345_elements(86) is bound as output of CP function.
    -- CP-element group 87:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: successors 
    -- CP-element group 87:  members (4) 
      -- CP-element group 87: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_next_count_inp1_123_sample_completed__ps
      -- CP-element group 87: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_next_count_inp1_123_Sample/ack
      -- CP-element group 87: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_next_count_inp1_123_Sample/$exit
      -- CP-element group 87: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_next_count_inp1_123_sample_completed_
      -- 
    ack_549_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_count_inp1_176_123_buf_ack_0, ack => concat_core_CP_345_elements(87)); -- 
    -- CP-element group 88:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	86 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (4) 
      -- CP-element group 88: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_next_count_inp1_123_Update/ack
      -- CP-element group 88: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_next_count_inp1_123_Update/$exit
      -- CP-element group 88: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_next_count_inp1_123_update_completed_
      -- CP-element group 88: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/R_next_count_inp1_123_update_completed__ps
      -- 
    ack_554_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => next_count_inp1_176_123_buf_ack_1, ack => concat_core_CP_345_elements(88)); -- 
    -- CP-element group 89:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	37 
    -- CP-element group 89: 	75 
    -- CP-element group 89: marked-predecessors 
    -- CP-element group 89: 	91 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/call_stmt_135_Sample/crr
      -- CP-element group 89: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/call_stmt_135_Sample/$entry
      -- CP-element group 89: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/call_stmt_135_sample_start_
      -- 
    crr_563_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_563_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_core_CP_345_elements(89), ack => call_stmt_135_call_req_0); -- 
    concat_core_cp_element_group_89: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 31) := "concat_core_cp_element_group_89"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_core_CP_345_elements(37) & concat_core_CP_345_elements(75) & concat_core_CP_345_elements(91);
      gj_concat_core_cp_element_group_89 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_core_CP_345_elements(89), clk => clk, reset => reset); --
    end block;
    -- CP-element group 90:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: marked-predecessors 
    -- CP-element group 90: 	107 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	92 
    -- CP-element group 90:  members (3) 
      -- CP-element group 90: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/call_stmt_135_Update/ccr
      -- CP-element group 90: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/call_stmt_135_Update/$entry
      -- CP-element group 90: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/call_stmt_135_update_start_
      -- 
    ccr_568_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_568_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_core_CP_345_elements(90), ack => call_stmt_135_call_req_1); -- 
    concat_core_cp_element_group_90: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "concat_core_cp_element_group_90"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= concat_core_CP_345_elements(107);
      gj_concat_core_cp_element_group_90 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_core_CP_345_elements(90), clk => clk, reset => reset); --
    end block;
    -- CP-element group 91:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: successors 
    -- CP-element group 91: marked-successors 
    -- CP-element group 91: 	33 
    -- CP-element group 91: 	71 
    -- CP-element group 91: 	89 
    -- CP-element group 91:  members (3) 
      -- CP-element group 91: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/call_stmt_135_Sample/cra
      -- CP-element group 91: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/call_stmt_135_Sample/$exit
      -- CP-element group 91: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/call_stmt_135_sample_completed_
      -- 
    cra_564_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_135_call_ack_0, ack => concat_core_CP_345_elements(91)); -- 
    -- CP-element group 92:  transition  input  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	90 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	105 
    -- CP-element group 92:  members (3) 
      -- CP-element group 92: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/call_stmt_135_Update/cca
      -- CP-element group 92: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/call_stmt_135_Update/$exit
      -- CP-element group 92: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/call_stmt_135_update_completed_
      -- 
    cca_569_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_135_call_ack_1, ack => concat_core_CP_345_elements(92)); -- 
    -- CP-element group 93:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	56 
    -- CP-element group 93: 	75 
    -- CP-element group 93: marked-predecessors 
    -- CP-element group 93: 	95 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/call_stmt_141_sample_start_
      -- CP-element group 93: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/call_stmt_141_Sample/crr
      -- CP-element group 93: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/call_stmt_141_Sample/$entry
      -- 
    crr_577_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_577_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_core_CP_345_elements(93), ack => call_stmt_141_call_req_0); -- 
    concat_core_cp_element_group_93: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 31) := "concat_core_cp_element_group_93"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= concat_core_CP_345_elements(56) & concat_core_CP_345_elements(75) & concat_core_CP_345_elements(95);
      gj_concat_core_cp_element_group_93 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_core_CP_345_elements(93), clk => clk, reset => reset); --
    end block;
    -- CP-element group 94:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: marked-predecessors 
    -- CP-element group 94: 	107 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	96 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/call_stmt_141_update_start_
      -- CP-element group 94: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/call_stmt_141_Update/ccr
      -- CP-element group 94: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/call_stmt_141_Update/$entry
      -- 
    ccr_582_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_582_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_core_CP_345_elements(94), ack => call_stmt_141_call_req_1); -- 
    concat_core_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "concat_core_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= concat_core_CP_345_elements(107);
      gj_concat_core_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_core_CP_345_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: successors 
    -- CP-element group 95: marked-successors 
    -- CP-element group 95: 	52 
    -- CP-element group 95: 	93 
    -- CP-element group 95: 	71 
    -- CP-element group 95:  members (3) 
      -- CP-element group 95: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/call_stmt_141_sample_completed_
      -- CP-element group 95: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/call_stmt_141_Sample/cra
      -- CP-element group 95: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/call_stmt_141_Sample/$exit
      -- 
    cra_578_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_141_call_ack_0, ack => concat_core_CP_345_elements(95)); -- 
    -- CP-element group 96:  transition  input  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	94 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	105 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/call_stmt_141_update_completed_
      -- CP-element group 96: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/call_stmt_141_Update/cca
      -- CP-element group 96: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/call_stmt_141_Update/$exit
      -- 
    cca_583_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_141_call_ack_1, ack => concat_core_CP_345_elements(96)); -- 
    -- CP-element group 97:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	75 
    -- CP-element group 97: marked-predecessors 
    -- CP-element group 97: 	99 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	99 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/assign_stmt_144_Sample/req
      -- CP-element group 97: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/assign_stmt_144_Sample/$entry
      -- CP-element group 97: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/assign_stmt_144_sample_start_
      -- 
    req_591_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_591_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_core_CP_345_elements(97), ack => W_cmp_143_delayed_15_0_142_inst_req_0); -- 
    concat_core_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "concat_core_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_core_CP_345_elements(75) & concat_core_CP_345_elements(99);
      gj_concat_core_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_core_CP_345_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: marked-predecessors 
    -- CP-element group 98: 	107 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	100 
    -- CP-element group 98:  members (3) 
      -- CP-element group 98: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/assign_stmt_144_update_start_
      -- CP-element group 98: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/assign_stmt_144_Update/req
      -- CP-element group 98: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/assign_stmt_144_Update/$entry
      -- 
    req_596_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_596_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_core_CP_345_elements(98), ack => W_cmp_143_delayed_15_0_142_inst_req_1); -- 
    concat_core_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "concat_core_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= concat_core_CP_345_elements(107);
      gj_concat_core_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_core_CP_345_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	97 
    -- CP-element group 99: successors 
    -- CP-element group 99: marked-successors 
    -- CP-element group 99: 	97 
    -- CP-element group 99: 	71 
    -- CP-element group 99:  members (3) 
      -- CP-element group 99: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/assign_stmt_144_Sample/ack
      -- CP-element group 99: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/assign_stmt_144_Sample/$exit
      -- CP-element group 99: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/assign_stmt_144_sample_completed_
      -- 
    ack_592_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_cmp_143_delayed_15_0_142_inst_ack_0, ack => concat_core_CP_345_elements(99)); -- 
    -- CP-element group 100:  transition  input  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	98 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	105 
    -- CP-element group 100:  members (3) 
      -- CP-element group 100: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/assign_stmt_144_update_completed_
      -- CP-element group 100: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/assign_stmt_144_Update/ack
      -- CP-element group 100: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/assign_stmt_144_Update/$exit
      -- 
    ack_597_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_cmp_143_delayed_15_0_142_inst_ack_1, ack => concat_core_CP_345_elements(100)); -- 
    -- CP-element group 101:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	18 
    -- CP-element group 101: marked-predecessors 
    -- CP-element group 101: 	103 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	103 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/assign_stmt_153_Sample/req
      -- CP-element group 101: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/assign_stmt_153_Sample/$entry
      -- CP-element group 101: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/assign_stmt_153_sample_start_
      -- 
    req_605_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_605_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_core_CP_345_elements(101), ack => W_add_out_149_delayed_15_0_151_inst_req_0); -- 
    concat_core_cp_element_group_101: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 32) := "concat_core_cp_element_group_101"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_core_CP_345_elements(18) & concat_core_CP_345_elements(103);
      gj_concat_core_cp_element_group_101 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_core_CP_345_elements(101), clk => clk, reset => reset); --
    end block;
    -- CP-element group 102:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: marked-predecessors 
    -- CP-element group 102: 	107 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	104 
    -- CP-element group 102:  members (3) 
      -- CP-element group 102: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/assign_stmt_153_Update/req
      -- CP-element group 102: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/assign_stmt_153_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/assign_stmt_153_update_start_
      -- 
    req_610_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_610_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_core_CP_345_elements(102), ack => W_add_out_149_delayed_15_0_151_inst_req_1); -- 
    concat_core_cp_element_group_102: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 32) := "concat_core_cp_element_group_102"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= concat_core_CP_345_elements(107);
      gj_concat_core_cp_element_group_102 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_core_CP_345_elements(102), clk => clk, reset => reset); --
    end block;
    -- CP-element group 103:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	101 
    -- CP-element group 103: successors 
    -- CP-element group 103: marked-successors 
    -- CP-element group 103: 	16 
    -- CP-element group 103: 	101 
    -- CP-element group 103:  members (3) 
      -- CP-element group 103: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/assign_stmt_153_Sample/ack
      -- CP-element group 103: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/assign_stmt_153_Sample/$exit
      -- CP-element group 103: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/assign_stmt_153_sample_completed_
      -- 
    ack_606_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_add_out_149_delayed_15_0_151_inst_ack_0, ack => concat_core_CP_345_elements(103)); -- 
    -- CP-element group 104:  transition  input  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	102 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	105 
    -- CP-element group 104:  members (3) 
      -- CP-element group 104: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/assign_stmt_153_Update/ack
      -- CP-element group 104: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/assign_stmt_153_Update/$exit
      -- CP-element group 104: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/assign_stmt_153_update_completed_
      -- 
    ack_611_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_add_out_149_delayed_15_0_151_inst_ack_1, ack => concat_core_CP_345_elements(104)); -- 
    -- CP-element group 105:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	92 
    -- CP-element group 105: 	96 
    -- CP-element group 105: 	100 
    -- CP-element group 105: 	104 
    -- CP-element group 105: marked-predecessors 
    -- CP-element group 105: 	107 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	107 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/call_stmt_158_Sample/crr
      -- CP-element group 105: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/call_stmt_158_Sample/$entry
      -- CP-element group 105: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/call_stmt_158_sample_start_
      -- 
    crr_619_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_619_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_core_CP_345_elements(105), ack => call_stmt_158_call_req_0); -- 
    concat_core_cp_element_group_105: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 32) := "concat_core_cp_element_group_105"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= concat_core_CP_345_elements(92) & concat_core_CP_345_elements(96) & concat_core_CP_345_elements(100) & concat_core_CP_345_elements(104) & concat_core_CP_345_elements(107);
      gj_concat_core_cp_element_group_105 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_core_CP_345_elements(105), clk => clk, reset => reset); --
    end block;
    -- CP-element group 106:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: marked-predecessors 
    -- CP-element group 106: 	108 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	108 
    -- CP-element group 106:  members (3) 
      -- CP-element group 106: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/call_stmt_158_update_start_
      -- CP-element group 106: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/call_stmt_158_Update/ccr
      -- CP-element group 106: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/call_stmt_158_Update/$entry
      -- 
    ccr_624_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_624_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_core_CP_345_elements(106), ack => call_stmt_158_call_req_1); -- 
    concat_core_cp_element_group_106: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 32) := "concat_core_cp_element_group_106"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= concat_core_CP_345_elements(108);
      gj_concat_core_cp_element_group_106 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_core_CP_345_elements(106), clk => clk, reset => reset); --
    end block;
    -- CP-element group 107:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	105 
    -- CP-element group 107: successors 
    -- CP-element group 107: marked-successors 
    -- CP-element group 107: 	94 
    -- CP-element group 107: 	98 
    -- CP-element group 107: 	102 
    -- CP-element group 107: 	105 
    -- CP-element group 107: 	90 
    -- CP-element group 107:  members (3) 
      -- CP-element group 107: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/call_stmt_158_Sample/cra
      -- CP-element group 107: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/call_stmt_158_Sample/$exit
      -- CP-element group 107: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/call_stmt_158_sample_completed_
      -- 
    cra_620_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_158_call_ack_0, ack => concat_core_CP_345_elements(107)); -- 
    -- CP-element group 108:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	106 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	118 
    -- CP-element group 108: marked-successors 
    -- CP-element group 108: 	106 
    -- CP-element group 108:  members (3) 
      -- CP-element group 108: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/call_stmt_158_Update/cca
      -- CP-element group 108: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/call_stmt_158_update_completed_
      -- CP-element group 108: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/call_stmt_158_Update/$exit
      -- 
    cca_625_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_158_call_ack_1, ack => concat_core_CP_345_elements(108)); -- 
    -- CP-element group 109:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	9 
    -- CP-element group 109: marked-predecessors 
    -- CP-element group 109: 	111 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/SUB_u16_u16_162_sample_start_
      -- CP-element group 109: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/SUB_u16_u16_162_Sample/rr
      -- CP-element group 109: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/SUB_u16_u16_162_Sample/$entry
      -- 
    rr_633_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_633_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_core_CP_345_elements(109), ack => SUB_u16_u16_162_inst_req_0); -- 
    concat_core_cp_element_group_109: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 32) := "concat_core_cp_element_group_109"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_core_CP_345_elements(9) & concat_core_CP_345_elements(111);
      gj_concat_core_cp_element_group_109 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_core_CP_345_elements(109), clk => clk, reset => reset); --
    end block;
    -- CP-element group 110:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	12 
    -- CP-element group 110: marked-predecessors 
    -- CP-element group 110: 	112 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	112 
    -- CP-element group 110:  members (3) 
      -- CP-element group 110: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/SUB_u16_u16_162_update_start_
      -- CP-element group 110: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/SUB_u16_u16_162_Update/cr
      -- CP-element group 110: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/SUB_u16_u16_162_Update/$entry
      -- 
    cr_638_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_638_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_core_CP_345_elements(110), ack => SUB_u16_u16_162_inst_req_1); -- 
    concat_core_cp_element_group_110: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "concat_core_cp_element_group_110"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_core_CP_345_elements(12) & concat_core_CP_345_elements(112);
      gj_concat_core_cp_element_group_110 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_core_CP_345_elements(110), clk => clk, reset => reset); --
    end block;
    -- CP-element group 111:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: successors 
    -- CP-element group 111: marked-successors 
    -- CP-element group 111: 	109 
    -- CP-element group 111:  members (3) 
      -- CP-element group 111: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/SUB_u16_u16_162_sample_completed_
      -- CP-element group 111: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/SUB_u16_u16_162_Sample/ra
      -- CP-element group 111: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/SUB_u16_u16_162_Sample/$exit
      -- 
    ra_634_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_162_inst_ack_0, ack => concat_core_CP_345_elements(111)); -- 
    -- CP-element group 112:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	110 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	10 
    -- CP-element group 112: marked-successors 
    -- CP-element group 112: 	110 
    -- CP-element group 112: 	70 
    -- CP-element group 112:  members (3) 
      -- CP-element group 112: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/SUB_u16_u16_162_update_completed_
      -- CP-element group 112: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/SUB_u16_u16_162_Update/ca
      -- CP-element group 112: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/SUB_u16_u16_162_Update/$exit
      -- 
    ca_639_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_162_inst_ack_1, ack => concat_core_CP_345_elements(112)); -- 
    -- CP-element group 113:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	9 
    -- CP-element group 113: marked-predecessors 
    -- CP-element group 113: 	115 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/SUB_u32_u32_201_Sample/rr
      -- CP-element group 113: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/SUB_u32_u32_201_Sample/$entry
      -- CP-element group 113: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/SUB_u32_u32_201_sample_start_
      -- 
    rr_647_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_647_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_core_CP_345_elements(113), ack => SUB_u32_u32_201_inst_req_0); -- 
    concat_core_cp_element_group_113: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 32) := "concat_core_cp_element_group_113"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_core_CP_345_elements(9) & concat_core_CP_345_elements(115);
      gj_concat_core_cp_element_group_113 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_core_CP_345_elements(113), clk => clk, reset => reset); --
    end block;
    -- CP-element group 114:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: marked-predecessors 
    -- CP-element group 114: 	116 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	116 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/SUB_u32_u32_201_update_start_
      -- CP-element group 114: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/SUB_u32_u32_201_Update/cr
      -- CP-element group 114: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/SUB_u32_u32_201_Update/$entry
      -- 
    cr_652_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_652_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => concat_core_CP_345_elements(114), ack => SUB_u32_u32_201_inst_req_1); -- 
    concat_core_cp_element_group_114: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 32) := "concat_core_cp_element_group_114"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= concat_core_CP_345_elements(116);
      gj_concat_core_cp_element_group_114 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_core_CP_345_elements(114), clk => clk, reset => reset); --
    end block;
    -- CP-element group 115:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: successors 
    -- CP-element group 115: marked-successors 
    -- CP-element group 115: 	113 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/SUB_u32_u32_201_Sample/$exit
      -- CP-element group 115: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/SUB_u32_u32_201_sample_completed_
      -- CP-element group 115: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/SUB_u32_u32_201_Sample/ra
      -- 
    ra_648_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u32_u32_201_inst_ack_0, ack => concat_core_CP_345_elements(115)); -- 
    -- CP-element group 116:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	114 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	10 
    -- CP-element group 116: marked-successors 
    -- CP-element group 116: 	114 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/SUB_u32_u32_201_update_completed_
      -- CP-element group 116: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/SUB_u32_u32_201_Update/ca
      -- CP-element group 116: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/SUB_u32_u32_201_Update/$exit
      -- 
    ca_653_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u32_u32_201_inst_ack_1, ack => concat_core_CP_345_elements(116)); -- 
    -- CP-element group 117:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	9 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	10 
    -- CP-element group 117:  members (1) 
      -- CP-element group 117: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group concat_core_CP_345_elements(117) is a control-delay.
    cp_element_117_delay: control_delay_element  generic map(name => " 117_delay", delay_value => 1)  port map(req => concat_core_CP_345_elements(9), ack => concat_core_CP_345_elements(117), clk => clk, reset =>reset);
    -- CP-element group 118:  join  transition  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	12 
    -- CP-element group 118: 	108 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	6 
    -- CP-element group 118:  members (1) 
      -- CP-element group 118: 	 branch_block_stmt_69/do_while_stmt_106/do_while_stmt_106_loop_body/$exit
      -- 
    concat_core_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "concat_core_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= concat_core_CP_345_elements(12) & concat_core_CP_345_elements(108);
      gj_concat_core_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => concat_core_CP_345_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  transition  input  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	5 
    -- CP-element group 119: successors 
    -- CP-element group 119:  members (2) 
      -- CP-element group 119: 	 branch_block_stmt_69/do_while_stmt_106/loop_exit/ack
      -- CP-element group 119: 	 branch_block_stmt_69/do_while_stmt_106/loop_exit/$exit
      -- 
    ack_658_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_106_branch_ack_0, ack => concat_core_CP_345_elements(119)); -- 
    -- CP-element group 120:  transition  input  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	5 
    -- CP-element group 120: successors 
    -- CP-element group 120:  members (2) 
      -- CP-element group 120: 	 branch_block_stmt_69/do_while_stmt_106/loop_taken/ack
      -- CP-element group 120: 	 branch_block_stmt_69/do_while_stmt_106/loop_taken/$exit
      -- 
    ack_662_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_106_branch_ack_1, ack => concat_core_CP_345_elements(120)); -- 
    -- CP-element group 121:  transition  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	3 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	1 
    -- CP-element group 121:  members (1) 
      -- CP-element group 121: 	 branch_block_stmt_69/do_while_stmt_106/$exit
      -- 
    concat_core_CP_345_elements(121) <= concat_core_CP_345_elements(3);
    concat_core_do_while_stmt_106_terminator_663: loop_terminator -- 
      generic map (name => " concat_core_do_while_stmt_106_terminator_663", max_iterations_in_flight =>15) 
      port map(loop_body_exit => concat_core_CP_345_elements(6),loop_continue => concat_core_CP_345_elements(120),loop_terminate => concat_core_CP_345_elements(119),loop_back => concat_core_CP_345_elements(4),loop_exit => concat_core_CP_345_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_108_phi_seq_423_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= concat_core_CP_345_elements(21);
      concat_core_CP_345_elements(24)<= src_sample_reqs(0);
      src_sample_acks(0)  <= concat_core_CP_345_elements(24);
      concat_core_CP_345_elements(25)<= src_update_reqs(0);
      src_update_acks(0)  <= concat_core_CP_345_elements(26);
      concat_core_CP_345_elements(22) <= phi_mux_reqs(0);
      triggers(1)  <= concat_core_CP_345_elements(19);
      concat_core_CP_345_elements(28)<= src_sample_reqs(1);
      src_sample_acks(1)  <= concat_core_CP_345_elements(30);
      concat_core_CP_345_elements(29)<= src_update_reqs(1);
      src_update_acks(1)  <= concat_core_CP_345_elements(31);
      concat_core_CP_345_elements(20) <= phi_mux_reqs(1);
      phi_stmt_108_phi_seq_423 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_108_phi_seq_423") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => concat_core_CP_345_elements(11), 
          phi_sample_ack => concat_core_CP_345_elements(17), 
          phi_update_req => concat_core_CP_345_elements(13), 
          phi_update_ack => concat_core_CP_345_elements(18), 
          phi_mux_ack => concat_core_CP_345_elements(23), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_112_phi_seq_467_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= concat_core_CP_345_elements(40);
      concat_core_CP_345_elements(43)<= src_sample_reqs(0);
      src_sample_acks(0)  <= concat_core_CP_345_elements(43);
      concat_core_CP_345_elements(44)<= src_update_reqs(0);
      src_update_acks(0)  <= concat_core_CP_345_elements(45);
      concat_core_CP_345_elements(41) <= phi_mux_reqs(0);
      triggers(1)  <= concat_core_CP_345_elements(38);
      concat_core_CP_345_elements(47)<= src_sample_reqs(1);
      src_sample_acks(1)  <= concat_core_CP_345_elements(49);
      concat_core_CP_345_elements(48)<= src_update_reqs(1);
      src_update_acks(1)  <= concat_core_CP_345_elements(50);
      concat_core_CP_345_elements(39) <= phi_mux_reqs(1);
      phi_stmt_112_phi_seq_467 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_112_phi_seq_467") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => concat_core_CP_345_elements(34), 
          phi_sample_ack => concat_core_CP_345_elements(35), 
          phi_update_req => concat_core_CP_345_elements(36), 
          phi_update_ack => concat_core_CP_345_elements(37), 
          phi_mux_ack => concat_core_CP_345_elements(42), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_116_phi_seq_511_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= concat_core_CP_345_elements(59);
      concat_core_CP_345_elements(62)<= src_sample_reqs(0);
      src_sample_acks(0)  <= concat_core_CP_345_elements(62);
      concat_core_CP_345_elements(63)<= src_update_reqs(0);
      src_update_acks(0)  <= concat_core_CP_345_elements(64);
      concat_core_CP_345_elements(60) <= phi_mux_reqs(0);
      triggers(1)  <= concat_core_CP_345_elements(57);
      concat_core_CP_345_elements(66)<= src_sample_reqs(1);
      src_sample_acks(1)  <= concat_core_CP_345_elements(68);
      concat_core_CP_345_elements(67)<= src_update_reqs(1);
      src_update_acks(1)  <= concat_core_CP_345_elements(69);
      concat_core_CP_345_elements(58) <= phi_mux_reqs(1);
      phi_stmt_116_phi_seq_511 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_116_phi_seq_511") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => concat_core_CP_345_elements(53), 
          phi_sample_ack => concat_core_CP_345_elements(54), 
          phi_update_req => concat_core_CP_345_elements(55), 
          phi_update_ack => concat_core_CP_345_elements(56), 
          phi_mux_ack => concat_core_CP_345_elements(61), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_120_phi_seq_555_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= concat_core_CP_345_elements(78);
      concat_core_CP_345_elements(81)<= src_sample_reqs(0);
      src_sample_acks(0)  <= concat_core_CP_345_elements(81);
      concat_core_CP_345_elements(82)<= src_update_reqs(0);
      src_update_acks(0)  <= concat_core_CP_345_elements(83);
      concat_core_CP_345_elements(79) <= phi_mux_reqs(0);
      triggers(1)  <= concat_core_CP_345_elements(76);
      concat_core_CP_345_elements(85)<= src_sample_reqs(1);
      src_sample_acks(1)  <= concat_core_CP_345_elements(87);
      concat_core_CP_345_elements(86)<= src_update_reqs(1);
      src_update_acks(1)  <= concat_core_CP_345_elements(88);
      concat_core_CP_345_elements(77) <= phi_mux_reqs(1);
      phi_stmt_120_phi_seq_555 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_120_phi_seq_555") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => concat_core_CP_345_elements(72), 
          phi_sample_ack => concat_core_CP_345_elements(73), 
          phi_update_req => concat_core_CP_345_elements(74), 
          phi_update_ack => concat_core_CP_345_elements(75), 
          phi_mux_ack => concat_core_CP_345_elements(80), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_375_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= concat_core_CP_345_elements(7);
        preds(1)  <= concat_core_CP_345_elements(8);
        entry_tmerge_375 : transition_merge -- 
          generic map(name => " entry_tmerge_375")
          port map (preds => preds, symbol_out => concat_core_CP_345_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u16_u16_174_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_181_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_190_wire : std_logic_vector(15 downto 0);
    signal NOT_u1_u1_205_wire : std_logic_vector(0 downto 0);
    signal SUB_u16_u16_157_157_delayed_1_0_163 : std_logic_vector(15 downto 0);
    signal SUB_u32_u32_195_195_delayed_1_0_202 : std_logic_vector(31 downto 0);
    signal ULT_u32_u1_208_wire : std_logic_vector(0 downto 0);
    signal add_inp1_112 : std_logic_vector(15 downto 0);
    signal add_inp1_init_92 : std_logic_vector(15 downto 0);
    signal add_inp2_116 : std_logic_vector(15 downto 0);
    signal add_inp2_init_96 : std_logic_vector(15 downto 0);
    signal add_out_108 : std_logic_vector(31 downto 0);
    signal add_out_149_delayed_15_0_153 : std_logic_vector(31 downto 0);
    signal add_out_init_88 : std_logic_vector(31 downto 0);
    signal cmp_129 : std_logic_vector(0 downto 0);
    signal cmp_143_delayed_15_0_144 : std_logic_vector(0 downto 0);
    signal continue_flag_210 : std_logic_vector(0 downto 0);
    signal count_inp1_120 : std_logic_vector(15 downto 0);
    signal count_inp1_init_100 : std_logic_vector(15 downto 0);
    signal done_158 : std_logic_vector(0 downto 0);
    signal i1_135 : std_logic_vector(63 downto 0);
    signal i2_141 : std_logic_vector(63 downto 0);
    signal index1_72 : std_logic_vector(7 downto 0);
    signal index2_75 : std_logic_vector(7 downto 0);
    signal index3_78 : std_logic_vector(7 downto 0);
    signal konst_161_wire_constant : std_logic_vector(15 downto 0);
    signal konst_171_wire_constant : std_logic_vector(15 downto 0);
    signal konst_173_wire_constant : std_logic_vector(15 downto 0);
    signal konst_180_wire_constant : std_logic_vector(15 downto 0);
    signal konst_189_wire_constant : std_logic_vector(15 downto 0);
    signal konst_195_wire_constant : std_logic_vector(31 downto 0);
    signal konst_200_wire_constant : std_logic_vector(31 downto 0);
    signal my_flag_168 : std_logic_vector(0 downto 0);
    signal next_add_inp1_184 : std_logic_vector(15 downto 0);
    signal next_add_inp1_184_115_buffered : std_logic_vector(15 downto 0);
    signal next_add_inp2_192 : std_logic_vector(15 downto 0);
    signal next_add_inp2_192_119_buffered : std_logic_vector(15 downto 0);
    signal next_add_out_197 : std_logic_vector(31 downto 0);
    signal next_add_out_197_111_buffered : std_logic_vector(31 downto 0);
    signal next_count_inp1_176 : std_logic_vector(15 downto 0);
    signal next_count_inp1_176_123_buffered : std_logic_vector(15 downto 0);
    signal o_150 : std_logic_vector(63 downto 0);
    signal out_concat_84 : std_logic_vector(31 downto 0);
    signal total_size_105 : std_logic_vector(15 downto 0);
    signal type_cast_133_wire : std_logic_vector(31 downto 0);
    signal type_cast_139_wire : std_logic_vector(31 downto 0);
    signal type_cast_82_wire_constant : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    add_inp1_init_92 <= "0000000000000000";
    add_inp2_init_96 <= "0000000000000000";
    add_out_init_88 <= "00000000000000000000000000000000";
    count_inp1_init_100 <= "0000000000000000";
    index1_72 <= "00000000";
    index2_75 <= "00000001";
    index3_78 <= "00000010";
    konst_161_wire_constant <= "0000000000000001";
    konst_171_wire_constant <= "0000000000000000";
    konst_173_wire_constant <= "0000000000000001";
    konst_180_wire_constant <= "0000000000000001";
    konst_189_wire_constant <= "0000000000000001";
    konst_195_wire_constant <= "00000000000000000000000000000001";
    konst_200_wire_constant <= "00000000000000000000000000000001";
    type_cast_82_wire_constant <= "00000000000000000000000000000011";
    phi_stmt_108: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= add_out_init_88 & next_add_out_197_111_buffered;
      req <= phi_stmt_108_req_0 & phi_stmt_108_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_108",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_108_ack_0,
          idata => idata,
          odata => add_out_108,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_108
    phi_stmt_112: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= add_inp1_init_92 & next_add_inp1_184_115_buffered;
      req <= phi_stmt_112_req_0 & phi_stmt_112_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_112",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_112_ack_0,
          idata => idata,
          odata => add_inp1_112,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_112
    phi_stmt_116: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= add_inp2_init_96 & next_add_inp2_192_119_buffered;
      req <= phi_stmt_116_req_0 & phi_stmt_116_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_116",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_116_ack_0,
          idata => idata,
          odata => add_inp2_116,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_116
    phi_stmt_120: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= count_inp1_init_100 & next_count_inp1_176_123_buffered;
      req <= phi_stmt_120_req_0 & phi_stmt_120_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_120",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_120_ack_0,
          idata => idata,
          odata => count_inp1_120,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_120
    -- flow-through select operator MUX_149_inst
    o_150 <= i1_135 when (cmp_143_delayed_15_0_144(0) /=  '0') else i2_141;
    -- flow-through select operator MUX_175_inst
    next_count_inp1_176 <= konst_171_wire_constant when (my_flag_168(0) /=  '0') else ADD_u16_u16_174_wire;
    -- flow-through select operator MUX_183_inst
    next_add_inp1_184 <= ADD_u16_u16_181_wire when (cmp_129(0) /=  '0') else add_inp1_112;
    -- flow-through select operator MUX_191_inst
    next_add_inp2_192 <= add_inp2_116 when (cmp_129(0) /=  '0') else ADD_u16_u16_190_wire;
    W_add_out_149_delayed_15_0_151_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_add_out_149_delayed_15_0_151_inst_req_0;
      W_add_out_149_delayed_15_0_151_inst_ack_0<= wack(0);
      rreq(0) <= W_add_out_149_delayed_15_0_151_inst_req_1;
      W_add_out_149_delayed_15_0_151_inst_ack_1<= rack(0);
      W_add_out_149_delayed_15_0_151_inst : InterlockBuffer generic map ( -- 
        name => "W_add_out_149_delayed_15_0_151_inst",
        buffer_size => 15,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add_out_108,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => add_out_149_delayed_15_0_153,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_cmp_143_delayed_15_0_142_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_cmp_143_delayed_15_0_142_inst_req_0;
      W_cmp_143_delayed_15_0_142_inst_ack_0<= wack(0);
      rreq(0) <= W_cmp_143_delayed_15_0_142_inst_req_1;
      W_cmp_143_delayed_15_0_142_inst_ack_1<= rack(0);
      W_cmp_143_delayed_15_0_142_inst : InterlockBuffer generic map ( -- 
        name => "W_cmp_143_delayed_15_0_142_inst",
        buffer_size => 15,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp_129,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => cmp_143_delayed_15_0_144,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_add_inp1_184_115_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_add_inp1_184_115_buf_req_0;
      next_add_inp1_184_115_buf_ack_0<= wack(0);
      rreq(0) <= next_add_inp1_184_115_buf_req_1;
      next_add_inp1_184_115_buf_ack_1<= rack(0);
      next_add_inp1_184_115_buf : InterlockBuffer generic map ( -- 
        name => "next_add_inp1_184_115_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_add_inp1_184,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_add_inp1_184_115_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_add_inp2_192_119_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_add_inp2_192_119_buf_req_0;
      next_add_inp2_192_119_buf_ack_0<= wack(0);
      rreq(0) <= next_add_inp2_192_119_buf_req_1;
      next_add_inp2_192_119_buf_ack_1<= rack(0);
      next_add_inp2_192_119_buf : InterlockBuffer generic map ( -- 
        name => "next_add_inp2_192_119_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_add_inp2_192,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_add_inp2_192_119_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_add_out_197_111_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_add_out_197_111_buf_req_0;
      next_add_out_197_111_buf_ack_0<= wack(0);
      rreq(0) <= next_add_out_197_111_buf_req_1;
      next_add_out_197_111_buf_ack_1<= rack(0);
      next_add_out_197_111_buf : InterlockBuffer generic map ( -- 
        name => "next_add_out_197_111_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_add_out_197,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_add_out_197_111_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    next_count_inp1_176_123_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= next_count_inp1_176_123_buf_req_0;
      next_count_inp1_176_123_buf_ack_0<= wack(0);
      rreq(0) <= next_count_inp1_176_123_buf_req_1;
      next_count_inp1_176_123_buf_ack_1<= rack(0);
      next_count_inp1_176_123_buf : InterlockBuffer generic map ( -- 
        name => "next_count_inp1_176_123_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_count_inp1_176,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_count_inp1_176_123_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_133_inst
    process(add_inp1_112) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := add_inp1_112(15 downto 0);
      type_cast_133_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_139_inst
    process(add_inp2_116) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := add_inp2_116(15 downto 0);
      type_cast_139_wire <= tmp_var; -- 
    end process;
    do_while_stmt_106_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= continue_flag_210;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_106_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_106_branch_req_0,
          ack0 => do_while_stmt_106_branch_ack_0,
          ack1 => do_while_stmt_106_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_104_inst
    process(input1_count_buffer, input2_count_buffer) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input1_count_buffer, input2_count_buffer, tmp_var);
      total_size_105 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_174_inst
    process(count_inp1_120) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(count_inp1_120, konst_173_wire_constant, tmp_var);
      ADD_u16_u16_174_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_181_inst
    process(add_inp1_112) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_inp1_112, konst_180_wire_constant, tmp_var);
      ADD_u16_u16_181_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_190_inst
    process(add_inp2_116) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_inp2_116, konst_189_wire_constant, tmp_var);
      ADD_u16_u16_190_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_196_inst
    process(add_out_108) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add_out_108, konst_195_wire_constant, tmp_var);
      next_add_out_197 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_167_inst
    process(count_inp1_120, SUB_u16_u16_157_157_delayed_1_0_163) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(count_inp1_120, SUB_u16_u16_157_157_delayed_1_0_163, tmp_var);
      my_flag_168 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_83_inst
    process(output_size_buffer) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(output_size_buffer, type_cast_82_wire_constant, tmp_var);
      out_concat_84 <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_205_inst
    process(my_flag_168) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", my_flag_168, tmp_var);
      NOT_u1_u1_205_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_209_inst
    process(NOT_u1_u1_205_wire, ULT_u32_u1_208_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_205_wire, ULT_u32_u1_208_wire, tmp_var);
      continue_flag_210 <= tmp_var; --
    end process;
    -- shared split operator group (9) : SUB_u16_u16_162_inst 
    ApIntSub_group_9: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= total_size_105;
      SUB_u16_u16_157_157_delayed_1_0_163 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u16_u16_162_inst_req_0;
      SUB_u16_u16_162_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u16_u16_162_inst_req_1;
      SUB_u16_u16_162_inst_ack_1 <= ackR_unguarded(0);
      ApIntSub_group_9_gI: SplitGuardInterface generic map(name => "ApIntSub_group_9_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_9",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 9
    -- shared split operator group (10) : SUB_u32_u32_201_inst 
    ApIntSub_group_10: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= out_concat_84;
      SUB_u32_u32_195_195_delayed_1_0_202 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u32_u32_201_inst_req_0;
      SUB_u32_u32_201_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u32_u32_201_inst_req_1;
      SUB_u32_u32_201_inst_ack_1 <= ackR_unguarded(0);
      ApIntSub_group_10_gI: SplitGuardInterface generic map(name => "ApIntSub_group_10_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_10",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 10
    -- binary operator ULT_u16_u1_128_inst
    process(count_inp1_120, input1_count_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(count_inp1_120, input1_count_buffer, tmp_var);
      cmp_129 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_208_inst
    process(add_out_108, SUB_u32_u32_195_195_delayed_1_0_202) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add_out_108, SUB_u32_u32_195_195_delayed_1_0_202, tmp_var);
      ULT_u32_u1_208_wire <= tmp_var; --
    end process;
    -- shared call operator group (0) : call_stmt_135_call call_stmt_141_call 
    readModule1_call_group_0: Block -- 
      signal data_in: std_logic_vector(79 downto 0);
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => true, 1 => true);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 15, 1 => 15);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_135_call_req_0;
      reqL_unguarded(0) <= call_stmt_141_call_req_0;
      call_stmt_135_call_ack_0 <= ackL_unguarded(1);
      call_stmt_141_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_135_call_req_1;
      reqR_unguarded(0) <= call_stmt_141_call_req_1;
      call_stmt_135_call_ack_1 <= ackR_unguarded(1);
      call_stmt_141_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not cmp_129(0);
      guard_vector(1)  <= cmp_129(0);
      readModule1_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "readModule1_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      readModule1_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "readModule1_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      readModule1_call_group_0_gI: SplitGuardInterface generic map(name => "readModule1_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= index1_72 & type_cast_133_wire & index2_75 & type_cast_139_wire;
      i1_135 <= data_out(127 downto 64);
      i2_141 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 80,
        owidth => 40,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 2,
        nreqs => 2,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => readModule1_call_reqs(0),
          ackR => readModule1_call_acks(0),
          dataR => readModule1_call_data(39 downto 0),
          tagR => readModule1_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => readModule1_return_acks(0), -- cross-over
          ackL => readModule1_return_reqs(0), -- cross-over
          dataL => readModule1_return_data(63 downto 0),
          tagL => readModule1_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_158_call 
    writeModule1_call_group_1: Block -- 
      signal data_in: std_logic_vector(103 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 9);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_158_call_req_0;
      call_stmt_158_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_158_call_req_1;
      call_stmt_158_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      writeModule1_call_group_1_gI: SplitGuardInterface generic map(name => "writeModule1_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= index3_78 & add_out_149_delayed_15_0_153 & o_150;
      done_158 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 104,
        owidth => 104,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => writeModule1_call_reqs(0),
          ackR => writeModule1_call_acks(0),
          dataR => writeModule1_call_data(103 downto 0),
          tagR => writeModule1_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 1,
          owidth => 1,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => writeModule1_return_acks(0), -- cross-over
          ackL => writeModule1_return_reqs(0), -- cross-over
          dataL => writeModule1_return_data(0 downto 0),
          tagL => writeModule1_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- 
  end Block; -- data_path
  -- 
end concat_core_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity readModule1 is -- 
  generic (tag_length : integer); 
  port ( -- 
    index : in  std_logic_vector(7 downto 0);
    address : in  std_logic_vector(31 downto 0);
    data : out  std_logic_vector(63 downto 0);
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(15 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity readModule1;
architecture readModule1_arch of readModule1 is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 40)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal index_buffer :  std_logic_vector(7 downto 0);
  signal index_update_enable: Boolean;
  signal address_buffer :  std_logic_vector(31 downto 0);
  signal address_update_enable: Boolean;
  -- output port buffer signals
  signal data_buffer :  std_logic_vector(63 downto 0);
  signal data_update_enable: Boolean;
  signal readModule1_CP_34_start: Boolean;
  signal readModule1_CP_34_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal array_obj_ref_32_index_0_scale_req_0 : boolean;
  signal ptr_deref_37_load_0_req_0 : boolean;
  signal array_obj_ref_32_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_32_index_0_scale_req_1 : boolean;
  signal array_obj_ref_32_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_32_index_sum_1_req_0 : boolean;
  signal array_obj_ref_32_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_32_index_sum_1_req_1 : boolean;
  signal array_obj_ref_32_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_32_index_offset_req_0 : boolean;
  signal array_obj_ref_32_index_offset_ack_0 : boolean;
  signal array_obj_ref_32_index_offset_req_1 : boolean;
  signal array_obj_ref_32_index_offset_ack_1 : boolean;
  signal addr_of_33_final_reg_req_0 : boolean;
  signal addr_of_33_final_reg_ack_0 : boolean;
  signal addr_of_33_final_reg_req_1 : boolean;
  signal addr_of_33_final_reg_ack_1 : boolean;
  signal ptr_deref_37_load_0_ack_0 : boolean;
  signal ptr_deref_37_load_0_req_1 : boolean;
  signal ptr_deref_37_load_0_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "readModule1_input_buffer", -- 
      buffer_size => 2,
      bypass_flag => false,
      data_width => tag_length + 40) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(7 downto 0) <= index;
  index_buffer <= in_buffer_data_out(7 downto 0);
  in_buffer_data_in(39 downto 8) <= address;
  address_buffer <= in_buffer_data_out(39 downto 8);
  in_buffer_data_in(tag_length + 39 downto 40) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 39 downto 40);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 3) := (0 => 8,1 => 8,2 => 1,3 => 8);
    constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 1,3 => 8);
    constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 4); -- 
  begin -- 
    preds <= index_update_enable & address_update_enable & in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  readModule1_CP_34_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "readModule1_out_buffer", -- 
      buffer_size => 2,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= data_buffer;
  data <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 8,1 => 1,2 => 8);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= readModule1_CP_34_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  data_update_enable_join: block -- 
    constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
    constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
    constant place_delays: IntegerArray(0 to 0) := (0 => 0);
    constant joinName: string(1 to 23) := "data_update_enable_join"; 
    signal preds: BooleanArray(1 to 1); -- 
  begin -- 
    preds(1) <= out_buffer_write_ack_symbol;
    gj_data_update_enable_join : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => data_update_enable, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 8,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 8,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= readModule1_CP_34_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 8,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= readModule1_CP_34_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  readModule1_CP_34: Block -- control-path 
    signal readModule1_CP_34_elements: BooleanArray(30 downto 0);
    -- 
  begin -- 
    readModule1_CP_34_elements(0) <= readModule1_CP_34_start;
    readModule1_CP_34_symbol <= readModule1_CP_34_elements(30);
    -- CP-element group 0:  transition  bypass  pipeline-parent 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (1) 
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	9 
    -- CP-element group 1: 	10 
    -- CP-element group 1: 	13 
    -- CP-element group 1: 	14 
    -- CP-element group 1: 	17 
    -- CP-element group 1: 	6 
    -- CP-element group 1:  members (18) 
      -- CP-element group 1: 	 assign_stmt_34_to_assign_stmt_38/$entry
      -- CP-element group 1: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_index_resized_0
      -- CP-element group 1: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_index_computed_0
      -- CP-element group 1: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_index_resize_0/$entry
      -- CP-element group 1: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_index_resize_0/$exit
      -- CP-element group 1: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_index_resize_0/index_resize_req
      -- CP-element group 1: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_index_resize_0/index_resize_ack
      -- CP-element group 1: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_index_resized_2
      -- CP-element group 1: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_index_scaled_2
      -- CP-element group 1: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_index_computed_2
      -- CP-element group 1: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_index_resize_2/$entry
      -- CP-element group 1: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_index_resize_2/$exit
      -- CP-element group 1: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_index_resize_2/index_resize_req
      -- CP-element group 1: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_index_resize_2/index_resize_ack
      -- CP-element group 1: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_index_scale_2/$entry
      -- CP-element group 1: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_index_scale_2/$exit
      -- CP-element group 1: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_index_scale_2/scale_rename_req
      -- CP-element group 1: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_index_scale_2/scale_rename_ack
      -- 
    readModule1_CP_34_elements(1) <= readModule1_CP_34_elements(0);
    -- CP-element group 2:  join  transition  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: marked-predecessors 
    -- CP-element group 2: 	8 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	27 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 assign_stmt_34_to_assign_stmt_38/index_update_enable
      -- CP-element group 2: 	 assign_stmt_34_to_assign_stmt_38/index_update_enable_out
      -- 
    readModule1_cp_element_group_2: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 30) := "readModule1_cp_element_group_2"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= readModule1_CP_34_elements(8);
      gj_readModule1_cp_element_group_2 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readModule1_CP_34_elements(2), clk => clk, reset => reset); --
    end block;
    -- CP-element group 3:  join  transition  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: marked-predecessors 
    -- CP-element group 3: 	15 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	28 
    -- CP-element group 3:  members (2) 
      -- CP-element group 3: 	 assign_stmt_34_to_assign_stmt_38/address_update_enable
      -- CP-element group 3: 	 assign_stmt_34_to_assign_stmt_38/address_update_enable_out
      -- 
    readModule1_cp_element_group_3: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 1);
      constant joinName: string(1 to 30) := "readModule1_cp_element_group_3"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= readModule1_CP_34_elements(15);
      gj_readModule1_cp_element_group_3 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readModule1_CP_34_elements(3), clk => clk, reset => reset); --
    end block;
    -- CP-element group 4:  transition  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	29 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	23 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 assign_stmt_34_to_assign_stmt_38/data_update_enable
      -- CP-element group 4: 	 assign_stmt_34_to_assign_stmt_38/data_update_enable_in
      -- 
    readModule1_CP_34_elements(4) <= readModule1_CP_34_elements(29);
    -- CP-element group 5:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	7 
    -- CP-element group 5: marked-predecessors 
    -- CP-element group 5: 	20 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	20 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 assign_stmt_34_to_assign_stmt_38/addr_of_33_sample_start_
      -- CP-element group 5: 	 assign_stmt_34_to_assign_stmt_38/addr_of_33_request/$entry
      -- CP-element group 5: 	 assign_stmt_34_to_assign_stmt_38/addr_of_33_request/req
      -- 
    req_121_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_121_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readModule1_CP_34_elements(5), ack => addr_of_33_final_reg_req_0); -- 
    readModule1_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "readModule1_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= readModule1_CP_34_elements(7) & readModule1_CP_34_elements(20);
      gj_readModule1_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readModule1_CP_34_elements(5), clk => clk, reset => reset); --
    end block;
    -- CP-element group 6:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	1 
    -- CP-element group 6: marked-predecessors 
    -- CP-element group 6: 	21 
    -- CP-element group 6: 	24 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	21 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 assign_stmt_34_to_assign_stmt_38/addr_of_33_update_start_
      -- CP-element group 6: 	 assign_stmt_34_to_assign_stmt_38/addr_of_33_complete/$entry
      -- CP-element group 6: 	 assign_stmt_34_to_assign_stmt_38/addr_of_33_complete/req
      -- 
    req_126_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_126_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readModule1_CP_34_elements(6), ack => addr_of_33_final_reg_req_1); -- 
    readModule1_cp_element_group_6: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 8,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "readModule1_cp_element_group_6"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= readModule1_CP_34_elements(1) & readModule1_CP_34_elements(21) & readModule1_CP_34_elements(24);
      gj_readModule1_cp_element_group_6 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readModule1_CP_34_elements(6), clk => clk, reset => reset); --
    end block;
    -- CP-element group 7:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	16 
    -- CP-element group 7: 	19 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	5 
    -- CP-element group 7: marked-successors 
    -- CP-element group 7: 	17 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_root_address_calculated
      -- CP-element group 7: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_offset_calculated
      -- CP-element group 7: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_base_plus_offset/$entry
      -- CP-element group 7: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_base_plus_offset/$exit
      -- CP-element group 7: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_base_plus_offset/sum_rename_req
      -- CP-element group 7: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_base_plus_offset/sum_rename_ack
      -- 
    readModule1_cp_element_group_7: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 8,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "readModule1_cp_element_group_7"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= readModule1_CP_34_elements(16) & readModule1_CP_34_elements(19);
      gj_readModule1_cp_element_group_7 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readModule1_CP_34_elements(7), clk => clk, reset => reset); --
    end block;
    -- CP-element group 8:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	12 
    -- CP-element group 8: marked-predecessors 
    -- CP-element group 8: 	15 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	13 
    -- CP-element group 8: marked-successors 
    -- CP-element group 8: 	2 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_index_scaled_0
      -- 
    readModule1_cp_element_group_8: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 8,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "readModule1_cp_element_group_8"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= readModule1_CP_34_elements(12) & readModule1_CP_34_elements(15);
      gj_readModule1_cp_element_group_8 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readModule1_CP_34_elements(8), clk => clk, reset => reset); --
    end block;
    -- CP-element group 9:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	1 
    -- CP-element group 9: marked-predecessors 
    -- CP-element group 9: 	11 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_index_scale_0_Sample/$entry
      -- CP-element group 9: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_index_scale_0_Sample/rr
      -- CP-element group 9: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_index_scale_0_sample_start
      -- 
    rr_67_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_67_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readModule1_CP_34_elements(9), ack => array_obj_ref_32_index_0_scale_req_0); -- 
    readModule1_cp_element_group_9: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 8,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "readModule1_cp_element_group_9"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= readModule1_CP_34_elements(1) & readModule1_CP_34_elements(11);
      gj_readModule1_cp_element_group_9 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readModule1_CP_34_elements(9), clk => clk, reset => reset); --
    end block;
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	1 
    -- CP-element group 10: marked-predecessors 
    -- CP-element group 10: 	12 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	12 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_index_scale_0_update_start
      -- CP-element group 10: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_index_scale_0_Update/$entry
      -- CP-element group 10: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_index_scale_0_Update/cr
      -- 
    cr_72_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_72_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readModule1_CP_34_elements(10), ack => array_obj_ref_32_index_0_scale_req_1); -- 
    readModule1_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 8,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "readModule1_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= readModule1_CP_34_elements(1) & readModule1_CP_34_elements(12);
      gj_readModule1_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readModule1_CP_34_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	26 
    -- CP-element group 11: marked-successors 
    -- CP-element group 11: 	9 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_index_scale_0_Sample/$exit
      -- CP-element group 11: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_index_scale_0_sample_complete
      -- CP-element group 11: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_index_scale_0_Sample/ra
      -- 
    ra_68_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_32_index_0_scale_ack_0, ack => readModule1_CP_34_elements(11)); -- 
    -- CP-element group 12:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	10 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	8 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	10 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_index_scale_0_update_complete
      -- CP-element group 12: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_index_scale_0_Update/$exit
      -- CP-element group 12: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_index_scale_0_Update/ca
      -- 
    ca_73_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_32_index_0_scale_ack_1, ack => readModule1_CP_34_elements(12)); -- 
    -- CP-element group 13:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	1 
    -- CP-element group 13: 	8 
    -- CP-element group 13: marked-predecessors 
    -- CP-element group 13: 	15 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	15 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_partial_sum_1_sample_start
      -- CP-element group 13: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_partial_sum_1_Sample/$entry
      -- CP-element group 13: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_partial_sum_1_Sample/rr
      -- 
    rr_94_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_94_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readModule1_CP_34_elements(13), ack => array_obj_ref_32_index_sum_1_req_0); -- 
    readModule1_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 8,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 31) := "readModule1_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= readModule1_CP_34_elements(1) & readModule1_CP_34_elements(8) & readModule1_CP_34_elements(15);
      gj_readModule1_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readModule1_CP_34_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	1 
    -- CP-element group 14: marked-predecessors 
    -- CP-element group 14: 	16 
    -- CP-element group 14: 	18 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	16 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_partial_sum_1_update_start
      -- CP-element group 14: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_partial_sum_1_Update/$entry
      -- CP-element group 14: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_partial_sum_1_Update/cr
      -- 
    cr_99_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_99_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readModule1_CP_34_elements(14), ack => array_obj_ref_32_index_sum_1_req_1); -- 
    readModule1_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 8,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 31) := "readModule1_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= readModule1_CP_34_elements(1) & readModule1_CP_34_elements(16) & readModule1_CP_34_elements(18);
      gj_readModule1_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readModule1_CP_34_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	13 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	26 
    -- CP-element group 15: marked-successors 
    -- CP-element group 15: 	13 
    -- CP-element group 15: 	3 
    -- CP-element group 15: 	8 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_partial_sum_1_sample_complete
      -- CP-element group 15: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_partial_sum_1_Sample/$exit
      -- CP-element group 15: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_partial_sum_1_Sample/ra
      -- 
    ra_95_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_32_index_sum_1_ack_0, ack => readModule1_CP_34_elements(15)); -- 
    -- CP-element group 16:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	14 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	18 
    -- CP-element group 16: 	7 
    -- CP-element group 16: marked-successors 
    -- CP-element group 16: 	14 
    -- CP-element group 16:  members (5) 
      -- CP-element group 16: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_partial_sum_1_update_complete
      -- CP-element group 16: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_partial_sum_1_Update/$exit
      -- CP-element group 16: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_partial_sum_1_Update/ca
      -- CP-element group 16: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_final_index_sum_regn_Sample/$entry
      -- CP-element group 16: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_final_index_sum_regn_Sample/req
      -- 
    ca_100_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_32_index_sum_1_ack_1, ack => readModule1_CP_34_elements(16)); -- 
    req_106_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_106_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readModule1_CP_34_elements(16), ack => array_obj_ref_32_index_offset_req_0); -- 
    -- CP-element group 17:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	1 
    -- CP-element group 17: marked-predecessors 
    -- CP-element group 17: 	20 
    -- CP-element group 17: 	7 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	19 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_final_index_sum_regn_update_start
      -- CP-element group 17: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_final_index_sum_regn_Update/$entry
      -- CP-element group 17: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_final_index_sum_regn_Update/req
      -- 
    req_111_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_111_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readModule1_CP_34_elements(17), ack => array_obj_ref_32_index_offset_req_1); -- 
    readModule1_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 8,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "readModule1_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= readModule1_CP_34_elements(1) & readModule1_CP_34_elements(20) & readModule1_CP_34_elements(7);
      gj_readModule1_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readModule1_CP_34_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	16 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	26 
    -- CP-element group 18: marked-successors 
    -- CP-element group 18: 	14 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_final_index_sum_regn_sample_complete
      -- CP-element group 18: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_final_index_sum_regn_Sample/$exit
      -- CP-element group 18: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_final_index_sum_regn_Sample/ack
      -- 
    ack_107_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_32_index_offset_ack_0, ack => readModule1_CP_34_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	17 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	7 
    -- CP-element group 19:  members (2) 
      -- CP-element group 19: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_final_index_sum_regn_Update/$exit
      -- CP-element group 19: 	 assign_stmt_34_to_assign_stmt_38/array_obj_ref_32_final_index_sum_regn_Update/ack
      -- 
    ack_112_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_32_index_offset_ack_1, ack => readModule1_CP_34_elements(19)); -- 
    -- CP-element group 20:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	5 
    -- CP-element group 20: successors 
    -- CP-element group 20: marked-successors 
    -- CP-element group 20: 	17 
    -- CP-element group 20: 	5 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 assign_stmt_34_to_assign_stmt_38/addr_of_33_sample_completed_
      -- CP-element group 20: 	 assign_stmt_34_to_assign_stmt_38/addr_of_33_request/$exit
      -- CP-element group 20: 	 assign_stmt_34_to_assign_stmt_38/addr_of_33_request/ack
      -- 
    ack_122_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_33_final_reg_ack_0, ack => readModule1_CP_34_elements(20)); -- 
    -- CP-element group 21:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	6 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21: marked-successors 
    -- CP-element group 21: 	6 
    -- CP-element group 21:  members (19) 
      -- CP-element group 21: 	 assign_stmt_34_to_assign_stmt_38/addr_of_33_update_completed_
      -- CP-element group 21: 	 assign_stmt_34_to_assign_stmt_38/addr_of_33_complete/$exit
      -- CP-element group 21: 	 assign_stmt_34_to_assign_stmt_38/addr_of_33_complete/ack
      -- CP-element group 21: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_base_address_calculated
      -- CP-element group 21: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_word_address_calculated
      -- CP-element group 21: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_root_address_calculated
      -- CP-element group 21: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_base_address_resized
      -- CP-element group 21: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_base_addr_resize/$entry
      -- CP-element group 21: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_base_addr_resize/$exit
      -- CP-element group 21: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_base_addr_resize/base_resize_req
      -- CP-element group 21: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_base_addr_resize/base_resize_ack
      -- CP-element group 21: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_base_plus_offset/$entry
      -- CP-element group 21: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_base_plus_offset/$exit
      -- CP-element group 21: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_base_plus_offset/sum_rename_req
      -- CP-element group 21: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_base_plus_offset/sum_rename_ack
      -- CP-element group 21: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_word_addrgen/$entry
      -- CP-element group 21: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_word_addrgen/$exit
      -- CP-element group 21: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_word_addrgen/root_register_req
      -- CP-element group 21: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_word_addrgen/root_register_ack
      -- 
    ack_127_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_33_final_reg_ack_1, ack => readModule1_CP_34_elements(21)); -- 
    -- CP-element group 22:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: marked-predecessors 
    -- CP-element group 22: 	24 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	24 
    -- CP-element group 22:  members (5) 
      -- CP-element group 22: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_Sample/$entry
      -- CP-element group 22: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_Sample/word_access_start/$entry
      -- CP-element group 22: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_Sample/word_access_start/word_0/$entry
      -- CP-element group 22: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_Sample/word_access_start/word_0/rr
      -- CP-element group 22: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_sample_start_
      -- 
    rr_160_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_160_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readModule1_CP_34_elements(22), ack => ptr_deref_37_load_0_req_0); -- 
    readModule1_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "readModule1_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= readModule1_CP_34_elements(21) & readModule1_CP_34_elements(24);
      gj_readModule1_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readModule1_CP_34_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	4 
    -- CP-element group 23: marked-predecessors 
    -- CP-element group 23: 	25 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	25 
    -- CP-element group 23:  members (5) 
      -- CP-element group 23: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_update_start_
      -- CP-element group 23: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_Update/$entry
      -- CP-element group 23: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_Update/word_access_complete/$entry
      -- CP-element group 23: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_Update/word_access_complete/word_0/$entry
      -- CP-element group 23: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_Update/word_access_complete/word_0/cr
      -- 
    cr_171_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_171_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readModule1_CP_34_elements(23), ack => ptr_deref_37_load_0_req_1); -- 
    readModule1_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 8,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "readModule1_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= readModule1_CP_34_elements(4) & readModule1_CP_34_elements(25);
      gj_readModule1_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readModule1_CP_34_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	22 
    -- CP-element group 24: successors 
    -- CP-element group 24: marked-successors 
    -- CP-element group 24: 	22 
    -- CP-element group 24: 	6 
    -- CP-element group 24:  members (5) 
      -- CP-element group 24: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_Sample/$exit
      -- CP-element group 24: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_Sample/word_access_start/$exit
      -- CP-element group 24: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_Sample/word_access_start/word_0/$exit
      -- CP-element group 24: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_sample_completed_
      -- CP-element group 24: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_Sample/word_access_start/word_0/ra
      -- 
    ra_161_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_37_load_0_ack_0, ack => readModule1_CP_34_elements(24)); -- 
    -- CP-element group 25:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	23 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25: marked-successors 
    -- CP-element group 25: 	23 
    -- CP-element group 25:  members (9) 
      -- CP-element group 25: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_update_completed_
      -- CP-element group 25: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_Update/$exit
      -- CP-element group 25: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_Update/word_access_complete/$exit
      -- CP-element group 25: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_Update/word_access_complete/word_0/$exit
      -- CP-element group 25: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_Update/word_access_complete/word_0/ca
      -- CP-element group 25: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_Update/ptr_deref_37_Merge/$entry
      -- CP-element group 25: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_Update/ptr_deref_37_Merge/$exit
      -- CP-element group 25: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_Update/ptr_deref_37_Merge/merge_req
      -- CP-element group 25: 	 assign_stmt_34_to_assign_stmt_38/ptr_deref_37_Update/ptr_deref_37_Merge/merge_ack
      -- 
    ca_172_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_37_load_0_ack_1, ack => readModule1_CP_34_elements(25)); -- 
    -- CP-element group 26:  join  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	11 
    -- CP-element group 26: 	15 
    -- CP-element group 26: 	18 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	30 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 assign_stmt_34_to_assign_stmt_38/$exit
      -- 
    readModule1_cp_element_group_26: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 8,1 => 8,2 => 8,3 => 8);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 31) := "readModule1_cp_element_group_26"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= readModule1_CP_34_elements(11) & readModule1_CP_34_elements(15) & readModule1_CP_34_elements(18) & readModule1_CP_34_elements(25);
      gj_readModule1_cp_element_group_26 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readModule1_CP_34_elements(26), clk => clk, reset => reset); --
    end block;
    -- CP-element group 27:  place  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	2 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 index_update_enable
      -- 
    readModule1_CP_34_elements(27) <= readModule1_CP_34_elements(2);
    -- CP-element group 28:  place  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	3 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 address_update_enable
      -- 
    readModule1_CP_34_elements(28) <= readModule1_CP_34_elements(3);
    -- CP-element group 29:  place  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	4 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 data_update_enable
      -- 
    -- CP-element group 30:  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	26 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 $exit
      -- 
    readModule1_CP_34_elements(30) <= readModule1_CP_34_elements(26);
    --  hookup: inputs to control-path 
    readModule1_CP_34_elements(29) <= data_update_enable;
    -- hookup: output from control-path 
    index_update_enable <= readModule1_CP_34_elements(27);
    address_update_enable <= readModule1_CP_34_elements(28);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_address_31_resized : std_logic_vector(15 downto 0);
    signal R_address_31_scaled : std_logic_vector(15 downto 0);
    signal array_obj_ref_32_constant_part_of_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_32_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_32_index_partial_sum_1 : std_logic_vector(15 downto 0);
    signal array_obj_ref_32_offset_scale_factor_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_32_offset_scale_factor_1 : std_logic_vector(15 downto 0);
    signal array_obj_ref_32_offset_scale_factor_2 : std_logic_vector(15 downto 0);
    signal array_obj_ref_32_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_32_root_address : std_logic_vector(15 downto 0);
    signal ptr_34 : std_logic_vector(31 downto 0);
    signal ptr_deref_37_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_37_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_37_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_37_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_37_word_offset_0 : std_logic_vector(15 downto 0);
    signal type_cast_28_resized : std_logic_vector(15 downto 0);
    signal type_cast_28_scaled : std_logic_vector(15 downto 0);
    signal type_cast_28_wire : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    array_obj_ref_32_constant_part_of_offset <= "0000000000000000";
    array_obj_ref_32_offset_scale_factor_0 <= "0100000000000000";
    array_obj_ref_32_offset_scale_factor_1 <= "0100000000000000";
    array_obj_ref_32_offset_scale_factor_2 <= "0000000000000001";
    array_obj_ref_32_resized_base_address <= "0000000000000000";
    ptr_deref_37_word_offset_0 <= "0000000000000000";
    addr_of_33_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_33_final_reg_req_0;
      addr_of_33_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_33_final_reg_req_1;
      addr_of_33_final_reg_ack_1<= rack(0);
      addr_of_33_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_33_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_32_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ptr_34,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_28_inst
    process(index_buffer) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := index_buffer(7 downto 0);
      type_cast_28_wire <= tmp_var; -- 
    end process;
    -- equivalence array_obj_ref_32_index_0_resize
    process(type_cast_28_wire) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_28_wire;
      ov := iv(15 downto 0);
      type_cast_28_resized <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_32_index_2_rename
    process(R_address_31_resized) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_address_31_resized;
      ov(15 downto 0) := iv;
      R_address_31_scaled <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_32_index_2_resize
    process(address_buffer) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := address_buffer;
      ov := iv(15 downto 0);
      R_address_31_resized <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_32_root_address_inst
    process(array_obj_ref_32_final_offset) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_32_final_offset;
      ov(15 downto 0) := iv;
      array_obj_ref_32_root_address <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_37_addr_0
    process(ptr_deref_37_root_address) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_37_root_address;
      ov(15 downto 0) := iv;
      ptr_deref_37_word_address_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_37_base_resize
    process(ptr_34) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_34;
      ov := iv(15 downto 0);
      ptr_deref_37_resized_base_address <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_37_gather_scatter
    process(ptr_deref_37_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_37_data_0;
      ov(63 downto 0) := iv;
      data_buffer <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_37_root_address_inst
    process(ptr_deref_37_resized_base_address) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_37_resized_base_address;
      ov(15 downto 0) := iv;
      ptr_deref_37_root_address <= ov(15 downto 0);
      --
    end process;
    -- shared split operator group (0) : array_obj_ref_32_index_0_scale 
    ApIntMul_group_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= type_cast_28_resized;
      type_cast_28_scaled <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_32_index_0_scale_req_0;
      array_obj_ref_32_index_0_scale_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_32_index_0_scale_req_1;
      array_obj_ref_32_index_0_scale_ack_1 <= ackR_unguarded(0);
      ApIntMul_group_0_gI: SplitGuardInterface generic map(name => "ApIntMul_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntMul",
          name => "ApIntMul_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0100000000000000",
          constant_width => 16,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : array_obj_ref_32_index_offset 
    ApIntAdd_group_1: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= array_obj_ref_32_index_partial_sum_1;
      array_obj_ref_32_final_offset <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_32_index_offset_req_0;
      array_obj_ref_32_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_32_index_offset_req_1;
      array_obj_ref_32_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_1_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_1",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : array_obj_ref_32_index_sum_1 
    ApIntAdd_group_2: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_address_31_scaled & type_cast_28_scaled;
      array_obj_ref_32_index_partial_sum_1 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_32_index_sum_1_req_0;
      array_obj_ref_32_index_sum_1_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_32_index_sum_1_req_1;
      array_obj_ref_32_index_sum_1_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_2_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_2",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- shared load operator group (0) : ptr_deref_37_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 6);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_37_load_0_req_0;
      ptr_deref_37_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_37_load_0_req_1;
      ptr_deref_37_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_37_word_address_0;
      ptr_deref_37_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 16,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(15 downto 0),
          mtag => memory_space_0_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- 
  end Block; -- data_path
  -- 
end readModule1_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timer is -- 
  generic (tag_length : integer); 
  port ( -- 
    T : out  std_logic_vector(63 downto 0);
    timer_resp_pipe_read_req : out  std_logic_vector(0 downto 0);
    timer_resp_pipe_read_ack : in   std_logic_vector(0 downto 0);
    timer_resp_pipe_read_data : in   std_logic_vector(63 downto 0);
    timer_req_pipe_write_req : out  std_logic_vector(0 downto 0);
    timer_req_pipe_write_ack : in   std_logic_vector(0 downto 0);
    timer_req_pipe_write_data : out  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timer;
architecture timer_arch of timer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal T_buffer :  std_logic_vector(63 downto 0);
  signal T_update_enable: Boolean;
  signal timer_CP_0_start: Boolean;
  signal timer_CP_0_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal WPIPE_timer_req_13_inst_req_0 : boolean;
  signal WPIPE_timer_req_13_inst_ack_0 : boolean;
  signal WPIPE_timer_req_13_inst_req_1 : boolean;
  signal WPIPE_timer_req_13_inst_ack_1 : boolean;
  signal RPIPE_timer_resp_18_inst_req_0 : boolean;
  signal RPIPE_timer_resp_18_inst_ack_0 : boolean;
  signal RPIPE_timer_resp_18_inst_req_1 : boolean;
  signal RPIPE_timer_resp_18_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timer_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timer_CP_0_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timer_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= T_buffer;
  T <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_0_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timer_CP_0_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_0_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timer_CP_0: Block -- control-path 
    signal timer_CP_0_elements: BooleanArray(5 downto 0);
    -- 
  begin -- 
    timer_CP_0_elements(0) <= timer_CP_0_start;
    timer_CP_0_symbol <= timer_CP_0_elements(5);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	3 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 assign_stmt_16_to_assign_stmt_19/RPIPE_timer_resp_18_sample_start_
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_16_to_assign_stmt_19/$entry
      -- CP-element group 0: 	 assign_stmt_16_to_assign_stmt_19/WPIPE_timer_req_13_sample_start_
      -- CP-element group 0: 	 assign_stmt_16_to_assign_stmt_19/WPIPE_timer_req_13_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_16_to_assign_stmt_19/WPIPE_timer_req_13_Sample/req
      -- CP-element group 0: 	 assign_stmt_16_to_assign_stmt_19/RPIPE_timer_resp_18_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_16_to_assign_stmt_19/RPIPE_timer_resp_18_Sample/rr
      -- 
    req_13_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_13_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_0_elements(0), ack => WPIPE_timer_req_13_inst_req_0); -- 
    rr_27_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_27_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_0_elements(0), ack => RPIPE_timer_resp_18_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 assign_stmt_16_to_assign_stmt_19/WPIPE_timer_req_13_sample_completed_
      -- CP-element group 1: 	 assign_stmt_16_to_assign_stmt_19/WPIPE_timer_req_13_update_start_
      -- CP-element group 1: 	 assign_stmt_16_to_assign_stmt_19/WPIPE_timer_req_13_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_16_to_assign_stmt_19/WPIPE_timer_req_13_Sample/ack
      -- CP-element group 1: 	 assign_stmt_16_to_assign_stmt_19/WPIPE_timer_req_13_Update/$entry
      -- CP-element group 1: 	 assign_stmt_16_to_assign_stmt_19/WPIPE_timer_req_13_Update/req
      -- 
    ack_14_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_req_13_inst_ack_0, ack => timer_CP_0_elements(1)); -- 
    req_18_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_18_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_0_elements(1), ack => WPIPE_timer_req_13_inst_req_1); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (3) 
      -- CP-element group 2: 	 assign_stmt_16_to_assign_stmt_19/WPIPE_timer_req_13_update_completed_
      -- CP-element group 2: 	 assign_stmt_16_to_assign_stmt_19/WPIPE_timer_req_13_Update/$exit
      -- CP-element group 2: 	 assign_stmt_16_to_assign_stmt_19/WPIPE_timer_req_13_Update/ack
      -- 
    ack_19_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_req_13_inst_ack_1, ack => timer_CP_0_elements(2)); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	0 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 assign_stmt_16_to_assign_stmt_19/RPIPE_timer_resp_18_sample_completed_
      -- CP-element group 3: 	 assign_stmt_16_to_assign_stmt_19/RPIPE_timer_resp_18_update_start_
      -- CP-element group 3: 	 assign_stmt_16_to_assign_stmt_19/RPIPE_timer_resp_18_Sample/$exit
      -- CP-element group 3: 	 assign_stmt_16_to_assign_stmt_19/RPIPE_timer_resp_18_Sample/ra
      -- CP-element group 3: 	 assign_stmt_16_to_assign_stmt_19/RPIPE_timer_resp_18_Update/$entry
      -- CP-element group 3: 	 assign_stmt_16_to_assign_stmt_19/RPIPE_timer_resp_18_Update/cr
      -- 
    ra_28_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_resp_18_inst_ack_0, ack => timer_CP_0_elements(3)); -- 
    cr_32_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_32_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_0_elements(3), ack => RPIPE_timer_resp_18_inst_req_1); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 assign_stmt_16_to_assign_stmt_19/RPIPE_timer_resp_18_update_completed_
      -- CP-element group 4: 	 assign_stmt_16_to_assign_stmt_19/RPIPE_timer_resp_18_Update/$exit
      -- CP-element group 4: 	 assign_stmt_16_to_assign_stmt_19/RPIPE_timer_resp_18_Update/ca
      -- 
    ca_33_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_resp_18_inst_ack_1, ack => timer_CP_0_elements(4)); -- 
    -- CP-element group 5:  join  transition  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 $exit
      -- CP-element group 5: 	 assign_stmt_16_to_assign_stmt_19/$exit
      -- 
    timer_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 24) := "timer_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timer_CP_0_elements(4) & timer_CP_0_elements(2);
      gj_timer_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timer_CP_0_elements(5), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal type_cast_15_wire_constant : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    type_cast_15_wire_constant <= "1";
    -- shared inport operator group (0) : RPIPE_timer_resp_18_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(63 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_timer_resp_18_inst_req_0;
      RPIPE_timer_resp_18_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_timer_resp_18_inst_req_1;
      RPIPE_timer_resp_18_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      T_buffer <= data_out(63 downto 0);
      timer_resp_read_0_gI: SplitGuardInterface generic map(name => "timer_resp_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      timer_resp_read_0: InputPortRevised -- 
        generic map ( name => "timer_resp_read_0", data_width => 64,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => timer_resp_pipe_read_req(0),
          oack => timer_resp_pipe_read_ack(0),
          odata => timer_resp_pipe_read_data(63 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_timer_req_13_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_timer_req_13_inst_req_0;
      WPIPE_timer_req_13_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_timer_req_13_inst_req_1;
      WPIPE_timer_req_13_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_15_wire_constant;
      timer_req_write_0_gI: SplitGuardInterface generic map(name => "timer_req_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      timer_req_write_0: OutputPortRevised -- 
        generic map ( name => "timer_req", data_width => 1, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => timer_req_pipe_write_req(0),
          oack => timer_req_pipe_write_ack(0),
          odata => timer_req_pipe_write_data(0 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end timer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timerDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    timer_req_pipe_read_req : out  std_logic_vector(0 downto 0);
    timer_req_pipe_read_ack : in   std_logic_vector(0 downto 0);
    timer_req_pipe_read_data : in   std_logic_vector(0 downto 0);
    timer_resp_pipe_write_req : out  std_logic_vector(0 downto 0);
    timer_resp_pipe_write_ack : in   std_logic_vector(0 downto 0);
    timer_resp_pipe_write_data : out  std_logic_vector(63 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timerDaemon;
architecture timerDaemon_arch of timerDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal timerDaemon_CP_2963_start: Boolean;
  signal timerDaemon_CP_2963_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal WPIPE_timer_resp_1276_inst_ack_1 : boolean;
  signal phi_stmt_1261_req_0 : boolean;
  signal RPIPE_timer_req_1268_inst_ack_0 : boolean;
  signal phi_stmt_1261_ack_0 : boolean;
  signal RPIPE_timer_req_1268_inst_ack_1 : boolean;
  signal do_while_stmt_1259_branch_req_0 : boolean;
  signal WPIPE_timer_resp_1276_inst_req_1 : boolean;
  signal RPIPE_timer_req_1268_inst_req_1 : boolean;
  signal WPIPE_timer_resp_1276_inst_ack_0 : boolean;
  signal do_while_stmt_1259_branch_ack_0 : boolean;
  signal do_while_stmt_1259_branch_ack_1 : boolean;
  signal nCOUNTER_1274_1265_buf_req_0 : boolean;
  signal nCOUNTER_1274_1265_buf_ack_0 : boolean;
  signal nCOUNTER_1274_1265_buf_req_1 : boolean;
  signal nCOUNTER_1274_1265_buf_ack_1 : boolean;
  signal RPIPE_timer_req_1268_inst_req_0 : boolean;
  signal WPIPE_timer_resp_1276_inst_req_0 : boolean;
  signal phi_stmt_1261_req_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timerDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timerDaemon_CP_2963_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timerDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timerDaemon_CP_2963_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timerDaemon_CP_2963_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timerDaemon_CP_2963_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timerDaemon_CP_2963: Block -- control-path 
    signal timerDaemon_CP_2963_elements: BooleanArray(44 downto 0);
    -- 
  begin -- 
    timerDaemon_CP_2963_elements(0) <= timerDaemon_CP_2963_start;
    timerDaemon_CP_2963_symbol <= timerDaemon_CP_2963_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 branch_block_stmt_1258/$entry
      -- CP-element group 0: 	 branch_block_stmt_1258/branch_block_stmt_1258__entry__
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1258/do_while_stmt_1259__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	44 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 branch_block_stmt_1258/do_while_stmt_1259__exit__
      -- CP-element group 1: 	 branch_block_stmt_1258/branch_block_stmt_1258__exit__
      -- CP-element group 1: 	 branch_block_stmt_1258/$exit
      -- CP-element group 1: 	 $exit
      -- 
    timerDaemon_CP_2963_elements(1) <= timerDaemon_CP_2963_elements(44);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259__entry__
      -- CP-element group 2: 	 branch_block_stmt_1258/do_while_stmt_1259/$entry
      -- 
    timerDaemon_CP_2963_elements(2) <= timerDaemon_CP_2963_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	44 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259__exit__
      -- 
    -- Element group timerDaemon_CP_2963_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_1258/do_while_stmt_1259/loop_back
      -- 
    -- Element group timerDaemon_CP_2963_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	42 
    -- CP-element group 5: 	43 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1258/do_while_stmt_1259/condition_done
      -- CP-element group 5: 	 branch_block_stmt_1258/do_while_stmt_1259/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_1258/do_while_stmt_1259/loop_taken/$entry
      -- 
    timerDaemon_CP_2963_elements(5) <= timerDaemon_CP_2963_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	41 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_1258/do_while_stmt_1259/loop_body_done
      -- 
    timerDaemon_CP_2963_elements(6) <= timerDaemon_CP_2963_elements(41);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	19 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/back_edge_to_loop_body
      -- 
    timerDaemon_CP_2963_elements(7) <= timerDaemon_CP_2963_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	21 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/first_time_through_loop_body
      -- 
    timerDaemon_CP_2963_elements(8) <= timerDaemon_CP_2963_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	40 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	32 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	15 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/phi_stmt_1266_sample_start_
      -- 
    -- Element group timerDaemon_CP_2963_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	40 
    -- CP-element group 10: 	14 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/condition_evaluated
      -- 
    condition_evaluated_2987_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_2987_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_2963_elements(10), ack => do_while_stmt_1259_branch_req_0); -- 
    timerDaemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_2963_elements(40) & timerDaemon_CP_2963_elements(14);
      gj_timerDaemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_2963_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: 	15 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	33 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/phi_stmt_1261_sample_start__ps
      -- 
    timerDaemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= timerDaemon_CP_2963_elements(9) & timerDaemon_CP_2963_elements(15) & timerDaemon_CP_2963_elements(14);
      gj_timerDaemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_2963_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	35 
    -- CP-element group 12: 	17 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	41 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	15 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/phi_stmt_1261_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/phi_stmt_1266_sample_completed_
      -- 
    timerDaemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_2963_elements(35) & timerDaemon_CP_2963_elements(17);
      gj_timerDaemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_2963_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	16 
    -- CP-element group 13: 	32 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	34 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/phi_stmt_1261_update_start__ps
      -- 
    timerDaemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_2963_elements(16) & timerDaemon_CP_2963_elements(32);
      gj_timerDaemon_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_2963_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	36 
    -- CP-element group 14: 	18 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/aggregated_phi_update_ack
      -- 
    timerDaemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_2963_elements(36) & timerDaemon_CP_2963_elements(18);
      gj_timerDaemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_2963_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/phi_stmt_1261_sample_start_
      -- 
    timerDaemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_2963_elements(9) & timerDaemon_CP_2963_elements(12);
      gj_timerDaemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_2963_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	38 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/phi_stmt_1261_update_start_
      -- 
    timerDaemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_2963_elements(9) & timerDaemon_CP_2963_elements(38);
      gj_timerDaemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_2963_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	12 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/phi_stmt_1261_sample_completed__ps
      -- 
    -- Element group timerDaemon_CP_2963_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	37 
    -- CP-element group 18: 	14 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/phi_stmt_1261_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/phi_stmt_1261_update_completed__ps
      -- 
    -- Element group timerDaemon_CP_2963_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	7 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/phi_stmt_1261_loopback_trigger
      -- 
    timerDaemon_CP_2963_elements(19) <= timerDaemon_CP_2963_elements(7);
    -- CP-element group 20:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/phi_stmt_1261_loopback_sample_req_ps
      -- CP-element group 20: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/phi_stmt_1261_loopback_sample_req
      -- 
    phi_stmt_1261_loopback_sample_req_3002_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1261_loopback_sample_req_3002_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_2963_elements(20), ack => phi_stmt_1261_req_1); -- 
    -- Element group timerDaemon_CP_2963_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	8 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/phi_stmt_1261_entry_trigger
      -- 
    timerDaemon_CP_2963_elements(21) <= timerDaemon_CP_2963_elements(8);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/phi_stmt_1261_entry_sample_req
      -- CP-element group 22: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/phi_stmt_1261_entry_sample_req_ps
      -- 
    phi_stmt_1261_entry_sample_req_3005_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1261_entry_sample_req_3005_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_2963_elements(22), ack => phi_stmt_1261_req_0); -- 
    -- Element group timerDaemon_CP_2963_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/phi_stmt_1261_phi_mux_ack
      -- CP-element group 23: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/phi_stmt_1261_phi_mux_ack_ps
      -- 
    phi_stmt_1261_phi_mux_ack_3008_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1261_ack_0, ack => timerDaemon_CP_2963_elements(23)); -- 
    -- CP-element group 24:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (4) 
      -- CP-element group 24: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/type_cast_1264_sample_completed__ps
      -- CP-element group 24: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/type_cast_1264_sample_start__ps
      -- CP-element group 24: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/type_cast_1264_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/type_cast_1264_sample_start_
      -- 
    -- Element group timerDaemon_CP_2963_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/type_cast_1264_update_start__ps
      -- CP-element group 25: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/type_cast_1264_update_start_
      -- 
    -- Element group timerDaemon_CP_2963_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/type_cast_1264_update_completed__ps
      -- 
    timerDaemon_CP_2963_elements(26) <= timerDaemon_CP_2963_elements(27);
    -- CP-element group 27:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	26 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/type_cast_1264_update_completed_
      -- 
    -- Element group timerDaemon_CP_2963_elements(27) is a control-delay.
    cp_element_27_delay: control_delay_element  generic map(name => " 27_delay", delay_value => 1)  port map(req => timerDaemon_CP_2963_elements(25), ack => timerDaemon_CP_2963_elements(27), clk => clk, reset =>reset);
    -- CP-element group 28:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/R_nCOUNTER_1265_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/R_nCOUNTER_1265_sample_start__ps
      -- CP-element group 28: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/R_nCOUNTER_1265_Sample/$entry
      -- CP-element group 28: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/R_nCOUNTER_1265_Sample/req
      -- 
    req_3029_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3029_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_2963_elements(28), ack => nCOUNTER_1274_1265_buf_req_0); -- 
    -- Element group timerDaemon_CP_2963_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/R_nCOUNTER_1265_update_start__ps
      -- CP-element group 29: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/R_nCOUNTER_1265_update_start_
      -- CP-element group 29: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/R_nCOUNTER_1265_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/R_nCOUNTER_1265_Update/req
      -- 
    req_3034_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3034_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_2963_elements(29), ack => nCOUNTER_1274_1265_buf_req_1); -- 
    -- Element group timerDaemon_CP_2963_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/R_nCOUNTER_1265_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/R_nCOUNTER_1265_sample_completed__ps
      -- CP-element group 30: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/R_nCOUNTER_1265_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/R_nCOUNTER_1265_Sample/ack
      -- 
    ack_3030_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nCOUNTER_1274_1265_buf_ack_0, ack => timerDaemon_CP_2963_elements(30)); -- 
    -- CP-element group 31:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/R_nCOUNTER_1265_update_completed__ps
      -- CP-element group 31: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/R_nCOUNTER_1265_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/R_nCOUNTER_1265_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/R_nCOUNTER_1265_Update/ack
      -- 
    ack_3035_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nCOUNTER_1274_1265_buf_ack_1, ack => timerDaemon_CP_2963_elements(31)); -- 
    -- CP-element group 32:  join  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	9 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	38 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	13 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/phi_stmt_1266_update_start_
      -- 
    timerDaemon_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_2963_elements(9) & timerDaemon_CP_2963_elements(38);
      gj_timerDaemon_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_2963_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	11 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	36 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/RPIPE_timer_req_1268_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/RPIPE_timer_req_1268_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/RPIPE_timer_req_1268_Sample/rr
      -- 
    rr_3048_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3048_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_2963_elements(33), ack => RPIPE_timer_req_1268_inst_req_0); -- 
    timerDaemon_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_2963_elements(11) & timerDaemon_CP_2963_elements(36);
      gj_timerDaemon_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_2963_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	13 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/RPIPE_timer_req_1268_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/RPIPE_timer_req_1268_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/RPIPE_timer_req_1268_Update/cr
      -- 
    cr_3053_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3053_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_2963_elements(34), ack => RPIPE_timer_req_1268_inst_req_1); -- 
    timerDaemon_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_2963_elements(35) & timerDaemon_CP_2963_elements(13);
      gj_timerDaemon_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_2963_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: 	12 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/RPIPE_timer_req_1268_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/RPIPE_timer_req_1268_Sample/ra
      -- CP-element group 35: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/RPIPE_timer_req_1268_Sample/$exit
      -- 
    ra_3049_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_req_1268_inst_ack_0, ack => timerDaemon_CP_2963_elements(35)); -- 
    -- CP-element group 36:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	37 
    -- CP-element group 36: 	14 
    -- CP-element group 36: marked-successors 
    -- CP-element group 36: 	33 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/RPIPE_timer_req_1268_Update/ca
      -- CP-element group 36: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/RPIPE_timer_req_1268_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/RPIPE_timer_req_1268_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/phi_stmt_1266_update_completed_
      -- 
    ca_3054_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_req_1268_inst_ack_1, ack => timerDaemon_CP_2963_elements(36)); -- 
    -- CP-element group 37:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	36 
    -- CP-element group 37: 	18 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	39 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/WPIPE_timer_resp_1276_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/WPIPE_timer_resp_1276_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/WPIPE_timer_resp_1276_Sample/req
      -- 
    req_3062_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3062_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_2963_elements(37), ack => WPIPE_timer_resp_1276_inst_req_0); -- 
    timerDaemon_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 7,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= timerDaemon_CP_2963_elements(36) & timerDaemon_CP_2963_elements(18) & timerDaemon_CP_2963_elements(39);
      gj_timerDaemon_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_2963_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38: marked-successors 
    -- CP-element group 38: 	16 
    -- CP-element group 38: 	32 
    -- CP-element group 38:  members (6) 
      -- CP-element group 38: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/WPIPE_timer_resp_1276_Update/$entry
      -- CP-element group 38: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/WPIPE_timer_resp_1276_Update/req
      -- CP-element group 38: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/WPIPE_timer_resp_1276_Sample/ack
      -- CP-element group 38: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/WPIPE_timer_resp_1276_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/WPIPE_timer_resp_1276_update_start_
      -- CP-element group 38: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/WPIPE_timer_resp_1276_Sample/$exit
      -- 
    ack_3063_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_resp_1276_inst_ack_0, ack => timerDaemon_CP_2963_elements(38)); -- 
    req_3067_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3067_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_2963_elements(38), ack => WPIPE_timer_resp_1276_inst_req_1); -- 
    -- CP-element group 39:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	41 
    -- CP-element group 39: marked-successors 
    -- CP-element group 39: 	37 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/WPIPE_timer_resp_1276_Update/ack
      -- CP-element group 39: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/WPIPE_timer_resp_1276_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/WPIPE_timer_resp_1276_update_completed_
      -- 
    ack_3068_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_resp_1276_inst_ack_1, ack => timerDaemon_CP_2963_elements(39)); -- 
    -- CP-element group 40:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	9 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	10 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group timerDaemon_CP_2963_elements(40) is a control-delay.
    cp_element_40_delay: control_delay_element  generic map(name => " 40_delay", delay_value => 1)  port map(req => timerDaemon_CP_2963_elements(9), ack => timerDaemon_CP_2963_elements(40), clk => clk, reset =>reset);
    -- CP-element group 41:  join  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	39 
    -- CP-element group 41: 	12 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	6 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_1258/do_while_stmt_1259/do_while_stmt_1259_loop_body/$exit
      -- 
    timerDaemon_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_2963_elements(39) & timerDaemon_CP_2963_elements(12);
      gj_timerDaemon_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_2963_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  transition  input  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	5 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (2) 
      -- CP-element group 42: 	 branch_block_stmt_1258/do_while_stmt_1259/loop_exit/ack
      -- CP-element group 42: 	 branch_block_stmt_1258/do_while_stmt_1259/loop_exit/$exit
      -- 
    ack_3073_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1259_branch_ack_0, ack => timerDaemon_CP_2963_elements(42)); -- 
    -- CP-element group 43:  transition  input  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	5 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (2) 
      -- CP-element group 43: 	 branch_block_stmt_1258/do_while_stmt_1259/loop_taken/$exit
      -- CP-element group 43: 	 branch_block_stmt_1258/do_while_stmt_1259/loop_taken/ack
      -- 
    ack_3077_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1259_branch_ack_1, ack => timerDaemon_CP_2963_elements(43)); -- 
    -- CP-element group 44:  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	3 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	1 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 branch_block_stmt_1258/do_while_stmt_1259/$exit
      -- 
    timerDaemon_CP_2963_elements(44) <= timerDaemon_CP_2963_elements(3);
    timerDaemon_do_while_stmt_1259_terminator_3078: loop_terminator -- 
      generic map (name => " timerDaemon_do_while_stmt_1259_terminator_3078", max_iterations_in_flight =>7) 
      port map(loop_body_exit => timerDaemon_CP_2963_elements(6),loop_continue => timerDaemon_CP_2963_elements(43),loop_terminate => timerDaemon_CP_2963_elements(42),loop_back => timerDaemon_CP_2963_elements(4),loop_exit => timerDaemon_CP_2963_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_1261_phi_seq_3036_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= timerDaemon_CP_2963_elements(21);
      timerDaemon_CP_2963_elements(24)<= src_sample_reqs(0);
      src_sample_acks(0)  <= timerDaemon_CP_2963_elements(24);
      timerDaemon_CP_2963_elements(25)<= src_update_reqs(0);
      src_update_acks(0)  <= timerDaemon_CP_2963_elements(26);
      timerDaemon_CP_2963_elements(22) <= phi_mux_reqs(0);
      triggers(1)  <= timerDaemon_CP_2963_elements(19);
      timerDaemon_CP_2963_elements(28)<= src_sample_reqs(1);
      src_sample_acks(1)  <= timerDaemon_CP_2963_elements(30);
      timerDaemon_CP_2963_elements(29)<= src_update_reqs(1);
      src_update_acks(1)  <= timerDaemon_CP_2963_elements(31);
      timerDaemon_CP_2963_elements(20) <= phi_mux_reqs(1);
      phi_stmt_1261_phi_seq_3036 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1261_phi_seq_3036") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => timerDaemon_CP_2963_elements(11), 
          phi_sample_ack => timerDaemon_CP_2963_elements(17), 
          phi_update_req => timerDaemon_CP_2963_elements(13), 
          phi_update_ack => timerDaemon_CP_2963_elements(18), 
          phi_mux_ack => timerDaemon_CP_2963_elements(23), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_2988_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= timerDaemon_CP_2963_elements(7);
        preds(1)  <= timerDaemon_CP_2963_elements(8);
        entry_tmerge_2988 : transition_merge -- 
          generic map(name => " entry_tmerge_2988")
          port map (preds => preds, symbol_out => timerDaemon_CP_2963_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal COUNTER_1261 : std_logic_vector(63 downto 0);
    signal RPIPE_timer_req_1268_wire : std_logic_vector(0 downto 0);
    signal konst_1272_wire_constant : std_logic_vector(63 downto 0);
    signal konst_1280_wire_constant : std_logic_vector(0 downto 0);
    signal nCOUNTER_1274 : std_logic_vector(63 downto 0);
    signal nCOUNTER_1274_1265_buffered : std_logic_vector(63 downto 0);
    signal req_1266 : std_logic_vector(0 downto 0);
    signal type_cast_1264_wire_constant : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    konst_1272_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    konst_1280_wire_constant <= "1";
    type_cast_1264_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    phi_stmt_1261: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1264_wire_constant & nCOUNTER_1274_1265_buffered;
      req <= phi_stmt_1261_req_0 & phi_stmt_1261_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1261",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1261_ack_0,
          idata => idata,
          odata => COUNTER_1261,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1261
    nCOUNTER_1274_1265_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nCOUNTER_1274_1265_buf_req_0;
      nCOUNTER_1274_1265_buf_ack_0<= wack(0);
      rreq(0) <= nCOUNTER_1274_1265_buf_req_1;
      nCOUNTER_1274_1265_buf_ack_1<= rack(0);
      nCOUNTER_1274_1265_buf : InterlockBuffer generic map ( -- 
        name => "nCOUNTER_1274_1265_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nCOUNTER_1274,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nCOUNTER_1274_1265_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock ssrc_phi_stmt_1266
    process(RPIPE_timer_req_1268_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := RPIPE_timer_req_1268_wire(0 downto 0);
      req_1266 <= tmp_var; -- 
    end process;
    do_while_stmt_1259_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_1280_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1259_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1259_branch_req_0,
          ack0 => do_while_stmt_1259_branch_ack_0,
          ack1 => do_while_stmt_1259_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u64_u64_1273_inst
    process(COUNTER_1261) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(COUNTER_1261, konst_1272_wire_constant, tmp_var);
      nCOUNTER_1274 <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_timer_req_1268_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(0 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_timer_req_1268_inst_req_0;
      RPIPE_timer_req_1268_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_timer_req_1268_inst_req_1;
      RPIPE_timer_req_1268_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_timer_req_1268_wire <= data_out(0 downto 0);
      timer_req_read_0_gI: SplitGuardInterface generic map(name => "timer_req_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      timer_req_read_0: InputPortRevised -- 
        generic map ( name => "timer_req_read_0", data_width => 1,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => timer_req_pipe_read_req(0),
          oack => timer_req_pipe_read_ack(0),
          odata => timer_req_pipe_read_data(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_timer_resp_1276_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_timer_resp_1276_inst_req_0;
      WPIPE_timer_resp_1276_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_timer_resp_1276_inst_req_1;
      WPIPE_timer_resp_1276_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= req_1266(0);
      data_in <= COUNTER_1261;
      timer_resp_write_0_gI: SplitGuardInterface generic map(name => "timer_resp_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      timer_resp_write_0: OutputPortRevised -- 
        generic map ( name => "timer_resp", data_width => 64, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => timer_resp_pipe_write_req(0),
          oack => timer_resp_pipe_write_ack(0),
          odata => timer_resp_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end timerDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity writeModule1 is -- 
  generic (tag_length : integer); 
  port ( -- 
    index : in  std_logic_vector(7 downto 0);
    address : in  std_logic_vector(31 downto 0);
    data : in  std_logic_vector(63 downto 0);
    done : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(15 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity writeModule1;
architecture writeModule1_arch of writeModule1 is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 104)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 1)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal index_buffer :  std_logic_vector(7 downto 0);
  signal index_update_enable: Boolean;
  signal address_buffer :  std_logic_vector(31 downto 0);
  signal address_update_enable: Boolean;
  signal data_buffer :  std_logic_vector(63 downto 0);
  signal data_update_enable: Boolean;
  -- output port buffer signals
  signal done_buffer :  std_logic_vector(0 downto 0);
  signal done_update_enable: Boolean;
  signal writeModule1_CP_181_start: Boolean;
  signal writeModule1_CP_181_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal array_obj_ref_51_index_0_scale_req_0 : boolean;
  signal array_obj_ref_51_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_51_index_0_scale_req_1 : boolean;
  signal array_obj_ref_51_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_51_index_sum_1_req_0 : boolean;
  signal array_obj_ref_51_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_51_index_sum_1_req_1 : boolean;
  signal array_obj_ref_51_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_51_index_offset_req_0 : boolean;
  signal array_obj_ref_51_index_offset_ack_0 : boolean;
  signal array_obj_ref_51_index_offset_req_1 : boolean;
  signal array_obj_ref_51_index_offset_ack_1 : boolean;
  signal addr_of_52_final_reg_req_0 : boolean;
  signal addr_of_52_final_reg_ack_0 : boolean;
  signal addr_of_52_final_reg_req_1 : boolean;
  signal addr_of_52_final_reg_ack_1 : boolean;
  signal ptr_deref_55_store_0_req_0 : boolean;
  signal ptr_deref_55_store_0_ack_0 : boolean;
  signal ptr_deref_55_store_0_req_1 : boolean;
  signal ptr_deref_55_store_0_ack_1 : boolean;
  signal BITSEL_u8_u1_61_inst_req_0 : boolean;
  signal BITSEL_u8_u1_61_inst_ack_0 : boolean;
  signal BITSEL_u8_u1_61_inst_req_1 : boolean;
  signal BITSEL_u8_u1_61_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "writeModule1_input_buffer", -- 
      buffer_size => 2,
      bypass_flag => false,
      data_width => tag_length + 104) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(7 downto 0) <= index;
  index_buffer <= in_buffer_data_out(7 downto 0);
  in_buffer_data_in(39 downto 8) <= address;
  address_buffer <= in_buffer_data_out(39 downto 8);
  in_buffer_data_in(103 downto 40) <= data;
  data_buffer <= in_buffer_data_out(103 downto 40);
  in_buffer_data_in(tag_length + 103 downto 104) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 103 downto 104);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 4) := (0 => 8,1 => 8,2 => 8,3 => 1,4 => 8);
    constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 8);
    constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 5); -- 
  begin -- 
    preds <= index_update_enable & address_update_enable & data_update_enable & in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  writeModule1_CP_181_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "writeModule1_out_buffer", -- 
      buffer_size => 2,
      full_rate => false,
      data_width => tag_length + 1) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(0 downto 0) <= done_buffer;
  done <= out_buffer_data_out(0 downto 0);
  out_buffer_data_in(tag_length + 0 downto 1) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 0 downto 1);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 8,1 => 1,2 => 8);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= writeModule1_CP_181_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  done_update_enable_join: block -- 
    constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
    constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
    constant place_delays: IntegerArray(0 to 0) := (0 => 0);
    constant joinName: string(1 to 23) := "done_update_enable_join"; 
    signal preds: BooleanArray(1 to 1); -- 
  begin -- 
    preds(1) <= out_buffer_write_ack_symbol;
    gj_done_update_enable_join : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => done_update_enable, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 8,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 8,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= writeModule1_CP_181_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 8,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= writeModule1_CP_181_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  writeModule1_CP_181: Block -- control-path 
    signal writeModule1_CP_181_elements: BooleanArray(36 downto 0);
    -- 
  begin -- 
    writeModule1_CP_181_elements(0) <= writeModule1_CP_181_start;
    writeModule1_CP_181_symbol <= writeModule1_CP_181_elements(36);
    -- CP-element group 0:  transition  bypass  pipeline-parent 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (1) 
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	18 
    -- CP-element group 1: 	27 
    -- CP-element group 1: 	15 
    -- CP-element group 1: 	14 
    -- CP-element group 1: 	10 
    -- CP-element group 1: 	7 
    -- CP-element group 1: 	23 
    -- CP-element group 1: 	11 
    -- CP-element group 1:  members (18) 
      -- CP-element group 1: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_index_resized_0
      -- CP-element group 1: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_index_computed_0
      -- CP-element group 1: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_index_resize_0/$entry
      -- CP-element group 1: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_index_resize_0/$exit
      -- CP-element group 1: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_index_resize_0/index_resize_req
      -- CP-element group 1: 	 assign_stmt_53_to_assign_stmt_62/$entry
      -- CP-element group 1: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_index_resize_0/index_resize_ack
      -- CP-element group 1: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_index_resized_2
      -- CP-element group 1: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_index_scaled_2
      -- CP-element group 1: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_index_computed_2
      -- CP-element group 1: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_index_resize_2/$entry
      -- CP-element group 1: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_index_resize_2/$exit
      -- CP-element group 1: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_index_resize_2/index_resize_req
      -- CP-element group 1: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_index_resize_2/index_resize_ack
      -- CP-element group 1: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_index_scale_2/$entry
      -- CP-element group 1: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_index_scale_2/$exit
      -- CP-element group 1: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_index_scale_2/scale_rename_req
      -- CP-element group 1: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_index_scale_2/scale_rename_ack
      -- 
    writeModule1_CP_181_elements(1) <= writeModule1_CP_181_elements(0);
    -- CP-element group 2:  join  transition  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: marked-predecessors 
    -- CP-element group 2: 	29 
    -- CP-element group 2: 	9 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	32 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 assign_stmt_53_to_assign_stmt_62/index_update_enable
      -- CP-element group 2: 	 assign_stmt_53_to_assign_stmt_62/index_update_enable_out
      -- 
    writeModule1_cp_element_group_2: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "writeModule1_cp_element_group_2"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeModule1_CP_181_elements(29) & writeModule1_CP_181_elements(9);
      gj_writeModule1_cp_element_group_2 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeModule1_CP_181_elements(2), clk => clk, reset => reset); --
    end block;
    -- CP-element group 3:  join  transition  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: marked-predecessors 
    -- CP-element group 3: 	16 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	33 
    -- CP-element group 3:  members (2) 
      -- CP-element group 3: 	 assign_stmt_53_to_assign_stmt_62/address_update_enable
      -- CP-element group 3: 	 assign_stmt_53_to_assign_stmt_62/address_update_enable_out
      -- 
    writeModule1_cp_element_group_3: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 1);
      constant joinName: string(1 to 31) := "writeModule1_cp_element_group_3"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= writeModule1_CP_181_elements(16);
      gj_writeModule1_cp_element_group_3 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeModule1_CP_181_elements(3), clk => clk, reset => reset); --
    end block;
    -- CP-element group 4:  join  transition  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: marked-predecessors 
    -- CP-element group 4: 	25 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	34 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 assign_stmt_53_to_assign_stmt_62/data_update_enable
      -- CP-element group 4: 	 assign_stmt_53_to_assign_stmt_62/data_update_enable_out
      -- 
    writeModule1_cp_element_group_4: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "writeModule1_cp_element_group_4"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= writeModule1_CP_181_elements(25);
      gj_writeModule1_cp_element_group_4 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeModule1_CP_181_elements(4), clk => clk, reset => reset); --
    end block;
    -- CP-element group 5:  transition  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	35 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	28 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 assign_stmt_53_to_assign_stmt_62/done_update_enable
      -- CP-element group 5: 	 assign_stmt_53_to_assign_stmt_62/done_update_enable_in
      -- 
    writeModule1_CP_181_elements(5) <= writeModule1_CP_181_elements(35);
    -- CP-element group 6:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	8 
    -- CP-element group 6: marked-predecessors 
    -- CP-element group 6: 	21 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	21 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 assign_stmt_53_to_assign_stmt_62/addr_of_52_sample_start_
      -- CP-element group 6: 	 assign_stmt_53_to_assign_stmt_62/addr_of_52_request/$entry
      -- CP-element group 6: 	 assign_stmt_53_to_assign_stmt_62/addr_of_52_request/req
      -- 
    req_270_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_270_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeModule1_CP_181_elements(6), ack => addr_of_52_final_reg_req_0); -- 
    writeModule1_cp_element_group_6: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "writeModule1_cp_element_group_6"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeModule1_CP_181_elements(8) & writeModule1_CP_181_elements(21);
      gj_writeModule1_cp_element_group_6 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeModule1_CP_181_elements(6), clk => clk, reset => reset); --
    end block;
    -- CP-element group 7:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	1 
    -- CP-element group 7: marked-predecessors 
    -- CP-element group 7: 	25 
    -- CP-element group 7: 	22 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	22 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 assign_stmt_53_to_assign_stmt_62/addr_of_52_update_start_
      -- CP-element group 7: 	 assign_stmt_53_to_assign_stmt_62/addr_of_52_complete/$entry
      -- CP-element group 7: 	 assign_stmt_53_to_assign_stmt_62/addr_of_52_complete/req
      -- 
    req_275_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_275_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeModule1_CP_181_elements(7), ack => addr_of_52_final_reg_req_1); -- 
    writeModule1_cp_element_group_7: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 8,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "writeModule1_cp_element_group_7"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= writeModule1_CP_181_elements(1) & writeModule1_CP_181_elements(25) & writeModule1_CP_181_elements(22);
      gj_writeModule1_cp_element_group_7 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeModule1_CP_181_elements(7), clk => clk, reset => reset); --
    end block;
    -- CP-element group 8:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	20 
    -- CP-element group 8: 	17 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	6 
    -- CP-element group 8: marked-successors 
    -- CP-element group 8: 	18 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_root_address_calculated
      -- CP-element group 8: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_offset_calculated
      -- CP-element group 8: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_base_plus_offset/$entry
      -- CP-element group 8: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_base_plus_offset/$exit
      -- CP-element group 8: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_base_plus_offset/sum_rename_req
      -- CP-element group 8: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_base_plus_offset/sum_rename_ack
      -- 
    writeModule1_cp_element_group_8: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 8);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "writeModule1_cp_element_group_8"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeModule1_CP_181_elements(20) & writeModule1_CP_181_elements(17);
      gj_writeModule1_cp_element_group_8 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeModule1_CP_181_elements(8), clk => clk, reset => reset); --
    end block;
    -- CP-element group 9:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	13 
    -- CP-element group 9: marked-predecessors 
    -- CP-element group 9: 	16 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	14 
    -- CP-element group 9: marked-successors 
    -- CP-element group 9: 	2 
    -- CP-element group 9:  members (1) 
      -- CP-element group 9: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_index_scaled_0
      -- 
    writeModule1_cp_element_group_9: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 8,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "writeModule1_cp_element_group_9"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeModule1_CP_181_elements(13) & writeModule1_CP_181_elements(16);
      gj_writeModule1_cp_element_group_9 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeModule1_CP_181_elements(9), clk => clk, reset => reset); --
    end block;
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	1 
    -- CP-element group 10: marked-predecessors 
    -- CP-element group 10: 	12 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	12 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_index_scale_0_sample_start
      -- CP-element group 10: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_index_scale_0_Sample/$entry
      -- CP-element group 10: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_index_scale_0_Sample/rr
      -- 
    rr_216_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_216_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeModule1_CP_181_elements(10), ack => array_obj_ref_51_index_0_scale_req_0); -- 
    writeModule1_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 8,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 32) := "writeModule1_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeModule1_CP_181_elements(1) & writeModule1_CP_181_elements(12);
      gj_writeModule1_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeModule1_CP_181_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	1 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	13 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	13 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_index_scale_0_update_start
      -- CP-element group 11: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_index_scale_0_Update/$entry
      -- CP-element group 11: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_index_scale_0_Update/cr
      -- 
    cr_221_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_221_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeModule1_CP_181_elements(11), ack => array_obj_ref_51_index_0_scale_req_1); -- 
    writeModule1_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 8,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "writeModule1_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeModule1_CP_181_elements(1) & writeModule1_CP_181_elements(13);
      gj_writeModule1_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeModule1_CP_181_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	10 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	31 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	10 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_index_scale_0_sample_complete
      -- CP-element group 12: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_index_scale_0_Sample/$exit
      -- CP-element group 12: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_index_scale_0_Sample/ra
      -- 
    ra_217_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_51_index_0_scale_ack_0, ack => writeModule1_CP_181_elements(12)); -- 
    -- CP-element group 13:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	11 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	9 
    -- CP-element group 13: marked-successors 
    -- CP-element group 13: 	11 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_index_scale_0_update_complete
      -- CP-element group 13: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_index_scale_0_Update/$exit
      -- CP-element group 13: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_index_scale_0_Update/ca
      -- 
    ca_222_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_51_index_0_scale_ack_1, ack => writeModule1_CP_181_elements(13)); -- 
    -- CP-element group 14:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	9 
    -- CP-element group 14: 	1 
    -- CP-element group 14: marked-predecessors 
    -- CP-element group 14: 	16 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	16 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_partial_sum_1_sample_start
      -- CP-element group 14: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_partial_sum_1_Sample/$entry
      -- CP-element group 14: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_partial_sum_1_Sample/rr
      -- 
    rr_243_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_243_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeModule1_CP_181_elements(14), ack => array_obj_ref_51_index_sum_1_req_0); -- 
    writeModule1_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 8,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 32) := "writeModule1_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= writeModule1_CP_181_elements(9) & writeModule1_CP_181_elements(1) & writeModule1_CP_181_elements(16);
      gj_writeModule1_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeModule1_CP_181_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	1 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	17 
    -- CP-element group 15: 	19 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	17 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_partial_sum_1_update_start
      -- CP-element group 15: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_partial_sum_1_Update/$entry
      -- CP-element group 15: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_partial_sum_1_Update/cr
      -- 
    cr_248_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_248_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeModule1_CP_181_elements(15), ack => array_obj_ref_51_index_sum_1_req_1); -- 
    writeModule1_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 8,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 32) := "writeModule1_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= writeModule1_CP_181_elements(1) & writeModule1_CP_181_elements(17) & writeModule1_CP_181_elements(19);
      gj_writeModule1_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeModule1_CP_181_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	14 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	31 
    -- CP-element group 16: marked-successors 
    -- CP-element group 16: 	14 
    -- CP-element group 16: 	3 
    -- CP-element group 16: 	9 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_partial_sum_1_sample_complete
      -- CP-element group 16: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_partial_sum_1_Sample/$exit
      -- CP-element group 16: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_partial_sum_1_Sample/ra
      -- 
    ra_244_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_51_index_sum_1_ack_0, ack => writeModule1_CP_181_elements(16)); -- 
    -- CP-element group 17:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	15 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	8 
    -- CP-element group 17: 	19 
    -- CP-element group 17: marked-successors 
    -- CP-element group 17: 	15 
    -- CP-element group 17:  members (5) 
      -- CP-element group 17: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_partial_sum_1_update_complete
      -- CP-element group 17: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_partial_sum_1_Update/$exit
      -- CP-element group 17: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_partial_sum_1_Update/ca
      -- CP-element group 17: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_final_index_sum_regn_Sample/$entry
      -- CP-element group 17: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_final_index_sum_regn_Sample/req
      -- 
    ca_249_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_51_index_sum_1_ack_1, ack => writeModule1_CP_181_elements(17)); -- 
    req_255_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_255_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeModule1_CP_181_elements(17), ack => array_obj_ref_51_index_offset_req_0); -- 
    -- CP-element group 18:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	1 
    -- CP-element group 18: marked-predecessors 
    -- CP-element group 18: 	21 
    -- CP-element group 18: 	8 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	20 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_final_index_sum_regn_update_start
      -- CP-element group 18: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_final_index_sum_regn_Update/$entry
      -- CP-element group 18: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_final_index_sum_regn_Update/req
      -- 
    req_260_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_260_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeModule1_CP_181_elements(18), ack => array_obj_ref_51_index_offset_req_1); -- 
    writeModule1_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 8,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "writeModule1_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= writeModule1_CP_181_elements(1) & writeModule1_CP_181_elements(21) & writeModule1_CP_181_elements(8);
      gj_writeModule1_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeModule1_CP_181_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	17 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	31 
    -- CP-element group 19: marked-successors 
    -- CP-element group 19: 	15 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_final_index_sum_regn_sample_complete
      -- CP-element group 19: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_final_index_sum_regn_Sample/$exit
      -- CP-element group 19: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_final_index_sum_regn_Sample/ack
      -- 
    ack_256_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_51_index_offset_ack_0, ack => writeModule1_CP_181_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	18 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	8 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_final_index_sum_regn_Update/$exit
      -- CP-element group 20: 	 assign_stmt_53_to_assign_stmt_62/array_obj_ref_51_final_index_sum_regn_Update/ack
      -- 
    ack_261_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_51_index_offset_ack_1, ack => writeModule1_CP_181_elements(20)); -- 
    -- CP-element group 21:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	6 
    -- CP-element group 21: successors 
    -- CP-element group 21: marked-successors 
    -- CP-element group 21: 	18 
    -- CP-element group 21: 	6 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 assign_stmt_53_to_assign_stmt_62/addr_of_52_sample_completed_
      -- CP-element group 21: 	 assign_stmt_53_to_assign_stmt_62/addr_of_52_request/$exit
      -- CP-element group 21: 	 assign_stmt_53_to_assign_stmt_62/addr_of_52_request/ack
      -- 
    ack_271_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_52_final_reg_ack_0, ack => writeModule1_CP_181_elements(21)); -- 
    -- CP-element group 22:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	7 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22: marked-successors 
    -- CP-element group 22: 	7 
    -- CP-element group 22:  members (19) 
      -- CP-element group 22: 	 assign_stmt_53_to_assign_stmt_62/addr_of_52_update_completed_
      -- CP-element group 22: 	 assign_stmt_53_to_assign_stmt_62/addr_of_52_complete/$exit
      -- CP-element group 22: 	 assign_stmt_53_to_assign_stmt_62/addr_of_52_complete/ack
      -- CP-element group 22: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_base_address_calculated
      -- CP-element group 22: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_word_address_calculated
      -- CP-element group 22: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_root_address_calculated
      -- CP-element group 22: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_base_address_resized
      -- CP-element group 22: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_base_addr_resize/$entry
      -- CP-element group 22: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_base_addr_resize/$exit
      -- CP-element group 22: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_base_addr_resize/base_resize_req
      -- CP-element group 22: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_base_addr_resize/base_resize_ack
      -- CP-element group 22: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_base_plus_offset/$entry
      -- CP-element group 22: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_base_plus_offset/$exit
      -- CP-element group 22: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_base_plus_offset/sum_rename_req
      -- CP-element group 22: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_base_plus_offset/sum_rename_ack
      -- CP-element group 22: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_word_addrgen/$entry
      -- CP-element group 22: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_word_addrgen/$exit
      -- CP-element group 22: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_word_addrgen/root_register_req
      -- CP-element group 22: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_word_addrgen/root_register_ack
      -- 
    ack_276_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_52_final_reg_ack_1, ack => writeModule1_CP_181_elements(22)); -- 
    -- CP-element group 23:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	1 
    -- CP-element group 23: 	22 
    -- CP-element group 23: marked-predecessors 
    -- CP-element group 23: 	25 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	25 
    -- CP-element group 23:  members (9) 
      -- CP-element group 23: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_sample_start_
      -- CP-element group 23: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_Sample/$entry
      -- CP-element group 23: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_Sample/ptr_deref_55_Split/$entry
      -- CP-element group 23: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_Sample/ptr_deref_55_Split/$exit
      -- CP-element group 23: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_Sample/ptr_deref_55_Split/split_req
      -- CP-element group 23: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_Sample/ptr_deref_55_Split/split_ack
      -- CP-element group 23: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_Sample/word_access_start/$entry
      -- CP-element group 23: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_Sample/word_access_start/word_0/$entry
      -- CP-element group 23: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_Sample/word_access_start/word_0/rr
      -- 
    rr_314_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_314_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeModule1_CP_181_elements(23), ack => ptr_deref_55_store_0_req_0); -- 
    writeModule1_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 8,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 32) := "writeModule1_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= writeModule1_CP_181_elements(1) & writeModule1_CP_181_elements(22) & writeModule1_CP_181_elements(25);
      gj_writeModule1_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeModule1_CP_181_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: marked-predecessors 
    -- CP-element group 24: 	26 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	26 
    -- CP-element group 24:  members (5) 
      -- CP-element group 24: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_update_start_
      -- CP-element group 24: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_Update/$entry
      -- CP-element group 24: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_Update/word_access_complete/$entry
      -- CP-element group 24: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_Update/word_access_complete/word_0/$entry
      -- CP-element group 24: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_Update/word_access_complete/word_0/cr
      -- 
    cr_325_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_325_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeModule1_CP_181_elements(24), ack => ptr_deref_55_store_0_req_1); -- 
    writeModule1_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 32) := "writeModule1_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= writeModule1_CP_181_elements(26);
      gj_writeModule1_cp_element_group_24 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeModule1_CP_181_elements(24), clk => clk, reset => reset); --
    end block;
    -- CP-element group 25:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	23 
    -- CP-element group 25: successors 
    -- CP-element group 25: marked-successors 
    -- CP-element group 25: 	4 
    -- CP-element group 25: 	7 
    -- CP-element group 25: 	23 
    -- CP-element group 25:  members (5) 
      -- CP-element group 25: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_sample_completed_
      -- CP-element group 25: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_Sample/$exit
      -- CP-element group 25: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_Sample/word_access_start/$exit
      -- CP-element group 25: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_Sample/word_access_start/word_0/$exit
      -- CP-element group 25: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_Sample/word_access_start/word_0/ra
      -- 
    ra_315_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_55_store_0_ack_0, ack => writeModule1_CP_181_elements(25)); -- 
    -- CP-element group 26:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	31 
    -- CP-element group 26: marked-successors 
    -- CP-element group 26: 	24 
    -- CP-element group 26:  members (5) 
      -- CP-element group 26: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_update_completed_
      -- CP-element group 26: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_Update/$exit
      -- CP-element group 26: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_Update/word_access_complete/$exit
      -- CP-element group 26: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_Update/word_access_complete/word_0/$exit
      -- CP-element group 26: 	 assign_stmt_53_to_assign_stmt_62/ptr_deref_55_Update/word_access_complete/word_0/ca
      -- 
    ca_326_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_55_store_0_ack_1, ack => writeModule1_CP_181_elements(26)); -- 
    -- CP-element group 27:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	1 
    -- CP-element group 27: marked-predecessors 
    -- CP-element group 27: 	29 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 assign_stmt_53_to_assign_stmt_62/BITSEL_u8_u1_61_sample_start_
      -- CP-element group 27: 	 assign_stmt_53_to_assign_stmt_62/BITSEL_u8_u1_61_Sample/$entry
      -- CP-element group 27: 	 assign_stmt_53_to_assign_stmt_62/BITSEL_u8_u1_61_Sample/rr
      -- 
    rr_334_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_334_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeModule1_CP_181_elements(27), ack => BITSEL_u8_u1_61_inst_req_0); -- 
    writeModule1_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 8,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 32) := "writeModule1_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeModule1_CP_181_elements(1) & writeModule1_CP_181_elements(29);
      gj_writeModule1_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeModule1_CP_181_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	5 
    -- CP-element group 28: marked-predecessors 
    -- CP-element group 28: 	30 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 assign_stmt_53_to_assign_stmt_62/BITSEL_u8_u1_61_update_start_
      -- CP-element group 28: 	 assign_stmt_53_to_assign_stmt_62/BITSEL_u8_u1_61_Update/$entry
      -- CP-element group 28: 	 assign_stmt_53_to_assign_stmt_62/BITSEL_u8_u1_61_Update/cr
      -- 
    cr_339_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_339_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeModule1_CP_181_elements(28), ack => BITSEL_u8_u1_61_inst_req_1); -- 
    writeModule1_cp_element_group_28: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 8,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "writeModule1_cp_element_group_28"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeModule1_CP_181_elements(5) & writeModule1_CP_181_elements(30);
      gj_writeModule1_cp_element_group_28 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeModule1_CP_181_elements(28), clk => clk, reset => reset); --
    end block;
    -- CP-element group 29:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29: marked-successors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: 	2 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 assign_stmt_53_to_assign_stmt_62/BITSEL_u8_u1_61_sample_completed_
      -- CP-element group 29: 	 assign_stmt_53_to_assign_stmt_62/BITSEL_u8_u1_61_Sample/$exit
      -- CP-element group 29: 	 assign_stmt_53_to_assign_stmt_62/BITSEL_u8_u1_61_Sample/ra
      -- 
    ra_335_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => BITSEL_u8_u1_61_inst_ack_0, ack => writeModule1_CP_181_elements(29)); -- 
    -- CP-element group 30:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30: marked-successors 
    -- CP-element group 30: 	28 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 assign_stmt_53_to_assign_stmt_62/BITSEL_u8_u1_61_update_completed_
      -- CP-element group 30: 	 assign_stmt_53_to_assign_stmt_62/BITSEL_u8_u1_61_Update/$exit
      -- CP-element group 30: 	 assign_stmt_53_to_assign_stmt_62/BITSEL_u8_u1_61_Update/ca
      -- 
    ca_340_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => BITSEL_u8_u1_61_inst_ack_1, ack => writeModule1_CP_181_elements(30)); -- 
    -- CP-element group 31:  join  transition  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	26 
    -- CP-element group 31: 	16 
    -- CP-element group 31: 	19 
    -- CP-element group 31: 	12 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	36 
    -- CP-element group 31:  members (1) 
      -- CP-element group 31: 	 assign_stmt_53_to_assign_stmt_62/$exit
      -- 
    writeModule1_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 8,1 => 8,2 => 8,3 => 8,4 => 8);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 32) := "writeModule1_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= writeModule1_CP_181_elements(26) & writeModule1_CP_181_elements(16) & writeModule1_CP_181_elements(19) & writeModule1_CP_181_elements(12) & writeModule1_CP_181_elements(30);
      gj_writeModule1_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeModule1_CP_181_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  place  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	2 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 index_update_enable
      -- 
    writeModule1_CP_181_elements(32) <= writeModule1_CP_181_elements(2);
    -- CP-element group 33:  place  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	3 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (1) 
      -- CP-element group 33: 	 address_update_enable
      -- 
    writeModule1_CP_181_elements(33) <= writeModule1_CP_181_elements(3);
    -- CP-element group 34:  place  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	4 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (1) 
      -- CP-element group 34: 	 data_update_enable
      -- 
    writeModule1_CP_181_elements(34) <= writeModule1_CP_181_elements(4);
    -- CP-element group 35:  place  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	5 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 done_update_enable
      -- 
    -- CP-element group 36:  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	31 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 $exit
      -- 
    writeModule1_CP_181_elements(36) <= writeModule1_CP_181_elements(31);
    --  hookup: inputs to control-path 
    writeModule1_CP_181_elements(35) <= done_update_enable;
    -- hookup: output from control-path 
    index_update_enable <= writeModule1_CP_181_elements(32);
    address_update_enable <= writeModule1_CP_181_elements(33);
    data_update_enable <= writeModule1_CP_181_elements(34);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_address_50_resized : std_logic_vector(15 downto 0);
    signal R_address_50_scaled : std_logic_vector(15 downto 0);
    signal array_obj_ref_51_constant_part_of_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_51_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_51_index_partial_sum_1 : std_logic_vector(15 downto 0);
    signal array_obj_ref_51_offset_scale_factor_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_51_offset_scale_factor_1 : std_logic_vector(15 downto 0);
    signal array_obj_ref_51_offset_scale_factor_2 : std_logic_vector(15 downto 0);
    signal array_obj_ref_51_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_51_root_address : std_logic_vector(15 downto 0);
    signal konst_60_wire_constant : std_logic_vector(7 downto 0);
    signal ptr_53 : std_logic_vector(31 downto 0);
    signal ptr_deref_55_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_55_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_55_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_55_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_55_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_55_word_offset_0 : std_logic_vector(15 downto 0);
    signal type_cast_47_resized : std_logic_vector(15 downto 0);
    signal type_cast_47_scaled : std_logic_vector(15 downto 0);
    signal type_cast_47_wire : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    array_obj_ref_51_constant_part_of_offset <= "0000000000000000";
    array_obj_ref_51_offset_scale_factor_0 <= "0100000000000000";
    array_obj_ref_51_offset_scale_factor_1 <= "0100000000000000";
    array_obj_ref_51_offset_scale_factor_2 <= "0000000000000001";
    array_obj_ref_51_resized_base_address <= "0000000000000000";
    konst_60_wire_constant <= "00000000";
    ptr_deref_55_word_offset_0 <= "0000000000000000";
    addr_of_52_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_52_final_reg_req_0;
      addr_of_52_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_52_final_reg_req_1;
      addr_of_52_final_reg_ack_1<= rack(0);
      addr_of_52_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_52_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_51_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ptr_53,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_47_inst
    process(index_buffer) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := index_buffer(7 downto 0);
      type_cast_47_wire <= tmp_var; -- 
    end process;
    -- equivalence array_obj_ref_51_index_0_resize
    process(type_cast_47_wire) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_47_wire;
      ov := iv(15 downto 0);
      type_cast_47_resized <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_51_index_2_rename
    process(R_address_50_resized) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_address_50_resized;
      ov(15 downto 0) := iv;
      R_address_50_scaled <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_51_index_2_resize
    process(address_buffer) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := address_buffer;
      ov := iv(15 downto 0);
      R_address_50_resized <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_51_root_address_inst
    process(array_obj_ref_51_final_offset) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_51_final_offset;
      ov(15 downto 0) := iv;
      array_obj_ref_51_root_address <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_55_addr_0
    process(ptr_deref_55_root_address) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_55_root_address;
      ov(15 downto 0) := iv;
      ptr_deref_55_word_address_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_55_base_resize
    process(ptr_53) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_53;
      ov := iv(15 downto 0);
      ptr_deref_55_resized_base_address <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_55_gather_scatter
    process(data_buffer) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := data_buffer;
      ov(63 downto 0) := iv;
      ptr_deref_55_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_55_root_address_inst
    process(ptr_deref_55_resized_base_address) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_55_resized_base_address;
      ov(15 downto 0) := iv;
      ptr_deref_55_root_address <= ov(15 downto 0);
      --
    end process;
    -- shared split operator group (0) : BITSEL_u8_u1_61_inst 
    ApBitsel_group_0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= index_buffer;
      done_buffer <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= BITSEL_u8_u1_61_inst_req_0;
      BITSEL_u8_u1_61_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= BITSEL_u8_u1_61_inst_req_1;
      BITSEL_u8_u1_61_inst_ack_1 <= ackR_unguarded(0);
      ApBitsel_group_0_gI: SplitGuardInterface generic map(name => "ApBitsel_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApBitsel",
          name => "ApBitsel_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000",
          constant_width => 8,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : array_obj_ref_51_index_0_scale 
    ApIntMul_group_1: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= type_cast_47_resized;
      type_cast_47_scaled <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_51_index_0_scale_req_0;
      array_obj_ref_51_index_0_scale_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_51_index_0_scale_req_1;
      array_obj_ref_51_index_0_scale_ack_1 <= ackR_unguarded(0);
      ApIntMul_group_1_gI: SplitGuardInterface generic map(name => "ApIntMul_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntMul",
          name => "ApIntMul_group_1",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0100000000000000",
          constant_width => 16,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : array_obj_ref_51_index_offset 
    ApIntAdd_group_2: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= array_obj_ref_51_index_partial_sum_1;
      array_obj_ref_51_final_offset <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_51_index_offset_req_0;
      array_obj_ref_51_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_51_index_offset_req_1;
      array_obj_ref_51_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_2_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_2",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- shared split operator group (3) : array_obj_ref_51_index_sum_1 
    ApIntAdd_group_3: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_address_50_scaled & type_cast_47_scaled;
      array_obj_ref_51_index_partial_sum_1 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_51_index_sum_1_req_0;
      array_obj_ref_51_index_sum_1_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_51_index_sum_1_req_1;
      array_obj_ref_51_index_sum_1_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_3_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_3",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- shared store operator group (0) : ptr_deref_55_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(15 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 8);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 6);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_55_store_0_req_0;
      ptr_deref_55_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_55_store_0_req_1;
      ptr_deref_55_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_55_word_address_0;
      data_in <= ptr_deref_55_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 16,
        data_width => 64,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(15 downto 0),
          mdata => memory_space_0_sr_data(63 downto 0),
          mtag => memory_space_0_sr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end writeModule1_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    Concat_input_pipe_pipe_write_data: in std_logic_vector(7 downto 0);
    Concat_input_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    Concat_input_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    Concat_output_pipe_pipe_read_data: out std_logic_vector(7 downto 0);
    Concat_output_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    Concat_output_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(1 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(1 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(31 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(39 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(1 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(127 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(1 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(1 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(31 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(127 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(39 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(1 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(3 downto 0);
  -- declarations related to module concat
  component concat is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(15 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(15 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
      Concat_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      Concat_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Concat_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      Concat_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      Concat_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Concat_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      timer_call_reqs : out  std_logic_vector(0 downto 0);
      timer_call_acks : in   std_logic_vector(0 downto 0);
      timer_call_tag  :  out  std_logic_vector(1 downto 0);
      timer_return_reqs : out  std_logic_vector(0 downto 0);
      timer_return_acks : in   std_logic_vector(0 downto 0);
      timer_return_data : in   std_logic_vector(63 downto 0);
      timer_return_tag :  in   std_logic_vector(1 downto 0);
      concat_core_call_reqs : out  std_logic_vector(0 downto 0);
      concat_core_call_acks : in   std_logic_vector(0 downto 0);
      concat_core_call_data : out  std_logic_vector(63 downto 0);
      concat_core_call_tag  :  out  std_logic_vector(0 downto 0);
      concat_core_return_reqs : out  std_logic_vector(0 downto 0);
      concat_core_return_acks : in   std_logic_vector(0 downto 0);
      concat_core_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module concat
  signal concat_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal concat_tag_out   : std_logic_vector(1 downto 0);
  signal concat_start_req : std_logic;
  signal concat_start_ack : std_logic;
  signal concat_fin_req   : std_logic;
  signal concat_fin_ack : std_logic;
  -- declarations related to module concat_core
  component concat_core is -- 
    generic (tag_length : integer); 
    port ( -- 
      input1_count : in  std_logic_vector(15 downto 0);
      input2_count : in  std_logic_vector(15 downto 0);
      output_size : in  std_logic_vector(31 downto 0);
      readModule1_call_reqs : out  std_logic_vector(0 downto 0);
      readModule1_call_acks : in   std_logic_vector(0 downto 0);
      readModule1_call_data : out  std_logic_vector(39 downto 0);
      readModule1_call_tag  :  out  std_logic_vector(1 downto 0);
      readModule1_return_reqs : out  std_logic_vector(0 downto 0);
      readModule1_return_acks : in   std_logic_vector(0 downto 0);
      readModule1_return_data : in   std_logic_vector(63 downto 0);
      readModule1_return_tag :  in   std_logic_vector(1 downto 0);
      writeModule1_call_reqs : out  std_logic_vector(0 downto 0);
      writeModule1_call_acks : in   std_logic_vector(0 downto 0);
      writeModule1_call_data : out  std_logic_vector(103 downto 0);
      writeModule1_call_tag  :  out  std_logic_vector(0 downto 0);
      writeModule1_return_reqs : out  std_logic_vector(0 downto 0);
      writeModule1_return_acks : in   std_logic_vector(0 downto 0);
      writeModule1_return_data : in   std_logic_vector(0 downto 0);
      writeModule1_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module concat_core
  signal concat_core_input1_count :  std_logic_vector(15 downto 0);
  signal concat_core_input2_count :  std_logic_vector(15 downto 0);
  signal concat_core_output_size :  std_logic_vector(31 downto 0);
  signal concat_core_in_args    : std_logic_vector(63 downto 0);
  signal concat_core_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal concat_core_tag_out   : std_logic_vector(1 downto 0);
  signal concat_core_start_req : std_logic;
  signal concat_core_start_ack : std_logic;
  signal concat_core_fin_req   : std_logic;
  signal concat_core_fin_ack : std_logic;
  -- caller side aggregated signals for module concat_core
  signal concat_core_call_reqs: std_logic_vector(0 downto 0);
  signal concat_core_call_acks: std_logic_vector(0 downto 0);
  signal concat_core_return_reqs: std_logic_vector(0 downto 0);
  signal concat_core_return_acks: std_logic_vector(0 downto 0);
  signal concat_core_call_data: std_logic_vector(63 downto 0);
  signal concat_core_call_tag: std_logic_vector(0 downto 0);
  signal concat_core_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module readModule1
  component readModule1 is -- 
    generic (tag_length : integer); 
    port ( -- 
      index : in  std_logic_vector(7 downto 0);
      address : in  std_logic_vector(31 downto 0);
      data : out  std_logic_vector(63 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(15 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module readModule1
  signal readModule1_index :  std_logic_vector(7 downto 0);
  signal readModule1_address :  std_logic_vector(31 downto 0);
  signal readModule1_data :  std_logic_vector(63 downto 0);
  signal readModule1_in_args    : std_logic_vector(39 downto 0);
  signal readModule1_out_args   : std_logic_vector(63 downto 0);
  signal readModule1_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal readModule1_tag_out   : std_logic_vector(2 downto 0);
  signal readModule1_start_req : std_logic;
  signal readModule1_start_ack : std_logic;
  signal readModule1_fin_req   : std_logic;
  signal readModule1_fin_ack : std_logic;
  -- caller side aggregated signals for module readModule1
  signal readModule1_call_reqs: std_logic_vector(0 downto 0);
  signal readModule1_call_acks: std_logic_vector(0 downto 0);
  signal readModule1_return_reqs: std_logic_vector(0 downto 0);
  signal readModule1_return_acks: std_logic_vector(0 downto 0);
  signal readModule1_call_data: std_logic_vector(39 downto 0);
  signal readModule1_call_tag: std_logic_vector(1 downto 0);
  signal readModule1_return_data: std_logic_vector(63 downto 0);
  signal readModule1_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module timer
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      T : out  std_logic_vector(63 downto 0);
      timer_resp_pipe_read_req : out  std_logic_vector(0 downto 0);
      timer_resp_pipe_read_ack : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_read_data : in   std_logic_vector(63 downto 0);
      timer_req_pipe_write_req : out  std_logic_vector(0 downto 0);
      timer_req_pipe_write_ack : in   std_logic_vector(0 downto 0);
      timer_req_pipe_write_data : out  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timer
  signal timer_T :  std_logic_vector(63 downto 0);
  signal timer_out_args   : std_logic_vector(63 downto 0);
  signal timer_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal timer_tag_out   : std_logic_vector(2 downto 0);
  signal timer_start_req : std_logic;
  signal timer_start_ack : std_logic;
  signal timer_fin_req   : std_logic;
  signal timer_fin_ack : std_logic;
  -- caller side aggregated signals for module timer
  signal timer_call_reqs: std_logic_vector(0 downto 0);
  signal timer_call_acks: std_logic_vector(0 downto 0);
  signal timer_return_reqs: std_logic_vector(0 downto 0);
  signal timer_return_acks: std_logic_vector(0 downto 0);
  signal timer_call_tag: std_logic_vector(1 downto 0);
  signal timer_return_data: std_logic_vector(63 downto 0);
  signal timer_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module timerDaemon
  component timerDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      timer_req_pipe_read_req : out  std_logic_vector(0 downto 0);
      timer_req_pipe_read_ack : in   std_logic_vector(0 downto 0);
      timer_req_pipe_read_data : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_write_req : out  std_logic_vector(0 downto 0);
      timer_resp_pipe_write_ack : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_write_data : out  std_logic_vector(63 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timerDaemon
  signal timerDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal timerDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal timerDaemon_start_req : std_logic;
  signal timerDaemon_start_ack : std_logic;
  signal timerDaemon_fin_req   : std_logic;
  signal timerDaemon_fin_ack : std_logic;
  -- declarations related to module writeModule1
  component writeModule1 is -- 
    generic (tag_length : integer); 
    port ( -- 
      index : in  std_logic_vector(7 downto 0);
      address : in  std_logic_vector(31 downto 0);
      data : in  std_logic_vector(63 downto 0);
      done : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(15 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module writeModule1
  signal writeModule1_index :  std_logic_vector(7 downto 0);
  signal writeModule1_address :  std_logic_vector(31 downto 0);
  signal writeModule1_data :  std_logic_vector(63 downto 0);
  signal writeModule1_done :  std_logic_vector(0 downto 0);
  signal writeModule1_in_args    : std_logic_vector(103 downto 0);
  signal writeModule1_out_args   : std_logic_vector(0 downto 0);
  signal writeModule1_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal writeModule1_tag_out   : std_logic_vector(1 downto 0);
  signal writeModule1_start_req : std_logic;
  signal writeModule1_start_ack : std_logic;
  signal writeModule1_fin_req   : std_logic;
  signal writeModule1_fin_ack : std_logic;
  -- caller side aggregated signals for module writeModule1
  signal writeModule1_call_reqs: std_logic_vector(0 downto 0);
  signal writeModule1_call_acks: std_logic_vector(0 downto 0);
  signal writeModule1_return_reqs: std_logic_vector(0 downto 0);
  signal writeModule1_return_acks: std_logic_vector(0 downto 0);
  signal writeModule1_call_data: std_logic_vector(103 downto 0);
  signal writeModule1_call_tag: std_logic_vector(0 downto 0);
  signal writeModule1_return_data: std_logic_vector(0 downto 0);
  signal writeModule1_return_tag: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Concat_input_pipe
  signal Concat_input_pipe_pipe_read_data: std_logic_vector(7 downto 0);
  signal Concat_input_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal Concat_input_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Concat_output_pipe
  signal Concat_output_pipe_pipe_write_data: std_logic_vector(7 downto 0);
  signal Concat_output_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal Concat_output_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe timer_req
  signal timer_req_pipe_write_data: std_logic_vector(0 downto 0);
  signal timer_req_pipe_write_req: std_logic_vector(0 downto 0);
  signal timer_req_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe timer_req
  signal timer_req_pipe_read_data: std_logic_vector(0 downto 0);
  signal timer_req_pipe_read_req: std_logic_vector(0 downto 0);
  signal timer_req_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe timer_resp
  signal timer_resp_pipe_write_data: std_logic_vector(63 downto 0);
  signal timer_resp_pipe_write_req: std_logic_vector(0 downto 0);
  signal timer_resp_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe timer_resp
  signal timer_resp_pipe_read_data: std_logic_vector(63 downto 0);
  signal timer_resp_pipe_read_req: std_logic_vector(0 downto 0);
  signal timer_resp_pipe_read_ack: std_logic_vector(0 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module concat
  concat_instance:concat-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => concat_start_req,
      start_ack => concat_start_ack,
      fin_req => concat_fin_req,
      fin_ack => concat_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(15 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(19 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(1 downto 0),
      memory_space_0_sr_req => memory_space_0_sr_req(1 downto 1),
      memory_space_0_sr_ack => memory_space_0_sr_ack(1 downto 1),
      memory_space_0_sr_addr => memory_space_0_sr_addr(31 downto 16),
      memory_space_0_sr_data => memory_space_0_sr_data(127 downto 64),
      memory_space_0_sr_tag => memory_space_0_sr_tag(39 downto 20),
      memory_space_0_sc_req => memory_space_0_sc_req(1 downto 1),
      memory_space_0_sc_ack => memory_space_0_sc_ack(1 downto 1),
      memory_space_0_sc_tag => memory_space_0_sc_tag(3 downto 2),
      Concat_input_pipe_pipe_read_req => Concat_input_pipe_pipe_read_req(0 downto 0),
      Concat_input_pipe_pipe_read_ack => Concat_input_pipe_pipe_read_ack(0 downto 0),
      Concat_input_pipe_pipe_read_data => Concat_input_pipe_pipe_read_data(7 downto 0),
      Concat_output_pipe_pipe_write_req => Concat_output_pipe_pipe_write_req(0 downto 0),
      Concat_output_pipe_pipe_write_ack => Concat_output_pipe_pipe_write_ack(0 downto 0),
      Concat_output_pipe_pipe_write_data => Concat_output_pipe_pipe_write_data(7 downto 0),
      timer_call_reqs => timer_call_reqs(0 downto 0),
      timer_call_acks => timer_call_acks(0 downto 0),
      timer_call_tag => timer_call_tag(1 downto 0),
      timer_return_reqs => timer_return_reqs(0 downto 0),
      timer_return_acks => timer_return_acks(0 downto 0),
      timer_return_data => timer_return_data(63 downto 0),
      timer_return_tag => timer_return_tag(1 downto 0),
      concat_core_call_reqs => concat_core_call_reqs(0 downto 0),
      concat_core_call_acks => concat_core_call_acks(0 downto 0),
      concat_core_call_data => concat_core_call_data(63 downto 0),
      concat_core_call_tag => concat_core_call_tag(0 downto 0),
      concat_core_return_reqs => concat_core_return_reqs(0 downto 0),
      concat_core_return_acks => concat_core_return_acks(0 downto 0),
      concat_core_return_tag => concat_core_return_tag(0 downto 0),
      tag_in => concat_tag_in,
      tag_out => concat_tag_out-- 
    ); -- 
  -- module will be run forever 
  concat_tag_in <= (others => '0');
  concat_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => concat_start_req, start_ack => concat_start_ack,  fin_req => concat_fin_req,  fin_ack => concat_fin_ack);
  -- module concat_core
  concat_core_input1_count <= concat_core_in_args(63 downto 48);
  concat_core_input2_count <= concat_core_in_args(47 downto 32);
  concat_core_output_size <= concat_core_in_args(31 downto 0);
  -- call arbiter for module concat_core
  concat_core_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => concat_core_call_reqs,
      call_acks => concat_core_call_acks,
      return_reqs => concat_core_return_reqs,
      return_acks => concat_core_return_acks,
      call_data  => concat_core_call_data,
      call_tag  => concat_core_call_tag,
      return_tag  => concat_core_return_tag,
      call_mtag => concat_core_tag_in,
      return_mtag => concat_core_tag_out,
      call_mreq => concat_core_start_req,
      call_mack => concat_core_start_ack,
      return_mreq => concat_core_fin_req,
      return_mack => concat_core_fin_ack,
      call_mdata => concat_core_in_args,
      clk => clk, 
      reset => reset --
    ); --
  concat_core_instance:concat_core-- 
    generic map(tag_length => 2)
    port map(-- 
      input1_count => concat_core_input1_count,
      input2_count => concat_core_input2_count,
      output_size => concat_core_output_size,
      start_req => concat_core_start_req,
      start_ack => concat_core_start_ack,
      fin_req => concat_core_fin_req,
      fin_ack => concat_core_fin_ack,
      clk => clk,
      reset => reset,
      readModule1_call_reqs => readModule1_call_reqs(0 downto 0),
      readModule1_call_acks => readModule1_call_acks(0 downto 0),
      readModule1_call_data => readModule1_call_data(39 downto 0),
      readModule1_call_tag => readModule1_call_tag(1 downto 0),
      readModule1_return_reqs => readModule1_return_reqs(0 downto 0),
      readModule1_return_acks => readModule1_return_acks(0 downto 0),
      readModule1_return_data => readModule1_return_data(63 downto 0),
      readModule1_return_tag => readModule1_return_tag(1 downto 0),
      writeModule1_call_reqs => writeModule1_call_reqs(0 downto 0),
      writeModule1_call_acks => writeModule1_call_acks(0 downto 0),
      writeModule1_call_data => writeModule1_call_data(103 downto 0),
      writeModule1_call_tag => writeModule1_call_tag(0 downto 0),
      writeModule1_return_reqs => writeModule1_return_reqs(0 downto 0),
      writeModule1_return_acks => writeModule1_return_acks(0 downto 0),
      writeModule1_return_data => writeModule1_return_data(0 downto 0),
      writeModule1_return_tag => writeModule1_return_tag(0 downto 0),
      tag_in => concat_core_tag_in,
      tag_out => concat_core_tag_out-- 
    ); -- 
  -- module readModule1
  readModule1_index <= readModule1_in_args(39 downto 32);
  readModule1_address <= readModule1_in_args(31 downto 0);
  readModule1_out_args <= readModule1_data ;
  -- call arbiter for module readModule1
  readModule1_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 40,
      return_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => readModule1_call_reqs,
      call_acks => readModule1_call_acks,
      return_reqs => readModule1_return_reqs,
      return_acks => readModule1_return_acks,
      call_data  => readModule1_call_data,
      call_tag  => readModule1_call_tag,
      return_tag  => readModule1_return_tag,
      call_mtag => readModule1_tag_in,
      return_mtag => readModule1_tag_out,
      return_data =>readModule1_return_data,
      call_mreq => readModule1_start_req,
      call_mack => readModule1_start_ack,
      return_mreq => readModule1_fin_req,
      return_mack => readModule1_fin_ack,
      call_mdata => readModule1_in_args,
      return_mdata => readModule1_out_args,
      clk => clk, 
      reset => reset --
    ); --
  readModule1_instance:readModule1-- 
    generic map(tag_length => 3)
    port map(-- 
      index => readModule1_index,
      address => readModule1_address,
      data => readModule1_data,
      start_req => readModule1_start_req,
      start_ack => readModule1_start_ack,
      fin_req => readModule1_fin_req,
      fin_ack => readModule1_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(1 downto 1),
      memory_space_0_lr_ack => memory_space_0_lr_ack(1 downto 1),
      memory_space_0_lr_addr => memory_space_0_lr_addr(31 downto 16),
      memory_space_0_lr_tag => memory_space_0_lr_tag(39 downto 20),
      memory_space_0_lc_req => memory_space_0_lc_req(1 downto 1),
      memory_space_0_lc_ack => memory_space_0_lc_ack(1 downto 1),
      memory_space_0_lc_data => memory_space_0_lc_data(127 downto 64),
      memory_space_0_lc_tag => memory_space_0_lc_tag(3 downto 2),
      tag_in => readModule1_tag_in,
      tag_out => readModule1_tag_out-- 
    ); -- 
  -- module timer
  timer_out_args <= timer_T ;
  -- call arbiter for module timer
  timer_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargs", num_reqs => 1,
      return_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => timer_call_reqs,
      call_acks => timer_call_acks,
      return_reqs => timer_return_reqs,
      return_acks => timer_return_acks,
      call_tag  => timer_call_tag,
      return_tag  => timer_return_tag,
      call_mtag => timer_tag_in,
      return_mtag => timer_tag_out,
      return_data =>timer_return_data,
      call_mreq => timer_start_req,
      call_mack => timer_start_ack,
      return_mreq => timer_fin_req,
      return_mack => timer_fin_ack,
      return_mdata => timer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  timer_instance:timer-- 
    generic map(tag_length => 3)
    port map(-- 
      T => timer_T,
      start_req => timer_start_req,
      start_ack => timer_start_ack,
      fin_req => timer_fin_req,
      fin_ack => timer_fin_ack,
      clk => clk,
      reset => reset,
      timer_resp_pipe_read_req => timer_resp_pipe_read_req(0 downto 0),
      timer_resp_pipe_read_ack => timer_resp_pipe_read_ack(0 downto 0),
      timer_resp_pipe_read_data => timer_resp_pipe_read_data(63 downto 0),
      timer_req_pipe_write_req => timer_req_pipe_write_req(0 downto 0),
      timer_req_pipe_write_ack => timer_req_pipe_write_ack(0 downto 0),
      timer_req_pipe_write_data => timer_req_pipe_write_data(0 downto 0),
      tag_in => timer_tag_in,
      tag_out => timer_tag_out-- 
    ); -- 
  -- module timerDaemon
  timerDaemon_instance:timerDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => timerDaemon_start_req,
      start_ack => timerDaemon_start_ack,
      fin_req => timerDaemon_fin_req,
      fin_ack => timerDaemon_fin_ack,
      clk => clk,
      reset => reset,
      timer_req_pipe_read_req => timer_req_pipe_read_req(0 downto 0),
      timer_req_pipe_read_ack => timer_req_pipe_read_ack(0 downto 0),
      timer_req_pipe_read_data => timer_req_pipe_read_data(0 downto 0),
      timer_resp_pipe_write_req => timer_resp_pipe_write_req(0 downto 0),
      timer_resp_pipe_write_ack => timer_resp_pipe_write_ack(0 downto 0),
      timer_resp_pipe_write_data => timer_resp_pipe_write_data(63 downto 0),
      tag_in => timerDaemon_tag_in,
      tag_out => timerDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  timerDaemon_tag_in <= (others => '0');
  timerDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => timerDaemon_start_req, start_ack => timerDaemon_start_ack,  fin_req => timerDaemon_fin_req,  fin_ack => timerDaemon_fin_ack);
  -- module writeModule1
  writeModule1_index <= writeModule1_in_args(103 downto 96);
  writeModule1_address <= writeModule1_in_args(95 downto 64);
  writeModule1_data <= writeModule1_in_args(63 downto 0);
  writeModule1_out_args <= writeModule1_done ;
  -- call arbiter for module writeModule1
  writeModule1_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 104,
      return_data_width => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => writeModule1_call_reqs,
      call_acks => writeModule1_call_acks,
      return_reqs => writeModule1_return_reqs,
      return_acks => writeModule1_return_acks,
      call_data  => writeModule1_call_data,
      call_tag  => writeModule1_call_tag,
      return_tag  => writeModule1_return_tag,
      call_mtag => writeModule1_tag_in,
      return_mtag => writeModule1_tag_out,
      return_data =>writeModule1_return_data,
      call_mreq => writeModule1_start_req,
      call_mack => writeModule1_start_ack,
      return_mreq => writeModule1_fin_req,
      return_mack => writeModule1_fin_ack,
      call_mdata => writeModule1_in_args,
      return_mdata => writeModule1_out_args,
      clk => clk, 
      reset => reset --
    ); --
  writeModule1_instance:writeModule1-- 
    generic map(tag_length => 2)
    port map(-- 
      index => writeModule1_index,
      address => writeModule1_address,
      data => writeModule1_data,
      done => writeModule1_done,
      start_req => writeModule1_start_req,
      start_ack => writeModule1_start_ack,
      fin_req => writeModule1_fin_req,
      fin_ack => writeModule1_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(15 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(63 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(19 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(1 downto 0),
      tag_in => writeModule1_tag_in,
      tag_out => writeModule1_tag_out-- 
    ); -- 
  Concat_input_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Concat_input_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Concat_input_pipe_pipe_read_req,
      read_ack => Concat_input_pipe_pipe_read_ack,
      read_data => Concat_input_pipe_pipe_read_data,
      write_req => Concat_input_pipe_pipe_write_req,
      write_ack => Concat_input_pipe_pipe_write_ack,
      write_data => Concat_input_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Concat_output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Concat_output_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Concat_output_pipe_pipe_read_req,
      read_ack => Concat_output_pipe_pipe_read_ack,
      read_data => Concat_output_pipe_pipe_read_data,
      write_req => Concat_output_pipe_pipe_write_req,
      write_ack => Concat_output_pipe_pipe_write_ack,
      write_data => Concat_output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  timer_req_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe timer_req",
      num_reads => 1,
      num_writes => 1,
      data_width => 1,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => timer_req_pipe_read_req,
      read_ack => timer_req_pipe_read_ack,
      read_data => timer_req_pipe_read_data,
      write_req => timer_req_pipe_write_req,
      write_ack => timer_req_pipe_write_ack,
      write_data => timer_req_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  timer_resp_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe timer_resp",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => timer_resp_pipe_read_req,
      read_ack => timer_resp_pipe_read_ack,
      read_data => timer_resp_pipe_read_data,
      write_req => timer_resp_pipe_write_req,
      write_ack => timer_resp_pipe_write_ack,
      write_data => timer_resp_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  MemorySpace_memory_space_0: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 2,
      num_stores => 2,
      addr_width => 16,
      data_width => 64,
      tag_width => 2,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 16,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
