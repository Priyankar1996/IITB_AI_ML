-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity fill_T is -- 
  generic (tag_length : integer); 
  port ( -- 
    addr : in  std_logic_vector(63 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(255 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(2 downto 0);
    maxpool_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity fill_T;
architecture fill_T_arch of fill_T is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal addr_buffer :  std_logic_vector(63 downto 0);
  signal addr_update_enable: Boolean;
  -- output port buffer signals
  signal fill_T_CP_0_start: Boolean;
  signal fill_T_CP_0_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_maxpool_input_pipe_35_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_35_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_35_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_35_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_39_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_39_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_39_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_39_inst_ack_1 : boolean;
  signal CONCAT_u8_u16_40_inst_req_0 : boolean;
  signal CONCAT_u8_u16_40_inst_ack_0 : boolean;
  signal CONCAT_u8_u16_40_inst_req_1 : boolean;
  signal CONCAT_u8_u16_40_inst_ack_1 : boolean;
  signal CONCAT_u240_u256_47_inst_req_0 : boolean;
  signal CONCAT_u240_u256_47_inst_ack_0 : boolean;
  signal CONCAT_u240_u256_47_inst_req_1 : boolean;
  signal CONCAT_u240_u256_47_inst_ack_1 : boolean;
  signal if_stmt_49_branch_req_0 : boolean;
  signal if_stmt_49_branch_ack_1 : boolean;
  signal if_stmt_49_branch_ack_0 : boolean;
  signal phi_stmt_17_req_0 : boolean;
  signal phi_stmt_23_req_1 : boolean;
  signal nmycount_33_22_buf_req_0 : boolean;
  signal nmycount_33_22_buf_ack_0 : boolean;
  signal nmycount_33_22_buf_req_1 : boolean;
  signal nmycount_33_22_buf_ack_1 : boolean;
  signal phi_stmt_17_req_1 : boolean;
  signal ninput_word_48_25_buf_req_0 : boolean;
  signal ninput_word_48_25_buf_ack_0 : boolean;
  signal ninput_word_48_25_buf_req_1 : boolean;
  signal ninput_word_48_25_buf_ack_1 : boolean;
  signal phi_stmt_23_req_0 : boolean;
  signal phi_stmt_17_ack_0 : boolean;
  signal phi_stmt_23_ack_0 : boolean;
  signal array_obj_ref_62_index_offset_req_0 : boolean;
  signal array_obj_ref_62_index_offset_ack_0 : boolean;
  signal array_obj_ref_62_index_offset_req_1 : boolean;
  signal array_obj_ref_62_index_offset_ack_1 : boolean;
  signal addr_of_63_final_reg_req_0 : boolean;
  signal addr_of_63_final_reg_ack_0 : boolean;
  signal addr_of_63_final_reg_req_1 : boolean;
  signal addr_of_63_final_reg_ack_1 : boolean;
  signal ptr_deref_66_store_0_req_0 : boolean;
  signal ptr_deref_66_store_0_ack_0 : boolean;
  signal ptr_deref_66_store_0_req_1 : boolean;
  signal ptr_deref_66_store_0_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "fill_T_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 64) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(63 downto 0) <= addr;
  addr_buffer <= in_buffer_data_out(63 downto 0);
  in_buffer_data_in(tag_length + 63 downto 64) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 63 downto 64);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  fill_T_CP_0_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "fill_T_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= fill_T_CP_0_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= fill_T_CP_0_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= fill_T_CP_0_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  fill_T_CP_0: Block -- control-path 
    signal fill_T_CP_0_elements: BooleanArray(33 downto 0);
    -- 
  begin -- 
    fill_T_CP_0_elements(0) <= fill_T_CP_0_start;
    fill_T_CP_0_symbol <= fill_T_CP_0_elements(33);
    -- CP-element group 0:  branch  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	12 
    -- CP-element group 0:  members (5) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_15/$entry
      -- CP-element group 0: 	 branch_block_stmt_15/branch_block_stmt_15__entry__
      -- CP-element group 0: 	 branch_block_stmt_15/merge_stmt_16__entry__
      -- CP-element group 0: 	 branch_block_stmt_15/merge_stmt_16_dead_link/$entry
      -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	26 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	7 
    -- CP-element group 1: 	2 
    -- CP-element group 1: 	9 
    -- CP-element group 1:  members (12) 
      -- CP-element group 1: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/RPIPE_maxpool_input_pipe_35_Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/CONCAT_u8_u16_40_update_start_
      -- CP-element group 1: 	 branch_block_stmt_15/merge_stmt_16__exit__
      -- CP-element group 1: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48__entry__
      -- CP-element group 1: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/$entry
      -- CP-element group 1: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/RPIPE_maxpool_input_pipe_35_sample_start_
      -- CP-element group 1: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/RPIPE_maxpool_input_pipe_35_Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/CONCAT_u8_u16_40_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/CONCAT_u8_u16_40_Update/cr
      -- CP-element group 1: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/CONCAT_u240_u256_47_update_start_
      -- CP-element group 1: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/CONCAT_u240_u256_47_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/CONCAT_u240_u256_47_Update/cr
      -- 
    rr_24_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_24_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(1), ack => RPIPE_maxpool_input_pipe_35_inst_req_0); -- 
    cr_57_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_57_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(1), ack => CONCAT_u8_u16_40_inst_req_1); -- 
    cr_71_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_71_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(1), ack => CONCAT_u240_u256_47_inst_req_1); -- 
    fill_T_CP_0_elements(1) <= fill_T_CP_0_elements(26);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/RPIPE_maxpool_input_pipe_35_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/RPIPE_maxpool_input_pipe_35_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/RPIPE_maxpool_input_pipe_35_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/RPIPE_maxpool_input_pipe_35_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/RPIPE_maxpool_input_pipe_35_update_start_
      -- CP-element group 2: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/RPIPE_maxpool_input_pipe_35_Sample/$exit
      -- 
    ra_25_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_35_inst_ack_0, ack => fill_T_CP_0_elements(2)); -- 
    cr_29_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_29_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(2), ack => RPIPE_maxpool_input_pipe_35_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/RPIPE_maxpool_input_pipe_35_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/RPIPE_maxpool_input_pipe_35_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/RPIPE_maxpool_input_pipe_35_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/RPIPE_maxpool_input_pipe_39_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/RPIPE_maxpool_input_pipe_39_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/RPIPE_maxpool_input_pipe_39_Sample/rr
      -- 
    ca_30_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_35_inst_ack_1, ack => fill_T_CP_0_elements(3)); -- 
    rr_42_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_42_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(3), ack => RPIPE_maxpool_input_pipe_39_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/RPIPE_maxpool_input_pipe_39_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/RPIPE_maxpool_input_pipe_39_update_start_
      -- CP-element group 4: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/RPIPE_maxpool_input_pipe_39_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/RPIPE_maxpool_input_pipe_39_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/RPIPE_maxpool_input_pipe_39_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/RPIPE_maxpool_input_pipe_39_Update/cr
      -- 
    ra_43_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_39_inst_ack_0, ack => fill_T_CP_0_elements(4)); -- 
    cr_47_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_47_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(4), ack => RPIPE_maxpool_input_pipe_39_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/CONCAT_u8_u16_40_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/RPIPE_maxpool_input_pipe_39_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/RPIPE_maxpool_input_pipe_39_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/RPIPE_maxpool_input_pipe_39_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/CONCAT_u8_u16_40_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/CONCAT_u8_u16_40_Sample/rr
      -- 
    ca_48_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_39_inst_ack_1, ack => fill_T_CP_0_elements(5)); -- 
    rr_52_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_52_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(5), ack => CONCAT_u8_u16_40_inst_req_0); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/CONCAT_u8_u16_40_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/CONCAT_u8_u16_40_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/CONCAT_u8_u16_40_Sample/ra
      -- 
    ra_53_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u8_u16_40_inst_ack_0, ack => fill_T_CP_0_elements(6)); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	1 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/CONCAT_u8_u16_40_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/CONCAT_u8_u16_40_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/CONCAT_u8_u16_40_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/CONCAT_u240_u256_47_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/CONCAT_u240_u256_47_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/CONCAT_u240_u256_47_Sample/rr
      -- 
    ca_58_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u8_u16_40_inst_ack_1, ack => fill_T_CP_0_elements(7)); -- 
    rr_66_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_66_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(7), ack => CONCAT_u240_u256_47_inst_req_0); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/CONCAT_u240_u256_47_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/CONCAT_u240_u256_47_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/CONCAT_u240_u256_47_Sample/ra
      -- 
    ra_67_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u240_u256_47_inst_ack_0, ack => fill_T_CP_0_elements(8)); -- 
    -- CP-element group 9:  branch  transition  place  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	1 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (27) 
      -- CP-element group 9: 	 branch_block_stmt_15/if_stmt_49_dead_link/$entry
      -- CP-element group 9: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48__exit__
      -- CP-element group 9: 	 branch_block_stmt_15/if_stmt_49__entry__
      -- CP-element group 9: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/$exit
      -- CP-element group 9: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/CONCAT_u240_u256_47_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/CONCAT_u240_u256_47_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_15/assign_stmt_33_to_assign_stmt_48/CONCAT_u240_u256_47_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_15/if_stmt_49_eval_test/$entry
      -- CP-element group 9: 	 branch_block_stmt_15/if_stmt_49_eval_test/$exit
      -- CP-element group 9: 	 branch_block_stmt_15/if_stmt_49_eval_test/ULT_u4_u1_52/$entry
      -- CP-element group 9: 	 branch_block_stmt_15/if_stmt_49_eval_test/ULT_u4_u1_52/$exit
      -- CP-element group 9: 	 branch_block_stmt_15/if_stmt_49_eval_test/ULT_u4_u1_52/ULT_u4_u1_52_inputs/$entry
      -- CP-element group 9: 	 branch_block_stmt_15/if_stmt_49_eval_test/ULT_u4_u1_52/ULT_u4_u1_52_inputs/$exit
      -- CP-element group 9: 	 branch_block_stmt_15/if_stmt_49_eval_test/ULT_u4_u1_52/SplitProtocol/$entry
      -- CP-element group 9: 	 branch_block_stmt_15/if_stmt_49_eval_test/ULT_u4_u1_52/SplitProtocol/$exit
      -- CP-element group 9: 	 branch_block_stmt_15/if_stmt_49_eval_test/ULT_u4_u1_52/SplitProtocol/Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_15/if_stmt_49_eval_test/ULT_u4_u1_52/SplitProtocol/Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_15/if_stmt_49_eval_test/ULT_u4_u1_52/SplitProtocol/Sample/rr
      -- CP-element group 9: 	 branch_block_stmt_15/if_stmt_49_eval_test/ULT_u4_u1_52/SplitProtocol/Sample/ra
      -- CP-element group 9: 	 branch_block_stmt_15/if_stmt_49_eval_test/ULT_u4_u1_52/SplitProtocol/Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_15/if_stmt_49_eval_test/ULT_u4_u1_52/SplitProtocol/Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_15/if_stmt_49_eval_test/ULT_u4_u1_52/SplitProtocol/Update/cr
      -- CP-element group 9: 	 branch_block_stmt_15/if_stmt_49_eval_test/ULT_u4_u1_52/SplitProtocol/Update/ca
      -- CP-element group 9: 	 branch_block_stmt_15/if_stmt_49_eval_test/branch_req
      -- CP-element group 9: 	 branch_block_stmt_15/ULT_u4_u1_52_place
      -- CP-element group 9: 	 branch_block_stmt_15/if_stmt_49_if_link/$entry
      -- CP-element group 9: 	 branch_block_stmt_15/if_stmt_49_else_link/$entry
      -- 
    ca_72_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u240_u256_47_inst_ack_1, ack => fill_T_CP_0_elements(9)); -- 
    branch_req_99_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_99_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(9), ack => if_stmt_49_branch_req_0); -- 
    -- CP-element group 10:  fork  transition  place  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	20 
    -- CP-element group 10: 	19 
    -- CP-element group 10: 	17 
    -- CP-element group 10: 	16 
    -- CP-element group 10:  members (18) 
      -- CP-element group 10: 	 branch_block_stmt_15/if_stmt_49_if_link/$exit
      -- CP-element group 10: 	 branch_block_stmt_15/if_stmt_49_if_link/if_choice_transition
      -- CP-element group 10: 	 branch_block_stmt_15/loopback
      -- CP-element group 10: 	 branch_block_stmt_15/loopback_PhiReq/$entry
      -- CP-element group 10: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_17/$entry
      -- CP-element group 10: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_17/phi_stmt_17_sources/$entry
      -- CP-element group 10: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_17/phi_stmt_17_sources/Interlock/$entry
      -- CP-element group 10: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_17/phi_stmt_17_sources/Interlock/Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_17/phi_stmt_17_sources/Interlock/Sample/req
      -- CP-element group 10: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_17/phi_stmt_17_sources/Interlock/Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_17/phi_stmt_17_sources/Interlock/Update/req
      -- CP-element group 10: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_23/$entry
      -- CP-element group 10: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_23/phi_stmt_23_sources/$entry
      -- CP-element group 10: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_23/phi_stmt_23_sources/Interlock/$entry
      -- CP-element group 10: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_23/phi_stmt_23_sources/Interlock/Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_23/phi_stmt_23_sources/Interlock/Sample/req
      -- CP-element group 10: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_23/phi_stmt_23_sources/Interlock/Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_23/phi_stmt_23_sources/Interlock/Update/req
      -- 
    if_choice_transition_104_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_49_branch_ack_1, ack => fill_T_CP_0_elements(10)); -- 
    req_148_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_148_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(10), ack => nmycount_33_22_buf_req_0); -- 
    req_153_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_153_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(10), ack => nmycount_33_22_buf_req_1); -- 
    req_168_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_168_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(10), ack => ninput_word_48_25_buf_req_0); -- 
    req_173_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_173_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(10), ack => ninput_word_48_25_buf_req_1); -- 
    -- CP-element group 11:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	32 
    -- CP-element group 11: 	27 
    -- CP-element group 11: 	28 
    -- CP-element group 11: 	30 
    -- CP-element group 11:  members (30) 
      -- CP-element group 11: 	 branch_block_stmt_15/$exit
      -- CP-element group 11: 	 branch_block_stmt_15/branch_block_stmt_15__exit__
      -- CP-element group 11: 	 branch_block_stmt_15/if_stmt_49__exit__
      -- CP-element group 11: 	 branch_block_stmt_15/if_stmt_49_else_link/$exit
      -- CP-element group 11: 	 branch_block_stmt_15/if_stmt_49_else_link/else_choice_transition
      -- CP-element group 11: 	 assign_stmt_64_to_assign_stmt_68/$entry
      -- CP-element group 11: 	 assign_stmt_64_to_assign_stmt_68/addr_of_63_update_start_
      -- CP-element group 11: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_index_resized_1
      -- CP-element group 11: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_index_scaled_1
      -- CP-element group 11: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_index_computed_1
      -- CP-element group 11: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_index_resize_1/$entry
      -- CP-element group 11: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_index_resize_1/$exit
      -- CP-element group 11: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_index_resize_1/index_resize_req
      -- CP-element group 11: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_index_resize_1/index_resize_ack
      -- CP-element group 11: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_index_scale_1/$entry
      -- CP-element group 11: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_index_scale_1/$exit
      -- CP-element group 11: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_index_scale_1/scale_rename_req
      -- CP-element group 11: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_index_scale_1/scale_rename_ack
      -- CP-element group 11: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_final_index_sum_regn_update_start
      -- CP-element group 11: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_final_index_sum_regn_Sample/$entry
      -- CP-element group 11: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_final_index_sum_regn_Sample/req
      -- CP-element group 11: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_final_index_sum_regn_Update/$entry
      -- CP-element group 11: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_final_index_sum_regn_Update/req
      -- CP-element group 11: 	 assign_stmt_64_to_assign_stmt_68/addr_of_63_complete/$entry
      -- CP-element group 11: 	 assign_stmt_64_to_assign_stmt_68/addr_of_63_complete/req
      -- CP-element group 11: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_update_start_
      -- CP-element group 11: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_Update/$entry
      -- CP-element group 11: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_Update/word_access_complete/$entry
      -- CP-element group 11: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_Update/word_access_complete/word_0/$entry
      -- CP-element group 11: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_Update/word_access_complete/word_0/cr
      -- 
    else_choice_transition_108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_49_branch_ack_0, ack => fill_T_CP_0_elements(11)); -- 
    req_209_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_209_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(11), ack => array_obj_ref_62_index_offset_req_0); -- 
    req_214_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_214_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(11), ack => array_obj_ref_62_index_offset_req_1); -- 
    req_229_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_229_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(11), ack => addr_of_63_final_reg_req_1); -- 
    cr_279_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_279_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(11), ack => ptr_deref_66_store_0_req_1); -- 
    -- CP-element group 12:  fork  transition  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	0 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	14 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (5) 
      -- CP-element group 12: 	 branch_block_stmt_15/merge_stmt_16__entry___PhiReq/$entry
      -- CP-element group 12: 	 branch_block_stmt_15/merge_stmt_16__entry___PhiReq/phi_stmt_17/$entry
      -- CP-element group 12: 	 branch_block_stmt_15/merge_stmt_16__entry___PhiReq/phi_stmt_17/phi_stmt_17_sources/$entry
      -- CP-element group 12: 	 branch_block_stmt_15/merge_stmt_16__entry___PhiReq/phi_stmt_23/$entry
      -- CP-element group 12: 	 branch_block_stmt_15/merge_stmt_16__entry___PhiReq/phi_stmt_23/phi_stmt_23_sources/$entry
      -- 
    fill_T_CP_0_elements(12) <= fill_T_CP_0_elements(0);
    -- CP-element group 13:  transition  output  delay-element  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	15 
    -- CP-element group 13:  members (4) 
      -- CP-element group 13: 	 branch_block_stmt_15/merge_stmt_16__entry___PhiReq/phi_stmt_17/$exit
      -- CP-element group 13: 	 branch_block_stmt_15/merge_stmt_16__entry___PhiReq/phi_stmt_17/phi_stmt_17_sources/$exit
      -- CP-element group 13: 	 branch_block_stmt_15/merge_stmt_16__entry___PhiReq/phi_stmt_17/phi_stmt_17_sources/type_cast_21_konst_delay_trans
      -- CP-element group 13: 	 branch_block_stmt_15/merge_stmt_16__entry___PhiReq/phi_stmt_17/phi_stmt_17_req
      -- 
    phi_stmt_17_req_124_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_17_req_124_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(13), ack => phi_stmt_17_req_0); -- 
    -- Element group fill_T_CP_0_elements(13) is a control-delay.
    cp_element_13_delay: control_delay_element  generic map(name => " 13_delay", delay_value => 1)  port map(req => fill_T_CP_0_elements(12), ack => fill_T_CP_0_elements(13), clk => clk, reset =>reset);
    -- CP-element group 14:  transition  output  delay-element  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	12 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (4) 
      -- CP-element group 14: 	 branch_block_stmt_15/merge_stmt_16__entry___PhiReq/phi_stmt_23/$exit
      -- CP-element group 14: 	 branch_block_stmt_15/merge_stmt_16__entry___PhiReq/phi_stmt_23/phi_stmt_23_sources/$exit
      -- CP-element group 14: 	 branch_block_stmt_15/merge_stmt_16__entry___PhiReq/phi_stmt_23/phi_stmt_23_sources/type_cast_27_konst_delay_trans
      -- CP-element group 14: 	 branch_block_stmt_15/merge_stmt_16__entry___PhiReq/phi_stmt_23/phi_stmt_23_req
      -- 
    phi_stmt_23_req_132_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_23_req_132_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(14), ack => phi_stmt_23_req_1); -- 
    -- Element group fill_T_CP_0_elements(14) is a control-delay.
    cp_element_14_delay: control_delay_element  generic map(name => " 14_delay", delay_value => 1)  port map(req => fill_T_CP_0_elements(12), ack => fill_T_CP_0_elements(14), clk => clk, reset =>reset);
    -- CP-element group 15:  join  transition  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: 	13 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	23 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_15/merge_stmt_16__entry___PhiReq/$exit
      -- 
    fill_T_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 26) := "fill_T_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= fill_T_CP_0_elements(14) & fill_T_CP_0_elements(13);
      gj_fill_T_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => fill_T_CP_0_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	10 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	18 
    -- CP-element group 16:  members (2) 
      -- CP-element group 16: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_17/phi_stmt_17_sources/Interlock/Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_17/phi_stmt_17_sources/Interlock/Sample/ack
      -- 
    ack_149_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmycount_33_22_buf_ack_0, ack => fill_T_CP_0_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	10 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (2) 
      -- CP-element group 17: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_17/phi_stmt_17_sources/Interlock/Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_17/phi_stmt_17_sources/Interlock/Update/ack
      -- 
    ack_154_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmycount_33_22_buf_ack_1, ack => fill_T_CP_0_elements(17)); -- 
    -- CP-element group 18:  join  transition  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: 	16 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	22 
    -- CP-element group 18:  members (4) 
      -- CP-element group 18: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_17/$exit
      -- CP-element group 18: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_17/phi_stmt_17_sources/$exit
      -- CP-element group 18: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_17/phi_stmt_17_sources/Interlock/$exit
      -- CP-element group 18: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_17/phi_stmt_17_req
      -- 
    phi_stmt_17_req_155_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_17_req_155_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(18), ack => phi_stmt_17_req_1); -- 
    fill_T_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 26) := "fill_T_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= fill_T_CP_0_elements(17) & fill_T_CP_0_elements(16);
      gj_fill_T_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => fill_T_CP_0_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	10 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	21 
    -- CP-element group 19:  members (2) 
      -- CP-element group 19: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_23/phi_stmt_23_sources/Interlock/Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_23/phi_stmt_23_sources/Interlock/Sample/ack
      -- 
    ack_169_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ninput_word_48_25_buf_ack_0, ack => fill_T_CP_0_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	10 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_23/phi_stmt_23_sources/Interlock/Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_23/phi_stmt_23_sources/Interlock/Update/ack
      -- 
    ack_174_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ninput_word_48_25_buf_ack_1, ack => fill_T_CP_0_elements(20)); -- 
    -- CP-element group 21:  join  transition  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: 	19 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (4) 
      -- CP-element group 21: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_23/$exit
      -- CP-element group 21: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_23/phi_stmt_23_sources/$exit
      -- CP-element group 21: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_23/phi_stmt_23_sources/Interlock/$exit
      -- CP-element group 21: 	 branch_block_stmt_15/loopback_PhiReq/phi_stmt_23/phi_stmt_23_req
      -- 
    phi_stmt_23_req_175_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_23_req_175_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(21), ack => phi_stmt_23_req_0); -- 
    fill_T_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 26) := "fill_T_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= fill_T_CP_0_elements(20) & fill_T_CP_0_elements(19);
      gj_fill_T_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => fill_T_CP_0_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  join  transition  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: 	18 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (1) 
      -- CP-element group 22: 	 branch_block_stmt_15/loopback_PhiReq/$exit
      -- 
    fill_T_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 26) := "fill_T_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= fill_T_CP_0_elements(21) & fill_T_CP_0_elements(18);
      gj_fill_T_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => fill_T_CP_0_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  merge  fork  transition  place  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	15 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23: 	25 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_15/merge_stmt_16_PhiReqMerge
      -- CP-element group 23: 	 branch_block_stmt_15/merge_stmt_16_PhiAck/$entry
      -- 
    fill_T_CP_0_elements(23) <= OrReduce(fill_T_CP_0_elements(15) & fill_T_CP_0_elements(22));
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	26 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_15/merge_stmt_16_PhiAck/phi_stmt_17_ack
      -- 
    phi_stmt_17_ack_180_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_17_ack_0, ack => fill_T_CP_0_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	23 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 branch_block_stmt_15/merge_stmt_16_PhiAck/phi_stmt_23_ack
      -- 
    phi_stmt_23_ack_181_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_23_ack_0, ack => fill_T_CP_0_elements(25)); -- 
    -- CP-element group 26:  join  transition  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	1 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_15/merge_stmt_16_PhiAck/$exit
      -- 
    fill_T_cp_element_group_26: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 26) := "fill_T_cp_element_group_26"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= fill_T_CP_0_elements(24) & fill_T_CP_0_elements(25);
      gj_fill_T_cp_element_group_26 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => fill_T_CP_0_elements(26), clk => clk, reset => reset); --
    end block;
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	11 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	33 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_final_index_sum_regn_sample_complete
      -- CP-element group 27: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_final_index_sum_regn_Sample/$exit
      -- CP-element group 27: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_final_index_sum_regn_Sample/ack
      -- 
    ack_210_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_62_index_offset_ack_0, ack => fill_T_CP_0_elements(27)); -- 
    -- CP-element group 28:  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	11 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (11) 
      -- CP-element group 28: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_base_plus_offset/$entry
      -- CP-element group 28: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_base_plus_offset/$exit
      -- CP-element group 28: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_base_plus_offset/sum_rename_req
      -- CP-element group 28: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_base_plus_offset/sum_rename_ack
      -- CP-element group 28: 	 assign_stmt_64_to_assign_stmt_68/addr_of_63_sample_start_
      -- CP-element group 28: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_root_address_calculated
      -- CP-element group 28: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_offset_calculated
      -- CP-element group 28: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_final_index_sum_regn_Update/$exit
      -- CP-element group 28: 	 assign_stmt_64_to_assign_stmt_68/array_obj_ref_62_final_index_sum_regn_Update/ack
      -- CP-element group 28: 	 assign_stmt_64_to_assign_stmt_68/addr_of_63_request/$entry
      -- CP-element group 28: 	 assign_stmt_64_to_assign_stmt_68/addr_of_63_request/req
      -- 
    ack_215_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_62_index_offset_ack_1, ack => fill_T_CP_0_elements(28)); -- 
    req_224_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_224_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(28), ack => addr_of_63_final_reg_req_0); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 assign_stmt_64_to_assign_stmt_68/addr_of_63_sample_completed_
      -- CP-element group 29: 	 assign_stmt_64_to_assign_stmt_68/addr_of_63_request/$exit
      -- CP-element group 29: 	 assign_stmt_64_to_assign_stmt_68/addr_of_63_request/ack
      -- 
    ack_225_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_63_final_reg_ack_0, ack => fill_T_CP_0_elements(29)); -- 
    -- CP-element group 30:  join  fork  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	11 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (28) 
      -- CP-element group 30: 	 assign_stmt_64_to_assign_stmt_68/addr_of_63_update_completed_
      -- CP-element group 30: 	 assign_stmt_64_to_assign_stmt_68/addr_of_63_complete/$exit
      -- CP-element group 30: 	 assign_stmt_64_to_assign_stmt_68/addr_of_63_complete/ack
      -- CP-element group 30: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_sample_start_
      -- CP-element group 30: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_base_address_calculated
      -- CP-element group 30: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_word_address_calculated
      -- CP-element group 30: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_root_address_calculated
      -- CP-element group 30: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_base_address_resized
      -- CP-element group 30: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_base_addr_resize/$entry
      -- CP-element group 30: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_base_addr_resize/$exit
      -- CP-element group 30: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_base_addr_resize/base_resize_req
      -- CP-element group 30: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_base_addr_resize/base_resize_ack
      -- CP-element group 30: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_base_plus_offset/$entry
      -- CP-element group 30: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_base_plus_offset/$exit
      -- CP-element group 30: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_base_plus_offset/sum_rename_req
      -- CP-element group 30: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_base_plus_offset/sum_rename_ack
      -- CP-element group 30: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_word_addrgen/$entry
      -- CP-element group 30: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_word_addrgen/$exit
      -- CP-element group 30: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_word_addrgen/root_register_req
      -- CP-element group 30: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_word_addrgen/root_register_ack
      -- CP-element group 30: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_Sample/$entry
      -- CP-element group 30: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_Sample/ptr_deref_66_Split/$entry
      -- CP-element group 30: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_Sample/ptr_deref_66_Split/$exit
      -- CP-element group 30: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_Sample/ptr_deref_66_Split/split_req
      -- CP-element group 30: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_Sample/ptr_deref_66_Split/split_ack
      -- CP-element group 30: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_Sample/word_access_start/$entry
      -- CP-element group 30: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_Sample/word_access_start/word_0/$entry
      -- CP-element group 30: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_Sample/word_access_start/word_0/rr
      -- 
    ack_230_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_63_final_reg_ack_1, ack => fill_T_CP_0_elements(30)); -- 
    rr_268_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_268_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => fill_T_CP_0_elements(30), ack => ptr_deref_66_store_0_req_0); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (5) 
      -- CP-element group 31: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_sample_completed_
      -- CP-element group 31: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_Sample/$exit
      -- CP-element group 31: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_Sample/word_access_start/$exit
      -- CP-element group 31: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_Sample/word_access_start/word_0/$exit
      -- CP-element group 31: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_Sample/word_access_start/word_0/ra
      -- 
    ra_269_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_66_store_0_ack_0, ack => fill_T_CP_0_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	11 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (5) 
      -- CP-element group 32: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_update_completed_
      -- CP-element group 32: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_Update/$exit
      -- CP-element group 32: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_Update/word_access_complete/$exit
      -- CP-element group 32: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_Update/word_access_complete/word_0/$exit
      -- CP-element group 32: 	 assign_stmt_64_to_assign_stmt_68/ptr_deref_66_Update/word_access_complete/word_0/ca
      -- 
    ca_280_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_66_store_0_ack_1, ack => fill_T_CP_0_elements(32)); -- 
    -- CP-element group 33:  join  transition  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: 	27 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (2) 
      -- CP-element group 33: 	 $exit
      -- CP-element group 33: 	 assign_stmt_64_to_assign_stmt_68/$exit
      -- 
    fill_T_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 26) := "fill_T_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= fill_T_CP_0_elements(32) & fill_T_CP_0_elements(27);
      gj_fill_T_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => fill_T_CP_0_elements(33), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal RPIPE_maxpool_input_pipe_39_wire : std_logic_vector(7 downto 0);
    signal R_addr_61_resized : std_logic_vector(13 downto 0);
    signal R_addr_61_scaled : std_logic_vector(13 downto 0);
    signal ULT_u4_u1_52_wire : std_logic_vector(0 downto 0);
    signal array_obj_ref_62_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_62_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_62_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_62_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_62_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_62_root_address : std_logic_vector(13 downto 0);
    signal input_word_23 : std_logic_vector(255 downto 0);
    signal konst_31_wire_constant : std_logic_vector(3 downto 0);
    signal konst_51_wire_constant : std_logic_vector(3 downto 0);
    signal mycount_17 : std_logic_vector(3 downto 0);
    signal ninput_word_48 : std_logic_vector(255 downto 0);
    signal ninput_word_48_25_buffered : std_logic_vector(255 downto 0);
    signal nmycount_33 : std_logic_vector(3 downto 0);
    signal nmycount_33_22_buffered : std_logic_vector(3 downto 0);
    signal ptr_64 : std_logic_vector(31 downto 0);
    signal ptr_deref_66_data_0 : std_logic_vector(255 downto 0);
    signal ptr_deref_66_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_66_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_66_wire : std_logic_vector(255 downto 0);
    signal ptr_deref_66_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_66_word_offset_0 : std_logic_vector(13 downto 0);
    signal slice_45_wire : std_logic_vector(239 downto 0);
    signal type_cast_21_wire_constant : std_logic_vector(3 downto 0);
    signal type_cast_27_wire_constant : std_logic_vector(255 downto 0);
    signal val1_36 : std_logic_vector(7 downto 0);
    signal val_41 : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_62_constant_part_of_offset <= "00000000000000";
    array_obj_ref_62_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_62_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_62_resized_base_address <= "00000000000000";
    konst_31_wire_constant <= "0001";
    konst_51_wire_constant <= "1111";
    ptr_deref_66_word_offset_0 <= "00000000000000";
    type_cast_21_wire_constant <= "0000";
    type_cast_27_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    phi_stmt_17: Block -- phi operator 
      signal idata: std_logic_vector(7 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_21_wire_constant & nmycount_33_22_buffered;
      req <= phi_stmt_17_req_0 & phi_stmt_17_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_17",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 4) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_17_ack_0,
          idata => idata,
          odata => mycount_17,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_17
    phi_stmt_23: Block -- phi operator 
      signal idata: std_logic_vector(511 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= ninput_word_48_25_buffered & type_cast_27_wire_constant;
      req <= phi_stmt_23_req_0 & phi_stmt_23_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_23",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 256) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_23_ack_0,
          idata => idata,
          odata => input_word_23,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_23
    -- flow-through slice operator slice_45_inst
    slice_45_wire <= input_word_23(239 downto 0);
    addr_of_63_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_63_final_reg_req_0;
      addr_of_63_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_63_final_reg_req_1;
      addr_of_63_final_reg_ack_1<= rack(0);
      addr_of_63_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_63_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_62_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ptr_64,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    ninput_word_48_25_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= ninput_word_48_25_buf_req_0;
      ninput_word_48_25_buf_ack_0<= wack(0);
      rreq(0) <= ninput_word_48_25_buf_req_1;
      ninput_word_48_25_buf_ack_1<= rack(0);
      ninput_word_48_25_buf : InterlockBuffer generic map ( -- 
        name => "ninput_word_48_25_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 256,
        out_data_width => 256,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ninput_word_48,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ninput_word_48_25_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nmycount_33_22_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nmycount_33_22_buf_req_0;
      nmycount_33_22_buf_ack_0<= wack(0);
      rreq(0) <= nmycount_33_22_buf_req_1;
      nmycount_33_22_buf_ack_1<= rack(0);
      nmycount_33_22_buf : InterlockBuffer generic map ( -- 
        name => "nmycount_33_22_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 4,
        out_data_width => 4,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nmycount_33,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nmycount_33_22_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_62_index_1_rename
    process(R_addr_61_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr_61_resized;
      ov(13 downto 0) := iv;
      R_addr_61_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_62_index_1_resize
    process(addr_buffer) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := addr_buffer;
      ov := iv(13 downto 0);
      R_addr_61_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_62_root_address_inst
    process(array_obj_ref_62_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_62_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_62_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_66_addr_0
    process(ptr_deref_66_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_66_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_66_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_66_base_resize
    process(ptr_64) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_64;
      ov := iv(13 downto 0);
      ptr_deref_66_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_66_gather_scatter
    process(ninput_word_48) --
      variable iv : std_logic_vector(255 downto 0);
      variable ov : std_logic_vector(255 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ninput_word_48;
      ov(255 downto 0) := iv;
      ptr_deref_66_data_0 <= ov(255 downto 0);
      --
    end process;
    -- equivalence ptr_deref_66_root_address_inst
    process(ptr_deref_66_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_66_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_66_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_49_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= ULT_u4_u1_52_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_49_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_49_branch_req_0,
          ack0 => if_stmt_49_branch_ack_0,
          ack1 => if_stmt_49_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u4_u4_32_inst
    process(mycount_17) -- 
      variable tmp_var : std_logic_vector(3 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mycount_17, konst_31_wire_constant, tmp_var);
      nmycount_33 <= tmp_var; --
    end process;
    -- shared split operator group (1) : CONCAT_u240_u256_47_inst 
    ApConcat_group_1: Block -- 
      signal data_in: std_logic_vector(255 downto 0);
      signal data_out: std_logic_vector(255 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= slice_45_wire & val_41;
      ninput_word_48 <= data_out(255 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u240_u256_47_inst_req_0;
      CONCAT_u240_u256_47_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u240_u256_47_inst_req_1;
      CONCAT_u240_u256_47_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_1_gI: SplitGuardInterface generic map(name => "ApConcat_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_1",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 240,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 256,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : CONCAT_u8_u16_40_inst 
    ApConcat_group_2: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= val1_36 & RPIPE_maxpool_input_pipe_39_wire;
      val_41 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u8_u16_40_inst_req_0;
      CONCAT_u8_u16_40_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u8_u16_40_inst_req_1;
      CONCAT_u8_u16_40_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_2_gI: SplitGuardInterface generic map(name => "ApConcat_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_2",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 8, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- binary operator ULT_u4_u1_52_inst
    process(mycount_17) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(mycount_17, konst_51_wire_constant, tmp_var);
      ULT_u4_u1_52_wire <= tmp_var; --
    end process;
    -- shared split operator group (4) : array_obj_ref_62_index_offset 
    ApIntAdd_group_4: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_addr_61_scaled;
      array_obj_ref_62_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_62_index_offset_req_0;
      array_obj_ref_62_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_62_index_offset_req_1;
      array_obj_ref_62_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_4_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_4",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- shared store operator group (0) : ptr_deref_66_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(255 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_66_store_0_req_0;
      ptr_deref_66_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_66_store_0_req_1;
      ptr_deref_66_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_66_word_address_0;
      data_in <= ptr_deref_66_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 256,
        num_reqs => 1,
        tag_length => 3,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(13 downto 0),
          mdata => memory_space_1_sr_data(255 downto 0),
          mtag => memory_space_1_sr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_maxpool_input_pipe_35_inst RPIPE_maxpool_input_pipe_39_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 1 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= RPIPE_maxpool_input_pipe_35_inst_req_0;
      reqL_unguarded(0) <= RPIPE_maxpool_input_pipe_39_inst_req_0;
      RPIPE_maxpool_input_pipe_35_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_maxpool_input_pipe_39_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= RPIPE_maxpool_input_pipe_35_inst_req_1;
      reqR_unguarded(0) <= RPIPE_maxpool_input_pipe_39_inst_req_1;
      RPIPE_maxpool_input_pipe_35_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_maxpool_input_pipe_39_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      val1_36 <= data_out(15 downto 8);
      RPIPE_maxpool_input_pipe_39_wire <= data_out(7 downto 0);
      maxpool_input_pipe_read_0_gI: SplitGuardInterface generic map(name => "maxpool_input_pipe_read_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      maxpool_input_pipe_read_0: InputPortRevised -- 
        generic map ( name => "maxpool_input_pipe_read_0", data_width => 8,  num_reqs => 2,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => maxpool_input_pipe_pipe_read_req(0),
          oack => maxpool_input_pipe_pipe_read_ack(0),
          odata => maxpool_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- 
  end Block; -- data_path
  -- 
end fill_T_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity maxPool3D is -- 
  generic (tag_length : integer); 
  port ( -- 
    maxpool_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    elapsed_time_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_write_data : out  std_logic_vector(63 downto 0);
    maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    fill_T_call_reqs : out  std_logic_vector(0 downto 0);
    fill_T_call_acks : in   std_logic_vector(0 downto 0);
    fill_T_call_data : out  std_logic_vector(63 downto 0);
    fill_T_call_tag  :  out  std_logic_vector(0 downto 0);
    fill_T_return_reqs : out  std_logic_vector(0 downto 0);
    fill_T_return_acks : in   std_logic_vector(0 downto 0);
    fill_T_return_tag :  in   std_logic_vector(0 downto 0);
    timer_call_reqs : out  std_logic_vector(0 downto 0);
    timer_call_acks : in   std_logic_vector(0 downto 0);
    timer_call_tag  :  out  std_logic_vector(1 downto 0);
    timer_return_reqs : out  std_logic_vector(0 downto 0);
    timer_return_acks : in   std_logic_vector(0 downto 0);
    timer_return_data : in   std_logic_vector(63 downto 0);
    timer_return_tag :  in   std_logic_vector(1 downto 0);
    maxPool4_call_reqs : out  std_logic_vector(0 downto 0);
    maxPool4_call_acks : in   std_logic_vector(0 downto 0);
    maxPool4_call_data : out  std_logic_vector(159 downto 0);
    maxPool4_call_tag  :  out  std_logic_vector(0 downto 0);
    maxPool4_return_reqs : out  std_logic_vector(0 downto 0);
    maxPool4_return_acks : in   std_logic_vector(0 downto 0);
    maxPool4_return_data : in   std_logic_vector(7 downto 0);
    maxPool4_return_tag :  in   std_logic_vector(0 downto 0);
    sendB_call_reqs : out  std_logic_vector(0 downto 0);
    sendB_call_acks : in   std_logic_vector(0 downto 0);
    sendB_call_data : out  std_logic_vector(31 downto 0);
    sendB_call_tag  :  out  std_logic_vector(0 downto 0);
    sendB_return_reqs : out  std_logic_vector(0 downto 0);
    sendB_return_acks : in   std_logic_vector(0 downto 0);
    sendB_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity maxPool3D;
architecture maxPool3D_arch of maxPool3D is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal maxPool3D_CP_2658_start: Boolean;
  signal maxPool3D_CP_2658_symbol: Boolean;
  -- volatile/operator module components. 
  component fill_T is -- 
    generic (tag_length : integer); 
    port ( -- 
      addr : in  std_logic_vector(63 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(255 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(2 downto 0);
      maxpool_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      maxpool_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      maxpool_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      c : out  std_logic_vector(63 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component maxPool4 is -- 
    generic (tag_length : integer); 
    port ( -- 
      addr : in  std_logic_vector(31 downto 0);
      addr1 : in  std_logic_vector(31 downto 0);
      addr2 : in  std_logic_vector(31 downto 0);
      addr3 : in  std_logic_vector(31 downto 0);
      addr4 : in  std_logic_vector(31 downto 0);
      output : out  std_logic_vector(7 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(255 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component sendB is -- 
    generic (tag_length : integer); 
    port ( -- 
      size : in  std_logic_vector(31 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
      maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal RPIPE_maxpool_input_pipe_1350_inst_ack_0 : boolean;
  signal type_cast_1354_inst_ack_1 : boolean;
  signal type_cast_1379_inst_ack_0 : boolean;
  signal type_cast_1341_inst_ack_1 : boolean;
  signal call_stmt_1745_call_ack_1 : boolean;
  signal type_cast_1404_inst_req_0 : boolean;
  signal type_cast_1404_inst_ack_0 : boolean;
  signal phi_stmt_1650_ack_0 : boolean;
  signal type_cast_1391_inst_req_1 : boolean;
  signal type_cast_1391_inst_ack_1 : boolean;
  signal call_stmt_1745_call_ack_0 : boolean;
  signal type_cast_1404_inst_req_1 : boolean;
  signal type_cast_1404_inst_ack_1 : boolean;
  signal type_cast_1391_inst_req_0 : boolean;
  signal type_cast_1366_inst_ack_1 : boolean;
  signal type_cast_1391_inst_ack_0 : boolean;
  signal do_while_stmt_1648_branch_req_0 : boolean;
  signal call_stmt_1745_call_req_0 : boolean;
  signal W_rowx_x1_1772_delayed_2_0_1785_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1375_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1375_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1350_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1387_inst_req_1 : boolean;
  signal type_cast_1668_inst_req_0 : boolean;
  signal type_cast_1653_inst_ack_1 : boolean;
  signal type_cast_1366_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1350_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1350_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1400_inst_ack_1 : boolean;
  signal type_cast_1653_inst_req_1 : boolean;
  signal type_cast_1341_inst_req_1 : boolean;
  signal type_cast_1354_inst_req_1 : boolean;
  signal type_cast_1366_inst_ack_0 : boolean;
  signal type_cast_1668_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1362_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1362_inst_req_1 : boolean;
  signal type_cast_1354_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1337_inst_ack_1 : boolean;
  signal call_stmt_1745_call_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1400_inst_ack_0 : boolean;
  signal type_cast_1366_inst_req_0 : boolean;
  signal type_cast_1658_inst_ack_0 : boolean;
  signal type_cast_1341_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1337_inst_req_1 : boolean;
  signal type_cast_1668_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1387_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1400_inst_req_0 : boolean;
  signal type_cast_1658_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1375_inst_ack_1 : boolean;
  signal type_cast_1379_inst_ack_1 : boolean;
  signal type_cast_1341_inst_req_0 : boolean;
  signal type_cast_1354_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1337_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1337_inst_req_0 : boolean;
  signal call_stmt_1824_call_req_0 : boolean;
  signal type_cast_1379_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1362_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1375_inst_req_1 : boolean;
  signal type_cast_1379_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1400_inst_req_1 : boolean;
  signal type_cast_1668_inst_ack_0 : boolean;
  signal type_cast_1783_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1387_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1362_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1387_inst_req_0 : boolean;
  signal W_rowx_x1_1772_delayed_2_0_1785_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1412_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1412_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1412_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1412_inst_ack_1 : boolean;
  signal type_cast_1416_inst_req_0 : boolean;
  signal type_cast_1416_inst_ack_0 : boolean;
  signal type_cast_1416_inst_req_1 : boolean;
  signal type_cast_1416_inst_ack_1 : boolean;
  signal W_colx_x1_1751_delayed_1_0_1761_inst_ack_1 : boolean;
  signal W_colx_x1_1751_delayed_1_0_1761_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1425_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1425_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1425_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1425_inst_ack_1 : boolean;
  signal type_cast_1837_inst_ack_0 : boolean;
  signal type_cast_1828_inst_ack_0 : boolean;
  signal type_cast_1676_inst_ack_1 : boolean;
  signal phi_stmt_1655_ack_0 : boolean;
  signal type_cast_1676_inst_req_1 : boolean;
  signal type_cast_1429_inst_req_0 : boolean;
  signal type_cast_1429_inst_ack_0 : boolean;
  signal type_cast_1429_inst_req_1 : boolean;
  signal type_cast_1429_inst_ack_1 : boolean;
  signal W_colx_x1_1751_delayed_1_0_1761_inst_ack_0 : boolean;
  signal W_colx_x1_1751_delayed_1_0_1761_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1437_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1437_inst_ack_0 : boolean;
  signal type_cast_1653_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1437_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1437_inst_ack_1 : boolean;
  signal type_cast_1837_inst_req_0 : boolean;
  signal type_cast_1828_inst_req_0 : boolean;
  signal if_stmt_1811_branch_ack_0 : boolean;
  signal type_cast_1676_inst_ack_0 : boolean;
  signal phi_stmt_1655_req_1 : boolean;
  signal type_cast_1441_inst_req_0 : boolean;
  signal type_cast_1441_inst_ack_0 : boolean;
  signal type_cast_1441_inst_req_1 : boolean;
  signal type_cast_1663_inst_ack_1 : boolean;
  signal type_cast_1441_inst_ack_1 : boolean;
  signal type_cast_1676_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1450_inst_req_0 : boolean;
  signal type_cast_1663_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1450_inst_ack_0 : boolean;
  signal type_cast_1653_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1450_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1450_inst_ack_1 : boolean;
  signal phi_stmt_1655_req_0 : boolean;
  signal if_stmt_1811_branch_ack_1 : boolean;
  signal type_cast_1454_inst_req_0 : boolean;
  signal type_cast_1454_inst_ack_0 : boolean;
  signal type_cast_1454_inst_req_1 : boolean;
  signal type_cast_1663_inst_ack_0 : boolean;
  signal type_cast_1454_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1462_inst_req_0 : boolean;
  signal type_cast_1663_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1462_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1462_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1462_inst_ack_1 : boolean;
  signal type_cast_1466_inst_req_0 : boolean;
  signal type_cast_1466_inst_ack_0 : boolean;
  signal type_cast_1466_inst_req_1 : boolean;
  signal type_cast_1466_inst_ack_1 : boolean;
  signal type_cast_1759_inst_ack_1 : boolean;
  signal call_stmt_1824_call_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1475_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1475_inst_ack_0 : boolean;
  signal call_stmt_1824_call_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1475_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1475_inst_ack_1 : boolean;
  signal type_cast_1672_inst_ack_1 : boolean;
  signal type_cast_1672_inst_req_1 : boolean;
  signal type_cast_1479_inst_req_0 : boolean;
  signal type_cast_1479_inst_ack_0 : boolean;
  signal type_cast_1479_inst_req_1 : boolean;
  signal type_cast_1479_inst_ack_1 : boolean;
  signal type_cast_1837_inst_ack_1 : boolean;
  signal type_cast_1783_inst_ack_1 : boolean;
  signal type_cast_1783_inst_req_1 : boolean;
  signal type_cast_1489_inst_req_0 : boolean;
  signal type_cast_1489_inst_ack_0 : boolean;
  signal type_cast_1489_inst_req_1 : boolean;
  signal type_cast_1489_inst_ack_1 : boolean;
  signal type_cast_1820_inst_ack_1 : boolean;
  signal type_cast_1837_inst_req_1 : boolean;
  signal type_cast_1820_inst_req_1 : boolean;
  signal type_cast_1759_inst_req_1 : boolean;
  signal if_stmt_1507_branch_req_0 : boolean;
  signal phi_stmt_1650_req_1 : boolean;
  signal if_stmt_1507_branch_ack_1 : boolean;
  signal if_stmt_1507_branch_ack_0 : boolean;
  signal type_cast_1672_inst_ack_0 : boolean;
  signal do_while_stmt_1648_branch_ack_1 : boolean;
  signal type_cast_1544_inst_req_0 : boolean;
  signal type_cast_1544_inst_ack_0 : boolean;
  signal type_cast_1544_inst_req_1 : boolean;
  signal phi_stmt_1660_ack_0 : boolean;
  signal type_cast_1544_inst_ack_1 : boolean;
  signal type_cast_1828_inst_ack_1 : boolean;
  signal type_cast_1672_inst_req_0 : boolean;
  signal call_stmt_1570_call_req_0 : boolean;
  signal call_stmt_1570_call_ack_0 : boolean;
  signal do_while_stmt_1648_branch_ack_0 : boolean;
  signal call_stmt_1570_call_req_1 : boolean;
  signal call_stmt_1570_call_ack_1 : boolean;
  signal type_cast_1828_inst_req_1 : boolean;
  signal phi_stmt_1650_req_0 : boolean;
  signal if_stmt_1582_branch_req_0 : boolean;
  signal if_stmt_1582_branch_ack_1 : boolean;
  signal if_stmt_1582_branch_ack_0 : boolean;
  signal if_stmt_1811_branch_req_0 : boolean;
  signal type_cast_1759_inst_ack_0 : boolean;
  signal call_stmt_1824_call_ack_0 : boolean;
  signal type_cast_1783_inst_ack_0 : boolean;
  signal call_stmt_1605_call_req_0 : boolean;
  signal phi_stmt_1660_req_1 : boolean;
  signal call_stmt_1605_call_ack_0 : boolean;
  signal type_cast_1658_inst_ack_1 : boolean;
  signal W_rowx_x1_1772_delayed_2_0_1785_inst_ack_1 : boolean;
  signal call_stmt_1605_call_req_1 : boolean;
  signal call_stmt_1605_call_ack_1 : boolean;
  signal type_cast_1820_inst_ack_0 : boolean;
  signal type_cast_1820_inst_req_0 : boolean;
  signal W_rowx_x1_1772_delayed_2_0_1785_inst_req_1 : boolean;
  signal type_cast_1609_inst_req_0 : boolean;
  signal type_cast_1609_inst_ack_0 : boolean;
  signal type_cast_1658_inst_req_1 : boolean;
  signal type_cast_1609_inst_req_1 : boolean;
  signal phi_stmt_1660_req_0 : boolean;
  signal type_cast_1609_inst_ack_1 : boolean;
  signal type_cast_1759_inst_req_0 : boolean;
  signal type_cast_1613_inst_req_0 : boolean;
  signal type_cast_1613_inst_ack_0 : boolean;
  signal type_cast_1613_inst_req_1 : boolean;
  signal type_cast_1613_inst_ack_1 : boolean;
  signal type_cast_1617_inst_req_0 : boolean;
  signal type_cast_1617_inst_ack_0 : boolean;
  signal type_cast_1617_inst_req_1 : boolean;
  signal type_cast_1617_inst_ack_1 : boolean;
  signal type_cast_1847_inst_req_0 : boolean;
  signal type_cast_1847_inst_ack_0 : boolean;
  signal type_cast_1847_inst_req_1 : boolean;
  signal type_cast_1847_inst_ack_1 : boolean;
  signal type_cast_1857_inst_req_0 : boolean;
  signal type_cast_1857_inst_ack_0 : boolean;
  signal type_cast_1857_inst_req_1 : boolean;
  signal type_cast_1857_inst_ack_1 : boolean;
  signal type_cast_1867_inst_req_0 : boolean;
  signal type_cast_1867_inst_ack_0 : boolean;
  signal type_cast_1867_inst_req_1 : boolean;
  signal type_cast_1867_inst_ack_1 : boolean;
  signal type_cast_1877_inst_req_0 : boolean;
  signal type_cast_1877_inst_ack_0 : boolean;
  signal type_cast_1877_inst_req_1 : boolean;
  signal type_cast_1877_inst_ack_1 : boolean;
  signal type_cast_1887_inst_req_0 : boolean;
  signal type_cast_1887_inst_ack_0 : boolean;
  signal type_cast_1887_inst_req_1 : boolean;
  signal type_cast_1887_inst_ack_1 : boolean;
  signal type_cast_1897_inst_req_0 : boolean;
  signal type_cast_1897_inst_ack_0 : boolean;
  signal type_cast_1897_inst_req_1 : boolean;
  signal type_cast_1897_inst_ack_1 : boolean;
  signal type_cast_1907_inst_req_0 : boolean;
  signal type_cast_1907_inst_ack_0 : boolean;
  signal type_cast_1907_inst_req_1 : boolean;
  signal type_cast_1907_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1909_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1909_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1909_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1909_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1912_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1912_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1912_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1912_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1915_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1915_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1915_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1915_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1918_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1918_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1918_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1918_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1921_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1921_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1921_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1921_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1924_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1924_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1924_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1924_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1927_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1927_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1927_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1927_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1930_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1930_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1930_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1930_inst_ack_1 : boolean;
  signal WPIPE_elapsed_time_pipe_1933_inst_req_0 : boolean;
  signal WPIPE_elapsed_time_pipe_1933_inst_ack_0 : boolean;
  signal WPIPE_elapsed_time_pipe_1933_inst_req_1 : boolean;
  signal WPIPE_elapsed_time_pipe_1933_inst_ack_1 : boolean;
  signal type_cast_1939_inst_req_0 : boolean;
  signal type_cast_1939_inst_ack_0 : boolean;
  signal type_cast_1939_inst_req_1 : boolean;
  signal type_cast_1939_inst_ack_1 : boolean;
  signal type_cast_1943_inst_req_0 : boolean;
  signal type_cast_1943_inst_ack_0 : boolean;
  signal type_cast_1943_inst_req_1 : boolean;
  signal type_cast_1943_inst_ack_1 : boolean;
  signal call_stmt_1956_call_req_0 : boolean;
  signal call_stmt_1956_call_ack_0 : boolean;
  signal call_stmt_1956_call_req_1 : boolean;
  signal call_stmt_1956_call_ack_1 : boolean;
  signal phi_stmt_1561_req_0 : boolean;
  signal type_cast_1567_inst_req_0 : boolean;
  signal type_cast_1567_inst_ack_0 : boolean;
  signal type_cast_1567_inst_req_1 : boolean;
  signal type_cast_1567_inst_ack_1 : boolean;
  signal phi_stmt_1561_req_1 : boolean;
  signal phi_stmt_1561_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "maxPool3D_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  maxPool3D_CP_2658_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "maxPool3D_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= maxPool3D_CP_2658_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= maxPool3D_CP_2658_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= maxPool3D_CP_2658_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  maxPool3D_CP_2658: Block -- control-path 
    signal maxPool3D_CP_2658_elements: BooleanArray(244 downto 0);
    -- 
  begin -- 
    maxPool3D_CP_2658_elements(0) <= maxPool3D_CP_2658_start;
    maxPool3D_CP_2658_symbol <= maxPool3D_CP_2658_elements(237);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	29 
    -- CP-element group 0: 	33 
    -- CP-element group 0: 	37 
    -- CP-element group 0: 	41 
    -- CP-element group 0: 	45 
    -- CP-element group 0: 	49 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	5 
    -- CP-element group 0: 	9 
    -- CP-element group 0: 	13 
    -- CP-element group 0: 	17 
    -- CP-element group 0: 	21 
    -- CP-element group 0: 	25 
    -- CP-element group 0:  members (44) 
      -- CP-element group 0: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1391_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1366_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485__entry__
      -- CP-element group 0: 	 branch_block_stmt_1335/branch_block_stmt_1335__entry__
      -- CP-element group 0: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1404_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1391_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1404_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1391_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1404_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1366_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1341_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1354_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1341_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1354_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1379_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1337_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1379_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1337_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1354_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1337_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1335/$entry
      -- CP-element group 0: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/$entry
      -- CP-element group 0: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1366_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1379_Update/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1341_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1416_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1416_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1416_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1429_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1429_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1429_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1441_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1441_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1441_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1454_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1454_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1454_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1466_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1466_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1466_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1479_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1479_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1479_Update/cr
      -- 
    cr_2849_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2849_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(0), ack => type_cast_1391_inst_req_1); -- 
    cr_2877_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2877_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(0), ack => type_cast_1404_inst_req_1); -- 
    cr_2793_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2793_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(0), ack => type_cast_1366_inst_req_1); -- 
    cr_2737_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2737_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(0), ack => type_cast_1341_inst_req_1); -- 
    cr_2765_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2765_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(0), ack => type_cast_1354_inst_req_1); -- 
    rr_2718_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2718_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(0), ack => RPIPE_maxpool_input_pipe_1337_inst_req_0); -- 
    cr_2821_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2821_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(0), ack => type_cast_1379_inst_req_1); -- 
    cr_2905_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2905_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(0), ack => type_cast_1416_inst_req_1); -- 
    cr_2933_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2933_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(0), ack => type_cast_1429_inst_req_1); -- 
    cr_2961_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2961_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(0), ack => type_cast_1441_inst_req_1); -- 
    cr_2989_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2989_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(0), ack => type_cast_1454_inst_req_1); -- 
    cr_3017_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3017_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(0), ack => type_cast_1466_inst_req_1); -- 
    cr_3045_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3045_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(0), ack => type_cast_1479_inst_req_1); -- 
    -- CP-element group 1:  branch  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	180 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	181 
    -- CP-element group 1: 	182 
    -- CP-element group 1:  members (9) 
      -- CP-element group 1: 	 branch_block_stmt_1335/do_while_stmt_1648__exit__
      -- CP-element group 1: 	 branch_block_stmt_1335/if_stmt_1811__entry__
      -- CP-element group 1: 	 branch_block_stmt_1335/if_stmt_1811_dead_link/$entry
      -- CP-element group 1: 	 branch_block_stmt_1335/if_stmt_1811_else_link/$entry
      -- CP-element group 1: 	 branch_block_stmt_1335/if_stmt_1811_if_link/$entry
      -- CP-element group 1: 	 branch_block_stmt_1335/R_whilex_xbody_whilex_xend_taken_1812_place
      -- CP-element group 1: 	 branch_block_stmt_1335/if_stmt_1811_eval_test/branch_req
      -- CP-element group 1: 	 branch_block_stmt_1335/if_stmt_1811_eval_test/$exit
      -- CP-element group 1: 	 branch_block_stmt_1335/if_stmt_1811_eval_test/$entry
      -- 
    branch_req_3482_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3482_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(1), ack => if_stmt_1811_branch_req_0); -- 
    maxPool3D_CP_2658_elements(1) <= maxPool3D_CP_2658_elements(180);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1337_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1337_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1337_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1337_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1337_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1337_sample_completed_
      -- 
    ra_2719_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1337_inst_ack_0, ack => maxPool3D_CP_2658_elements(2)); -- 
    cr_2723_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2723_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(2), ack => RPIPE_maxpool_input_pipe_1337_inst_req_1); -- 
    -- CP-element group 3:  fork  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3: 	6 
    -- CP-element group 3:  members (9) 
      -- CP-element group 3: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1350_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1341_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1350_Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1337_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1337_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1341_Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1341_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1350_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1337_update_completed_
      -- 
    ca_2724_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1337_inst_ack_1, ack => maxPool3D_CP_2658_elements(3)); -- 
    rr_2732_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2732_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(3), ack => type_cast_1341_inst_req_0); -- 
    rr_2746_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2746_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(3), ack => RPIPE_maxpool_input_pipe_1350_inst_req_0); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1341_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1341_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1341_Sample/$exit
      -- 
    ra_2733_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1341_inst_ack_0, ack => maxPool3D_CP_2658_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	50 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1341_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1341_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1341_update_completed_
      -- 
    ca_2738_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1341_inst_ack_1, ack => maxPool3D_CP_2658_elements(5)); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	3 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1350_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1350_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1350_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1350_Update/cr
      -- CP-element group 6: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1350_update_start_
      -- CP-element group 6: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1350_sample_completed_
      -- 
    ra_2747_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1350_inst_ack_0, ack => maxPool3D_CP_2658_elements(6)); -- 
    cr_2751_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2751_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(6), ack => RPIPE_maxpool_input_pipe_1350_inst_req_1); -- 
    -- CP-element group 7:  fork  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7: 	10 
    -- CP-element group 7:  members (9) 
      -- CP-element group 7: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1350_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1350_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1350_Update/ca
      -- CP-element group 7: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1354_Sample/rr
      -- CP-element group 7: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1354_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1362_Sample/rr
      -- CP-element group 7: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1362_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1354_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1362_sample_start_
      -- 
    ca_2752_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1350_inst_ack_1, ack => maxPool3D_CP_2658_elements(7)); -- 
    rr_2760_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2760_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(7), ack => type_cast_1354_inst_req_0); -- 
    rr_2774_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2774_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(7), ack => RPIPE_maxpool_input_pipe_1362_inst_req_0); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1354_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1354_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1354_sample_completed_
      -- 
    ra_2761_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1354_inst_ack_0, ack => maxPool3D_CP_2658_elements(8)); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	0 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	50 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1354_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1354_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1354_update_completed_
      -- 
    ca_2766_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1354_inst_ack_1, ack => maxPool3D_CP_2658_elements(9)); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	7 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (6) 
      -- CP-element group 10: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1362_Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1362_Update/cr
      -- CP-element group 10: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1362_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1362_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1362_update_start_
      -- CP-element group 10: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1362_sample_completed_
      -- 
    ra_2775_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1362_inst_ack_0, ack => maxPool3D_CP_2658_elements(10)); -- 
    cr_2779_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2779_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(10), ack => RPIPE_maxpool_input_pipe_1362_inst_req_1); -- 
    -- CP-element group 11:  fork  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11: 	14 
    -- CP-element group 11:  members (9) 
      -- CP-element group 11: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1375_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1366_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1362_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1362_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1366_Sample/rr
      -- CP-element group 11: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1375_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1366_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1375_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1362_update_completed_
      -- 
    ca_2780_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1362_inst_ack_1, ack => maxPool3D_CP_2658_elements(11)); -- 
    rr_2788_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2788_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(11), ack => type_cast_1366_inst_req_0); -- 
    rr_2802_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2802_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(11), ack => RPIPE_maxpool_input_pipe_1375_inst_req_0); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1366_Sample/ra
      -- CP-element group 12: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1366_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1366_sample_completed_
      -- 
    ra_2789_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1366_inst_ack_0, ack => maxPool3D_CP_2658_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	0 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	50 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1366_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1366_Update/ca
      -- CP-element group 13: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1366_update_completed_
      -- 
    ca_2794_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1366_inst_ack_1, ack => maxPool3D_CP_2658_elements(13)); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	11 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (6) 
      -- CP-element group 14: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1375_Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1375_Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1375_Update/cr
      -- CP-element group 14: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1375_update_start_
      -- CP-element group 14: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1375_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1375_Update/$entry
      -- 
    ra_2803_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1375_inst_ack_0, ack => maxPool3D_CP_2658_elements(14)); -- 
    cr_2807_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2807_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(14), ack => RPIPE_maxpool_input_pipe_1375_inst_req_1); -- 
    -- CP-element group 15:  fork  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15: 	18 
    -- CP-element group 15:  members (9) 
      -- CP-element group 15: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1379_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1387_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1387_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1375_Update/ca
      -- CP-element group 15: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1375_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1379_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1375_Update/$exit
      -- CP-element group 15: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1379_Sample/rr
      -- CP-element group 15: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1387_Sample/rr
      -- 
    ca_2808_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1375_inst_ack_1, ack => maxPool3D_CP_2658_elements(15)); -- 
    rr_2816_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2816_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(15), ack => type_cast_1379_inst_req_0); -- 
    rr_2830_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2830_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(15), ack => RPIPE_maxpool_input_pipe_1387_inst_req_0); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1379_Sample/ra
      -- CP-element group 16: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1379_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1379_Sample/$exit
      -- 
    ra_2817_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1379_inst_ack_0, ack => maxPool3D_CP_2658_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	0 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	50 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1379_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1379_Update/ca
      -- CP-element group 17: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1379_Update/$exit
      -- 
    ca_2822_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1379_inst_ack_1, ack => maxPool3D_CP_2658_elements(17)); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	15 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1387_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1387_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1387_update_start_
      -- CP-element group 18: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1387_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1387_Update/cr
      -- CP-element group 18: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1387_Sample/ra
      -- 
    ra_2831_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1387_inst_ack_0, ack => maxPool3D_CP_2658_elements(18)); -- 
    cr_2835_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2835_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(18), ack => RPIPE_maxpool_input_pipe_1387_inst_req_1); -- 
    -- CP-element group 19:  fork  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19: 	22 
    -- CP-element group 19:  members (9) 
      -- CP-element group 19: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1387_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1391_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1400_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1387_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1391_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1400_Sample/rr
      -- CP-element group 19: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1400_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1387_Update/ca
      -- CP-element group 19: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1391_sample_start_
      -- 
    ca_2836_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1387_inst_ack_1, ack => maxPool3D_CP_2658_elements(19)); -- 
    rr_2844_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2844_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(19), ack => type_cast_1391_inst_req_0); -- 
    rr_2858_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2858_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(19), ack => RPIPE_maxpool_input_pipe_1400_inst_req_0); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1391_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1391_Sample/ra
      -- CP-element group 20: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1391_sample_completed_
      -- 
    ra_2845_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1391_inst_ack_0, ack => maxPool3D_CP_2658_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	0 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	50 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1391_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1391_Update/ca
      -- CP-element group 21: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1391_Update/$exit
      -- 
    ca_2850_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1391_inst_ack_1, ack => maxPool3D_CP_2658_elements(21)); -- 
    -- CP-element group 22:  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	19 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (6) 
      -- CP-element group 22: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1400_update_start_
      -- CP-element group 22: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1400_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1400_Sample/ra
      -- CP-element group 22: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1400_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1400_Update/$entry
      -- CP-element group 22: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1400_Update/cr
      -- 
    ra_2859_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1400_inst_ack_0, ack => maxPool3D_CP_2658_elements(22)); -- 
    cr_2863_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2863_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(22), ack => RPIPE_maxpool_input_pipe_1400_inst_req_1); -- 
    -- CP-element group 23:  fork  transition  input  output  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	26 
    -- CP-element group 23: 	24 
    -- CP-element group 23:  members (9) 
      -- CP-element group 23: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1404_Sample/rr
      -- CP-element group 23: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1404_sample_start_
      -- CP-element group 23: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1400_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1404_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1400_Update/ca
      -- CP-element group 23: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1400_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1412_sample_start_
      -- CP-element group 23: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1412_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1412_Sample/rr
      -- 
    ca_2864_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1400_inst_ack_1, ack => maxPool3D_CP_2658_elements(23)); -- 
    rr_2872_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2872_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(23), ack => type_cast_1404_inst_req_0); -- 
    rr_2886_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2886_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(23), ack => RPIPE_maxpool_input_pipe_1412_inst_req_0); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1404_Sample/ra
      -- CP-element group 24: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1404_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1404_sample_completed_
      -- 
    ra_2873_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1404_inst_ack_0, ack => maxPool3D_CP_2658_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	0 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	50 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1404_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1404_Update/ca
      -- CP-element group 25: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1404_update_completed_
      -- 
    ca_2878_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1404_inst_ack_1, ack => maxPool3D_CP_2658_elements(25)); -- 
    -- CP-element group 26:  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	23 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (6) 
      -- CP-element group 26: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1412_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1412_update_start_
      -- CP-element group 26: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1412_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1412_Sample/ra
      -- CP-element group 26: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1412_Update/$entry
      -- CP-element group 26: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1412_Update/cr
      -- 
    ra_2887_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1412_inst_ack_0, ack => maxPool3D_CP_2658_elements(26)); -- 
    cr_2891_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2891_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(26), ack => RPIPE_maxpool_input_pipe_1412_inst_req_1); -- 
    -- CP-element group 27:  fork  transition  input  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27: 	30 
    -- CP-element group 27:  members (9) 
      -- CP-element group 27: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1412_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1412_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1412_Update/ca
      -- CP-element group 27: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1416_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1416_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1416_Sample/rr
      -- CP-element group 27: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1425_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1425_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1425_Sample/rr
      -- 
    ca_2892_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1412_inst_ack_1, ack => maxPool3D_CP_2658_elements(27)); -- 
    rr_2900_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2900_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(27), ack => type_cast_1416_inst_req_0); -- 
    rr_2914_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2914_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(27), ack => RPIPE_maxpool_input_pipe_1425_inst_req_0); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1416_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1416_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1416_Sample/ra
      -- 
    ra_2901_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1416_inst_ack_0, ack => maxPool3D_CP_2658_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	0 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	50 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1416_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1416_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1416_Update/ca
      -- 
    ca_2906_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1416_inst_ack_1, ack => maxPool3D_CP_2658_elements(29)); -- 
    -- CP-element group 30:  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	27 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (6) 
      -- CP-element group 30: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1425_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1425_update_start_
      -- CP-element group 30: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1425_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1425_Sample/ra
      -- CP-element group 30: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1425_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1425_Update/cr
      -- 
    ra_2915_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1425_inst_ack_0, ack => maxPool3D_CP_2658_elements(30)); -- 
    cr_2919_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2919_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(30), ack => RPIPE_maxpool_input_pipe_1425_inst_req_1); -- 
    -- CP-element group 31:  fork  transition  input  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31: 	34 
    -- CP-element group 31:  members (9) 
      -- CP-element group 31: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1425_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1425_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1425_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1429_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1429_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1429_Sample/rr
      -- CP-element group 31: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1437_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1437_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1437_Sample/rr
      -- 
    ca_2920_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1425_inst_ack_1, ack => maxPool3D_CP_2658_elements(31)); -- 
    rr_2928_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2928_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(31), ack => type_cast_1429_inst_req_0); -- 
    rr_2942_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2942_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(31), ack => RPIPE_maxpool_input_pipe_1437_inst_req_0); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1429_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1429_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1429_Sample/ra
      -- 
    ra_2929_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1429_inst_ack_0, ack => maxPool3D_CP_2658_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	0 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	50 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1429_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1429_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1429_Update/ca
      -- 
    ca_2934_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1429_inst_ack_1, ack => maxPool3D_CP_2658_elements(33)); -- 
    -- CP-element group 34:  transition  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	31 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34:  members (6) 
      -- CP-element group 34: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1437_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1437_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1437_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1437_Sample/ra
      -- CP-element group 34: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1437_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1437_Update/cr
      -- 
    ra_2943_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1437_inst_ack_0, ack => maxPool3D_CP_2658_elements(34)); -- 
    cr_2947_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2947_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(34), ack => RPIPE_maxpool_input_pipe_1437_inst_req_1); -- 
    -- CP-element group 35:  fork  transition  input  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35: 	38 
    -- CP-element group 35:  members (9) 
      -- CP-element group 35: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1437_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1437_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1437_Update/ca
      -- CP-element group 35: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1441_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1441_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1441_Sample/rr
      -- CP-element group 35: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1450_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1450_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1450_Sample/rr
      -- 
    ca_2948_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1437_inst_ack_1, ack => maxPool3D_CP_2658_elements(35)); -- 
    rr_2956_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2956_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(35), ack => type_cast_1441_inst_req_0); -- 
    rr_2970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(35), ack => RPIPE_maxpool_input_pipe_1450_inst_req_0); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1441_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1441_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1441_Sample/ra
      -- 
    ra_2957_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1441_inst_ack_0, ack => maxPool3D_CP_2658_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	0 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	50 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1441_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1441_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1441_Update/ca
      -- 
    ca_2962_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1441_inst_ack_1, ack => maxPool3D_CP_2658_elements(37)); -- 
    -- CP-element group 38:  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	35 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (6) 
      -- CP-element group 38: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1450_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1450_update_start_
      -- CP-element group 38: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1450_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1450_Sample/ra
      -- CP-element group 38: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1450_Update/$entry
      -- CP-element group 38: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1450_Update/cr
      -- 
    ra_2971_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1450_inst_ack_0, ack => maxPool3D_CP_2658_elements(38)); -- 
    cr_2975_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2975_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(38), ack => RPIPE_maxpool_input_pipe_1450_inst_req_1); -- 
    -- CP-element group 39:  fork  transition  input  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39: 	42 
    -- CP-element group 39:  members (9) 
      -- CP-element group 39: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1450_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1450_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1450_Update/ca
      -- CP-element group 39: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1454_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1454_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1454_Sample/rr
      -- CP-element group 39: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1462_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1462_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1462_Sample/rr
      -- 
    ca_2976_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1450_inst_ack_1, ack => maxPool3D_CP_2658_elements(39)); -- 
    rr_2984_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2984_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(39), ack => type_cast_1454_inst_req_0); -- 
    rr_2998_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2998_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(39), ack => RPIPE_maxpool_input_pipe_1462_inst_req_0); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1454_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1454_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1454_Sample/ra
      -- 
    ra_2985_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1454_inst_ack_0, ack => maxPool3D_CP_2658_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	0 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	50 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1454_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1454_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1454_Update/ca
      -- 
    ca_2990_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1454_inst_ack_1, ack => maxPool3D_CP_2658_elements(41)); -- 
    -- CP-element group 42:  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	39 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (6) 
      -- CP-element group 42: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1462_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1462_update_start_
      -- CP-element group 42: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1462_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1462_Sample/ra
      -- CP-element group 42: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1462_Update/$entry
      -- CP-element group 42: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1462_Update/cr
      -- 
    ra_2999_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1462_inst_ack_0, ack => maxPool3D_CP_2658_elements(42)); -- 
    cr_3003_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3003_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(42), ack => RPIPE_maxpool_input_pipe_1462_inst_req_1); -- 
    -- CP-element group 43:  fork  transition  input  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43: 	46 
    -- CP-element group 43:  members (9) 
      -- CP-element group 43: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1462_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1462_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1462_Update/ca
      -- CP-element group 43: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1466_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1466_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1466_Sample/rr
      -- CP-element group 43: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1475_sample_start_
      -- CP-element group 43: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1475_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1475_Sample/rr
      -- 
    ca_3004_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1462_inst_ack_1, ack => maxPool3D_CP_2658_elements(43)); -- 
    rr_3012_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3012_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(43), ack => type_cast_1466_inst_req_0); -- 
    rr_3026_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3026_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(43), ack => RPIPE_maxpool_input_pipe_1475_inst_req_0); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1466_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1466_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1466_Sample/ra
      -- 
    ra_3013_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1466_inst_ack_0, ack => maxPool3D_CP_2658_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	0 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	50 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1466_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1466_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1466_Update/ca
      -- 
    ca_3018_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1466_inst_ack_1, ack => maxPool3D_CP_2658_elements(45)); -- 
    -- CP-element group 46:  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	43 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (6) 
      -- CP-element group 46: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1475_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1475_update_start_
      -- CP-element group 46: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1475_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1475_Sample/ra
      -- CP-element group 46: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1475_Update/$entry
      -- CP-element group 46: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1475_Update/cr
      -- 
    ra_3027_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1475_inst_ack_0, ack => maxPool3D_CP_2658_elements(46)); -- 
    cr_3031_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3031_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(46), ack => RPIPE_maxpool_input_pipe_1475_inst_req_1); -- 
    -- CP-element group 47:  transition  input  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (6) 
      -- CP-element group 47: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1475_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1475_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/RPIPE_maxpool_input_pipe_1475_Update/ca
      -- CP-element group 47: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1479_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1479_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1479_Sample/rr
      -- 
    ca_3032_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1475_inst_ack_1, ack => maxPool3D_CP_2658_elements(47)); -- 
    rr_3040_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3040_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(47), ack => type_cast_1479_inst_req_0); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1479_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1479_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1479_Sample/ra
      -- 
    ra_3041_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1479_inst_ack_0, ack => maxPool3D_CP_2658_elements(48)); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	0 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1479_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1479_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/type_cast_1479_Update/ca
      -- 
    ca_3046_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1479_inst_ack_1, ack => maxPool3D_CP_2658_elements(49)); -- 
    -- CP-element group 50:  join  fork  transition  place  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	29 
    -- CP-element group 50: 	33 
    -- CP-element group 50: 	37 
    -- CP-element group 50: 	41 
    -- CP-element group 50: 	45 
    -- CP-element group 50: 	49 
    -- CP-element group 50: 	5 
    -- CP-element group 50: 	9 
    -- CP-element group 50: 	13 
    -- CP-element group 50: 	17 
    -- CP-element group 50: 	21 
    -- CP-element group 50: 	25 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (10) 
      -- CP-element group 50: 	 branch_block_stmt_1335/assign_stmt_1490_to_assign_stmt_1506__entry__
      -- CP-element group 50: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485__exit__
      -- CP-element group 50: 	 branch_block_stmt_1335/assign_stmt_1338_to_assign_stmt_1485/$exit
      -- CP-element group 50: 	 branch_block_stmt_1335/assign_stmt_1490_to_assign_stmt_1506/$entry
      -- CP-element group 50: 	 branch_block_stmt_1335/assign_stmt_1490_to_assign_stmt_1506/type_cast_1489_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_1335/assign_stmt_1490_to_assign_stmt_1506/type_cast_1489_update_start_
      -- CP-element group 50: 	 branch_block_stmt_1335/assign_stmt_1490_to_assign_stmt_1506/type_cast_1489_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_1335/assign_stmt_1490_to_assign_stmt_1506/type_cast_1489_Sample/rr
      -- CP-element group 50: 	 branch_block_stmt_1335/assign_stmt_1490_to_assign_stmt_1506/type_cast_1489_Update/$entry
      -- CP-element group 50: 	 branch_block_stmt_1335/assign_stmt_1490_to_assign_stmt_1506/type_cast_1489_Update/cr
      -- 
    rr_3057_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3057_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(50), ack => type_cast_1489_inst_req_0); -- 
    cr_3062_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3062_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(50), ack => type_cast_1489_inst_req_1); -- 
    maxPool3D_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 11) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1);
      constant place_markings: IntegerArray(0 to 11)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0);
      constant place_delays: IntegerArray(0 to 11) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0);
      constant joinName: string(1 to 29) := "maxPool3D_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 12); -- 
    begin -- 
      preds <= maxPool3D_CP_2658_elements(29) & maxPool3D_CP_2658_elements(33) & maxPool3D_CP_2658_elements(37) & maxPool3D_CP_2658_elements(41) & maxPool3D_CP_2658_elements(45) & maxPool3D_CP_2658_elements(49) & maxPool3D_CP_2658_elements(5) & maxPool3D_CP_2658_elements(9) & maxPool3D_CP_2658_elements(13) & maxPool3D_CP_2658_elements(17) & maxPool3D_CP_2658_elements(21) & maxPool3D_CP_2658_elements(25);
      gj_maxPool3D_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 12, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2658_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_1335/assign_stmt_1490_to_assign_stmt_1506/type_cast_1489_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_1335/assign_stmt_1490_to_assign_stmt_1506/type_cast_1489_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_1335/assign_stmt_1490_to_assign_stmt_1506/type_cast_1489_Sample/ra
      -- 
    ra_3058_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1489_inst_ack_0, ack => maxPool3D_CP_2658_elements(51)); -- 
    -- CP-element group 52:  branch  transition  place  input  output  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	53 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (13) 
      -- CP-element group 52: 	 branch_block_stmt_1335/assign_stmt_1490_to_assign_stmt_1506__exit__
      -- CP-element group 52: 	 branch_block_stmt_1335/if_stmt_1507__entry__
      -- CP-element group 52: 	 branch_block_stmt_1335/assign_stmt_1490_to_assign_stmt_1506/$exit
      -- CP-element group 52: 	 branch_block_stmt_1335/assign_stmt_1490_to_assign_stmt_1506/type_cast_1489_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_1335/assign_stmt_1490_to_assign_stmt_1506/type_cast_1489_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_1335/assign_stmt_1490_to_assign_stmt_1506/type_cast_1489_Update/ca
      -- CP-element group 52: 	 branch_block_stmt_1335/if_stmt_1507_dead_link/$entry
      -- CP-element group 52: 	 branch_block_stmt_1335/if_stmt_1507_eval_test/$entry
      -- CP-element group 52: 	 branch_block_stmt_1335/if_stmt_1507_eval_test/$exit
      -- CP-element group 52: 	 branch_block_stmt_1335/if_stmt_1507_eval_test/branch_req
      -- CP-element group 52: 	 branch_block_stmt_1335/R_cmp257_1508_place
      -- CP-element group 52: 	 branch_block_stmt_1335/if_stmt_1507_if_link/$entry
      -- CP-element group 52: 	 branch_block_stmt_1335/if_stmt_1507_else_link/$entry
      -- 
    ca_3063_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1489_inst_ack_1, ack => maxPool3D_CP_2658_elements(52)); -- 
    branch_req_3071_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3071_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(52), ack => if_stmt_1507_branch_req_0); -- 
    -- CP-element group 53:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	52 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53: 	56 
    -- CP-element group 53:  members (18) 
      -- CP-element group 53: 	 branch_block_stmt_1335/assign_stmt_1518_to_assign_stmt_1558__entry__
      -- CP-element group 53: 	 branch_block_stmt_1335/merge_stmt_1513__exit__
      -- CP-element group 53: 	 branch_block_stmt_1335/if_stmt_1507_if_link/$exit
      -- CP-element group 53: 	 branch_block_stmt_1335/if_stmt_1507_if_link/if_choice_transition
      -- CP-element group 53: 	 branch_block_stmt_1335/entry_bbx_xnph
      -- CP-element group 53: 	 branch_block_stmt_1335/assign_stmt_1518_to_assign_stmt_1558/$entry
      -- CP-element group 53: 	 branch_block_stmt_1335/assign_stmt_1518_to_assign_stmt_1558/type_cast_1544_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_1335/assign_stmt_1518_to_assign_stmt_1558/type_cast_1544_update_start_
      -- CP-element group 53: 	 branch_block_stmt_1335/assign_stmt_1518_to_assign_stmt_1558/type_cast_1544_Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_1335/assign_stmt_1518_to_assign_stmt_1558/type_cast_1544_Sample/rr
      -- CP-element group 53: 	 branch_block_stmt_1335/assign_stmt_1518_to_assign_stmt_1558/type_cast_1544_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_1335/assign_stmt_1518_to_assign_stmt_1558/type_cast_1544_Update/cr
      -- CP-element group 53: 	 branch_block_stmt_1335/entry_bbx_xnph_PhiReq/$entry
      -- CP-element group 53: 	 branch_block_stmt_1335/entry_bbx_xnph_PhiReq/$exit
      -- CP-element group 53: 	 branch_block_stmt_1335/merge_stmt_1513_PhiReqMerge
      -- CP-element group 53: 	 branch_block_stmt_1335/merge_stmt_1513_PhiAck/$entry
      -- CP-element group 53: 	 branch_block_stmt_1335/merge_stmt_1513_PhiAck/$exit
      -- CP-element group 53: 	 branch_block_stmt_1335/merge_stmt_1513_PhiAck/dummy
      -- 
    if_choice_transition_3076_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1507_branch_ack_1, ack => maxPool3D_CP_2658_elements(53)); -- 
    rr_3093_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3093_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(53), ack => type_cast_1544_inst_req_0); -- 
    cr_3098_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3098_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(53), ack => type_cast_1544_inst_req_1); -- 
    -- CP-element group 54:  transition  place  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	244 
    -- CP-element group 54:  members (5) 
      -- CP-element group 54: 	 branch_block_stmt_1335/if_stmt_1507_else_link/$exit
      -- CP-element group 54: 	 branch_block_stmt_1335/if_stmt_1507_else_link/else_choice_transition
      -- CP-element group 54: 	 branch_block_stmt_1335/entry_forx_xend
      -- CP-element group 54: 	 branch_block_stmt_1335/entry_forx_xend_PhiReq/$entry
      -- CP-element group 54: 	 branch_block_stmt_1335/entry_forx_xend_PhiReq/$exit
      -- 
    else_choice_transition_3080_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1507_branch_ack_0, ack => maxPool3D_CP_2658_elements(54)); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_1335/assign_stmt_1518_to_assign_stmt_1558/type_cast_1544_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_1335/assign_stmt_1518_to_assign_stmt_1558/type_cast_1544_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_1335/assign_stmt_1518_to_assign_stmt_1558/type_cast_1544_Sample/ra
      -- 
    ra_3094_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1544_inst_ack_0, ack => maxPool3D_CP_2658_elements(55)); -- 
    -- CP-element group 56:  transition  place  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	53 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	238 
    -- CP-element group 56:  members (9) 
      -- CP-element group 56: 	 branch_block_stmt_1335/bbx_xnph_forx_xbody
      -- CP-element group 56: 	 branch_block_stmt_1335/assign_stmt_1518_to_assign_stmt_1558__exit__
      -- CP-element group 56: 	 branch_block_stmt_1335/assign_stmt_1518_to_assign_stmt_1558/$exit
      -- CP-element group 56: 	 branch_block_stmt_1335/assign_stmt_1518_to_assign_stmt_1558/type_cast_1544_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_1335/assign_stmt_1518_to_assign_stmt_1558/type_cast_1544_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_1335/assign_stmt_1518_to_assign_stmt_1558/type_cast_1544_Update/ca
      -- CP-element group 56: 	 branch_block_stmt_1335/bbx_xnph_forx_xbody_PhiReq/$entry
      -- CP-element group 56: 	 branch_block_stmt_1335/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1561/$entry
      -- CP-element group 56: 	 branch_block_stmt_1335/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1561/phi_stmt_1561_sources/$entry
      -- 
    ca_3099_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1544_inst_ack_1, ack => maxPool3D_CP_2658_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	243 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_1335/call_stmt_1570_to_assign_stmt_1581/call_stmt_1570_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_1335/call_stmt_1570_to_assign_stmt_1581/call_stmt_1570_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_1335/call_stmt_1570_to_assign_stmt_1581/call_stmt_1570_Sample/cra
      -- 
    cra_3111_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1570_call_ack_0, ack => maxPool3D_CP_2658_elements(57)); -- 
    -- CP-element group 58:  branch  transition  place  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	243 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58: 	60 
    -- CP-element group 58:  members (13) 
      -- CP-element group 58: 	 branch_block_stmt_1335/call_stmt_1570_to_assign_stmt_1581__exit__
      -- CP-element group 58: 	 branch_block_stmt_1335/if_stmt_1582__entry__
      -- CP-element group 58: 	 branch_block_stmt_1335/call_stmt_1570_to_assign_stmt_1581/$exit
      -- CP-element group 58: 	 branch_block_stmt_1335/call_stmt_1570_to_assign_stmt_1581/call_stmt_1570_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_1335/call_stmt_1570_to_assign_stmt_1581/call_stmt_1570_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_1335/call_stmt_1570_to_assign_stmt_1581/call_stmt_1570_Update/cca
      -- CP-element group 58: 	 branch_block_stmt_1335/if_stmt_1582_dead_link/$entry
      -- CP-element group 58: 	 branch_block_stmt_1335/if_stmt_1582_eval_test/$entry
      -- CP-element group 58: 	 branch_block_stmt_1335/if_stmt_1582_eval_test/$exit
      -- CP-element group 58: 	 branch_block_stmt_1335/if_stmt_1582_eval_test/branch_req
      -- CP-element group 58: 	 branch_block_stmt_1335/R_exitcond1_1583_place
      -- CP-element group 58: 	 branch_block_stmt_1335/if_stmt_1582_if_link/$entry
      -- CP-element group 58: 	 branch_block_stmt_1335/if_stmt_1582_else_link/$entry
      -- 
    cca_3116_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1570_call_ack_1, ack => maxPool3D_CP_2658_elements(58)); -- 
    branch_req_3124_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3124_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(58), ack => if_stmt_1582_branch_req_0); -- 
    -- CP-element group 59:  merge  transition  place  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	244 
    -- CP-element group 59:  members (13) 
      -- CP-element group 59: 	 branch_block_stmt_1335/merge_stmt_1588__exit__
      -- CP-element group 59: 	 branch_block_stmt_1335/forx_xendx_xloopexit_forx_xend
      -- CP-element group 59: 	 branch_block_stmt_1335/if_stmt_1582_if_link/$exit
      -- CP-element group 59: 	 branch_block_stmt_1335/if_stmt_1582_if_link/if_choice_transition
      -- CP-element group 59: 	 branch_block_stmt_1335/forx_xbody_forx_xendx_xloopexit
      -- CP-element group 59: 	 branch_block_stmt_1335/forx_xbody_forx_xendx_xloopexit_PhiReq/$entry
      -- CP-element group 59: 	 branch_block_stmt_1335/forx_xbody_forx_xendx_xloopexit_PhiReq/$exit
      -- CP-element group 59: 	 branch_block_stmt_1335/merge_stmt_1588_PhiReqMerge
      -- CP-element group 59: 	 branch_block_stmt_1335/merge_stmt_1588_PhiAck/$entry
      -- CP-element group 59: 	 branch_block_stmt_1335/merge_stmt_1588_PhiAck/$exit
      -- CP-element group 59: 	 branch_block_stmt_1335/merge_stmt_1588_PhiAck/dummy
      -- CP-element group 59: 	 branch_block_stmt_1335/forx_xendx_xloopexit_forx_xend_PhiReq/$entry
      -- CP-element group 59: 	 branch_block_stmt_1335/forx_xendx_xloopexit_forx_xend_PhiReq/$exit
      -- 
    if_choice_transition_3129_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1582_branch_ack_1, ack => maxPool3D_CP_2658_elements(59)); -- 
    -- CP-element group 60:  fork  transition  place  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	58 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	239 
    -- CP-element group 60: 	240 
    -- CP-element group 60:  members (12) 
      -- CP-element group 60: 	 branch_block_stmt_1335/if_stmt_1582_else_link/$exit
      -- CP-element group 60: 	 branch_block_stmt_1335/if_stmt_1582_else_link/else_choice_transition
      -- CP-element group 60: 	 branch_block_stmt_1335/forx_xbody_forx_xbody
      -- CP-element group 60: 	 branch_block_stmt_1335/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 60: 	 branch_block_stmt_1335/forx_xbody_forx_xbody_PhiReq/phi_stmt_1561/$entry
      -- CP-element group 60: 	 branch_block_stmt_1335/forx_xbody_forx_xbody_PhiReq/phi_stmt_1561/phi_stmt_1561_sources/$entry
      -- CP-element group 60: 	 branch_block_stmt_1335/forx_xbody_forx_xbody_PhiReq/phi_stmt_1561/phi_stmt_1561_sources/type_cast_1567/$entry
      -- CP-element group 60: 	 branch_block_stmt_1335/forx_xbody_forx_xbody_PhiReq/phi_stmt_1561/phi_stmt_1561_sources/type_cast_1567/SplitProtocol/$entry
      -- CP-element group 60: 	 branch_block_stmt_1335/forx_xbody_forx_xbody_PhiReq/phi_stmt_1561/phi_stmt_1561_sources/type_cast_1567/SplitProtocol/Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_1335/forx_xbody_forx_xbody_PhiReq/phi_stmt_1561/phi_stmt_1561_sources/type_cast_1567/SplitProtocol/Sample/rr
      -- CP-element group 60: 	 branch_block_stmt_1335/forx_xbody_forx_xbody_PhiReq/phi_stmt_1561/phi_stmt_1561_sources/type_cast_1567/SplitProtocol/Update/$entry
      -- CP-element group 60: 	 branch_block_stmt_1335/forx_xbody_forx_xbody_PhiReq/phi_stmt_1561/phi_stmt_1561_sources/type_cast_1567/SplitProtocol/Update/cr
      -- 
    else_choice_transition_3133_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1582_branch_ack_0, ack => maxPool3D_CP_2658_elements(60)); -- 
    rr_3865_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3865_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(60), ack => type_cast_1567_inst_req_0); -- 
    cr_3870_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3870_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(60), ack => type_cast_1567_inst_req_1); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	244 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_1335/call_stmt_1605/call_stmt_1605_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_1335/call_stmt_1605/call_stmt_1605_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_1335/call_stmt_1605/call_stmt_1605_Sample/cra
      -- 
    cra_3150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1605_call_ack_0, ack => maxPool3D_CP_2658_elements(61)); -- 
    -- CP-element group 62:  fork  transition  place  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	244 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62: 	64 
    -- CP-element group 62: 	65 
    -- CP-element group 62: 	66 
    -- CP-element group 62: 	67 
    -- CP-element group 62: 	68 
    -- CP-element group 62:  members (25) 
      -- CP-element group 62: 	 branch_block_stmt_1335/call_stmt_1605__exit__
      -- CP-element group 62: 	 branch_block_stmt_1335/assign_stmt_1610_to_assign_stmt_1629__entry__
      -- CP-element group 62: 	 branch_block_stmt_1335/call_stmt_1605/$exit
      -- CP-element group 62: 	 branch_block_stmt_1335/call_stmt_1605/call_stmt_1605_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_1335/call_stmt_1605/call_stmt_1605_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_1335/call_stmt_1605/call_stmt_1605_Update/cca
      -- CP-element group 62: 	 branch_block_stmt_1335/assign_stmt_1610_to_assign_stmt_1629/$entry
      -- CP-element group 62: 	 branch_block_stmt_1335/assign_stmt_1610_to_assign_stmt_1629/type_cast_1609_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_1335/assign_stmt_1610_to_assign_stmt_1629/type_cast_1609_update_start_
      -- CP-element group 62: 	 branch_block_stmt_1335/assign_stmt_1610_to_assign_stmt_1629/type_cast_1609_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_1335/assign_stmt_1610_to_assign_stmt_1629/type_cast_1609_Sample/rr
      -- CP-element group 62: 	 branch_block_stmt_1335/assign_stmt_1610_to_assign_stmt_1629/type_cast_1609_Update/$entry
      -- CP-element group 62: 	 branch_block_stmt_1335/assign_stmt_1610_to_assign_stmt_1629/type_cast_1609_Update/cr
      -- CP-element group 62: 	 branch_block_stmt_1335/assign_stmt_1610_to_assign_stmt_1629/type_cast_1613_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_1335/assign_stmt_1610_to_assign_stmt_1629/type_cast_1613_update_start_
      -- CP-element group 62: 	 branch_block_stmt_1335/assign_stmt_1610_to_assign_stmt_1629/type_cast_1613_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_1335/assign_stmt_1610_to_assign_stmt_1629/type_cast_1613_Sample/rr
      -- CP-element group 62: 	 branch_block_stmt_1335/assign_stmt_1610_to_assign_stmt_1629/type_cast_1613_Update/$entry
      -- CP-element group 62: 	 branch_block_stmt_1335/assign_stmt_1610_to_assign_stmt_1629/type_cast_1613_Update/cr
      -- CP-element group 62: 	 branch_block_stmt_1335/assign_stmt_1610_to_assign_stmt_1629/type_cast_1617_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_1335/assign_stmt_1610_to_assign_stmt_1629/type_cast_1617_update_start_
      -- CP-element group 62: 	 branch_block_stmt_1335/assign_stmt_1610_to_assign_stmt_1629/type_cast_1617_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_1335/assign_stmt_1610_to_assign_stmt_1629/type_cast_1617_Sample/rr
      -- CP-element group 62: 	 branch_block_stmt_1335/assign_stmt_1610_to_assign_stmt_1629/type_cast_1617_Update/$entry
      -- CP-element group 62: 	 branch_block_stmt_1335/assign_stmt_1610_to_assign_stmt_1629/type_cast_1617_Update/cr
      -- 
    cca_3155_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1605_call_ack_1, ack => maxPool3D_CP_2658_elements(62)); -- 
    rr_3166_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3166_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(62), ack => type_cast_1609_inst_req_0); -- 
    cr_3171_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3171_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(62), ack => type_cast_1609_inst_req_1); -- 
    rr_3180_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3180_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(62), ack => type_cast_1613_inst_req_0); -- 
    cr_3185_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3185_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(62), ack => type_cast_1613_inst_req_1); -- 
    rr_3194_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3194_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(62), ack => type_cast_1617_inst_req_0); -- 
    cr_3199_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3199_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(62), ack => type_cast_1617_inst_req_1); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_1335/assign_stmt_1610_to_assign_stmt_1629/type_cast_1609_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_1335/assign_stmt_1610_to_assign_stmt_1629/type_cast_1609_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_1335/assign_stmt_1610_to_assign_stmt_1629/type_cast_1609_Sample/ra
      -- 
    ra_3167_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1609_inst_ack_0, ack => maxPool3D_CP_2658_elements(63)); -- 
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	62 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	69 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_1335/assign_stmt_1610_to_assign_stmt_1629/type_cast_1609_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_1335/assign_stmt_1610_to_assign_stmt_1629/type_cast_1609_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_1335/assign_stmt_1610_to_assign_stmt_1629/type_cast_1609_Update/ca
      -- 
    ca_3172_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1609_inst_ack_1, ack => maxPool3D_CP_2658_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	62 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_1335/assign_stmt_1610_to_assign_stmt_1629/type_cast_1613_sample_completed_
      -- CP-element group 65: 	 branch_block_stmt_1335/assign_stmt_1610_to_assign_stmt_1629/type_cast_1613_Sample/$exit
      -- CP-element group 65: 	 branch_block_stmt_1335/assign_stmt_1610_to_assign_stmt_1629/type_cast_1613_Sample/ra
      -- 
    ra_3181_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1613_inst_ack_0, ack => maxPool3D_CP_2658_elements(65)); -- 
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	62 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	69 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_1335/assign_stmt_1610_to_assign_stmt_1629/type_cast_1613_update_completed_
      -- CP-element group 66: 	 branch_block_stmt_1335/assign_stmt_1610_to_assign_stmt_1629/type_cast_1613_Update/$exit
      -- CP-element group 66: 	 branch_block_stmt_1335/assign_stmt_1610_to_assign_stmt_1629/type_cast_1613_Update/ca
      -- 
    ca_3186_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1613_inst_ack_1, ack => maxPool3D_CP_2658_elements(66)); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	62 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_1335/assign_stmt_1610_to_assign_stmt_1629/type_cast_1617_sample_completed_
      -- CP-element group 67: 	 branch_block_stmt_1335/assign_stmt_1610_to_assign_stmt_1629/type_cast_1617_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_1335/assign_stmt_1610_to_assign_stmt_1629/type_cast_1617_Sample/ra
      -- 
    ra_3195_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1617_inst_ack_0, ack => maxPool3D_CP_2658_elements(67)); -- 
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	62 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_1335/assign_stmt_1610_to_assign_stmt_1629/type_cast_1617_update_completed_
      -- CP-element group 68: 	 branch_block_stmt_1335/assign_stmt_1610_to_assign_stmt_1629/type_cast_1617_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_1335/assign_stmt_1610_to_assign_stmt_1629/type_cast_1617_Update/ca
      -- 
    ca_3200_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1617_inst_ack_1, ack => maxPool3D_CP_2658_elements(68)); -- 
    -- CP-element group 69:  join  transition  place  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	64 
    -- CP-element group 69: 	66 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69:  members (10) 
      -- CP-element group 69: 	 branch_block_stmt_1335/do_while_stmt_1648__entry__
      -- CP-element group 69: 	 branch_block_stmt_1335/merge_stmt_1631__exit__
      -- CP-element group 69: 	 branch_block_stmt_1335/forx_xend_whilex_xbody
      -- CP-element group 69: 	 branch_block_stmt_1335/assign_stmt_1610_to_assign_stmt_1629__exit__
      -- CP-element group 69: 	 branch_block_stmt_1335/assign_stmt_1610_to_assign_stmt_1629/$exit
      -- CP-element group 69: 	 branch_block_stmt_1335/forx_xend_whilex_xbody_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_1335/forx_xend_whilex_xbody_PhiReq/$exit
      -- CP-element group 69: 	 branch_block_stmt_1335/merge_stmt_1631_PhiReqMerge
      -- CP-element group 69: 	 branch_block_stmt_1335/merge_stmt_1631_PhiAck/$entry
      -- CP-element group 69: 	 branch_block_stmt_1335/merge_stmt_1631_PhiAck/$exit
      -- 
    maxPool3D_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool3D_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool3D_CP_2658_elements(64) & maxPool3D_CP_2658_elements(66) & maxPool3D_CP_2658_elements(68);
      gj_maxPool3D_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2658_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  transition  place  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	76 
    -- CP-element group 70:  members (2) 
      -- CP-element group 70: 	 branch_block_stmt_1335/do_while_stmt_1648/$entry
      -- CP-element group 70: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648__entry__
      -- 
    maxPool3D_CP_2658_elements(70) <= maxPool3D_CP_2658_elements(69);
    -- CP-element group 71:  merge  place  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	180 
    -- CP-element group 71:  members (1) 
      -- CP-element group 71: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648__exit__
      -- 
    -- Element group maxPool3D_CP_2658_elements(71) is bound as output of CP function.
    -- CP-element group 72:  merge  place  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	75 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_1335/do_while_stmt_1648/loop_back
      -- 
    -- Element group maxPool3D_CP_2658_elements(72) is bound as output of CP function.
    -- CP-element group 73:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	78 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	178 
    -- CP-element group 73: 	179 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_1335/do_while_stmt_1648/condition_done
      -- CP-element group 73: 	 branch_block_stmt_1335/do_while_stmt_1648/loop_taken/$entry
      -- CP-element group 73: 	 branch_block_stmt_1335/do_while_stmt_1648/loop_exit/$entry
      -- 
    maxPool3D_CP_2658_elements(73) <= maxPool3D_CP_2658_elements(78);
    -- CP-element group 74:  branch  place  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	177 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (1) 
      -- CP-element group 74: 	 branch_block_stmt_1335/do_while_stmt_1648/loop_body_done
      -- 
    maxPool3D_CP_2658_elements(74) <= maxPool3D_CP_2658_elements(177);
    -- CP-element group 75:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	72 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	87 
    -- CP-element group 75: 	108 
    -- CP-element group 75: 	129 
    -- CP-element group 75:  members (1) 
      -- CP-element group 75: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/back_edge_to_loop_body
      -- 
    maxPool3D_CP_2658_elements(75) <= maxPool3D_CP_2658_elements(72);
    -- CP-element group 76:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	70 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	89 
    -- CP-element group 76: 	110 
    -- CP-element group 76: 	131 
    -- CP-element group 76:  members (1) 
      -- CP-element group 76: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/first_time_through_loop_body
      -- 
    maxPool3D_CP_2658_elements(76) <= maxPool3D_CP_2658_elements(70);
    -- CP-element group 77:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	83 
    -- CP-element group 77: 	84 
    -- CP-element group 77: 	102 
    -- CP-element group 77: 	103 
    -- CP-element group 77: 	123 
    -- CP-element group 77: 	124 
    -- CP-element group 77: 	176 
    -- CP-element group 77:  members (2) 
      -- CP-element group 77: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/loop_body_start
      -- CP-element group 77: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/$entry
      -- 
    -- Element group maxPool3D_CP_2658_elements(77) is bound as output of CP function.
    -- CP-element group 78:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	82 
    -- CP-element group 78: 	171 
    -- CP-element group 78: 	175 
    -- CP-element group 78: 	176 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	73 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/condition_evaluated
      -- 
    condition_evaluated_3215_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_3215_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(78), ack => do_while_stmt_1648_branch_req_0); -- 
    maxPool3D_cp_element_group_78: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 15);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "maxPool3D_cp_element_group_78"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= maxPool3D_CP_2658_elements(82) & maxPool3D_CP_2658_elements(171) & maxPool3D_CP_2658_elements(175) & maxPool3D_CP_2658_elements(176);
      gj_maxPool3D_cp_element_group_78 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2658_elements(78), clk => clk, reset => reset); --
    end block;
    -- CP-element group 79:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	83 
    -- CP-element group 79: 	102 
    -- CP-element group 79: 	123 
    -- CP-element group 79: marked-predecessors 
    -- CP-element group 79: 	82 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	104 
    -- CP-element group 79: 	125 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/aggregated_phi_sample_req
      -- CP-element group 79: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/phi_stmt_1650_sample_start__ps
      -- 
    maxPool3D_cp_element_group_79: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "maxPool3D_cp_element_group_79"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= maxPool3D_CP_2658_elements(83) & maxPool3D_CP_2658_elements(102) & maxPool3D_CP_2658_elements(123) & maxPool3D_CP_2658_elements(82);
      gj_maxPool3D_cp_element_group_79 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2658_elements(79), clk => clk, reset => reset); --
    end block;
    -- CP-element group 80:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	85 
    -- CP-element group 80: 	105 
    -- CP-element group 80: 	126 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	161 
    -- CP-element group 80: 	165 
    -- CP-element group 80: 	169 
    -- CP-element group 80: 	173 
    -- CP-element group 80: 	177 
    -- CP-element group 80: marked-successors 
    -- CP-element group 80: 	83 
    -- CP-element group 80: 	102 
    -- CP-element group 80: 	123 
    -- CP-element group 80:  members (4) 
      -- CP-element group 80: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/phi_stmt_1650_sample_completed_
      -- CP-element group 80: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/aggregated_phi_sample_ack
      -- CP-element group 80: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/phi_stmt_1655_sample_completed_
      -- CP-element group 80: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/phi_stmt_1660_sample_completed_
      -- 
    maxPool3D_cp_element_group_80: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool3D_cp_element_group_80"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool3D_CP_2658_elements(85) & maxPool3D_CP_2658_elements(105) & maxPool3D_CP_2658_elements(126);
      gj_maxPool3D_cp_element_group_80 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2658_elements(80), clk => clk, reset => reset); --
    end block;
    -- CP-element group 81:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	84 
    -- CP-element group 81: 	103 
    -- CP-element group 81: 	124 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	106 
    -- CP-element group 81: 	127 
    -- CP-element group 81:  members (2) 
      -- CP-element group 81: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/aggregated_phi_update_req
      -- CP-element group 81: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/phi_stmt_1650_update_start__ps
      -- 
    maxPool3D_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool3D_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool3D_CP_2658_elements(84) & maxPool3D_CP_2658_elements(103) & maxPool3D_CP_2658_elements(124);
      gj_maxPool3D_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2658_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	86 
    -- CP-element group 82: 	107 
    -- CP-element group 82: 	128 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	78 
    -- CP-element group 82: marked-successors 
    -- CP-element group 82: 	79 
    -- CP-element group 82:  members (1) 
      -- CP-element group 82: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/aggregated_phi_update_ack
      -- 
    maxPool3D_cp_element_group_82: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool3D_cp_element_group_82"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool3D_CP_2658_elements(86) & maxPool3D_CP_2658_elements(107) & maxPool3D_CP_2658_elements(128);
      gj_maxPool3D_cp_element_group_82 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2658_elements(82), clk => clk, reset => reset); --
    end block;
    -- CP-element group 83:  join  transition  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	77 
    -- CP-element group 83: marked-predecessors 
    -- CP-element group 83: 	80 
    -- CP-element group 83: 	171 
    -- CP-element group 83: 	175 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	79 
    -- CP-element group 83:  members (1) 
      -- CP-element group 83: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/phi_stmt_1650_sample_start_
      -- 
    maxPool3D_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 1,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "maxPool3D_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= maxPool3D_CP_2658_elements(77) & maxPool3D_CP_2658_elements(80) & maxPool3D_CP_2658_elements(171) & maxPool3D_CP_2658_elements(175);
      gj_maxPool3D_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2658_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  join  transition  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	77 
    -- CP-element group 84: marked-predecessors 
    -- CP-element group 84: 	86 
    -- CP-element group 84: 	154 
    -- CP-element group 84: 	174 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	81 
    -- CP-element group 84:  members (1) 
      -- CP-element group 84: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/phi_stmt_1650_update_start_
      -- 
    maxPool3D_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "maxPool3D_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= maxPool3D_CP_2658_elements(77) & maxPool3D_CP_2658_elements(86) & maxPool3D_CP_2658_elements(154) & maxPool3D_CP_2658_elements(174);
      gj_maxPool3D_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2658_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  join  transition  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	80 
    -- CP-element group 85:  members (1) 
      -- CP-element group 85: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/phi_stmt_1650_sample_completed__ps
      -- 
    -- Element group maxPool3D_CP_2658_elements(85) is bound as output of CP function.
    -- CP-element group 86:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	82 
    -- CP-element group 86: 	152 
    -- CP-element group 86: 	172 
    -- CP-element group 86: marked-successors 
    -- CP-element group 86: 	84 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/phi_stmt_1650_update_completed_
      -- CP-element group 86: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/phi_stmt_1650_update_completed__ps
      -- 
    -- Element group maxPool3D_CP_2658_elements(86) is bound as output of CP function.
    -- CP-element group 87:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	75 
    -- CP-element group 87: successors 
    -- CP-element group 87:  members (1) 
      -- CP-element group 87: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/phi_stmt_1650_loopback_trigger
      -- 
    maxPool3D_CP_2658_elements(87) <= maxPool3D_CP_2658_elements(75);
    -- CP-element group 88:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (2) 
      -- CP-element group 88: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/phi_stmt_1650_loopback_sample_req_ps
      -- CP-element group 88: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/phi_stmt_1650_loopback_sample_req
      -- 
    phi_stmt_1650_loopback_sample_req_3230_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1650_loopback_sample_req_3230_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(88), ack => phi_stmt_1650_req_0); -- 
    -- Element group maxPool3D_CP_2658_elements(88) is bound as output of CP function.
    -- CP-element group 89:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	76 
    -- CP-element group 89: successors 
    -- CP-element group 89:  members (1) 
      -- CP-element group 89: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/phi_stmt_1650_entry_trigger
      -- 
    maxPool3D_CP_2658_elements(89) <= maxPool3D_CP_2658_elements(76);
    -- CP-element group 90:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: successors 
    -- CP-element group 90:  members (2) 
      -- CP-element group 90: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/phi_stmt_1650_entry_sample_req_ps
      -- CP-element group 90: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/phi_stmt_1650_entry_sample_req
      -- 
    phi_stmt_1650_entry_sample_req_3233_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1650_entry_sample_req_3233_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(90), ack => phi_stmt_1650_req_1); -- 
    -- Element group maxPool3D_CP_2658_elements(90) is bound as output of CP function.
    -- CP-element group 91:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: successors 
    -- CP-element group 91:  members (2) 
      -- CP-element group 91: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/phi_stmt_1650_phi_mux_ack
      -- CP-element group 91: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/phi_stmt_1650_phi_mux_ack_ps
      -- 
    phi_stmt_1650_phi_mux_ack_3236_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1650_ack_0, ack => maxPool3D_CP_2658_elements(91)); -- 
    -- CP-element group 92:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	94 
    -- CP-element group 92:  members (1) 
      -- CP-element group 92: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1653_sample_start__ps
      -- 
    -- Element group maxPool3D_CP_2658_elements(92) is bound as output of CP function.
    -- CP-element group 93:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (1) 
      -- CP-element group 93: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1653_update_start__ps
      -- 
    -- Element group maxPool3D_CP_2658_elements(93) is bound as output of CP function.
    -- CP-element group 94:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	92 
    -- CP-element group 94: marked-predecessors 
    -- CP-element group 94: 	96 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	96 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1653_sample_start_
      -- CP-element group 94: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1653_Sample/rr
      -- CP-element group 94: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1653_Sample/$entry
      -- 
    rr_3249_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3249_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(94), ack => type_cast_1653_inst_req_0); -- 
    maxPool3D_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool3D_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2658_elements(92) & maxPool3D_CP_2658_elements(96);
      gj_maxPool3D_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2658_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: marked-predecessors 
    -- CP-element group 95: 	97 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	97 
    -- CP-element group 95:  members (3) 
      -- CP-element group 95: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1653_Update/cr
      -- CP-element group 95: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1653_update_start_
      -- CP-element group 95: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1653_Update/$entry
      -- 
    cr_3254_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3254_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(95), ack => type_cast_1653_inst_req_1); -- 
    maxPool3D_cp_element_group_95: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool3D_cp_element_group_95"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2658_elements(93) & maxPool3D_CP_2658_elements(97);
      gj_maxPool3D_cp_element_group_95 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2658_elements(95), clk => clk, reset => reset); --
    end block;
    -- CP-element group 96:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	94 
    -- CP-element group 96: successors 
    -- CP-element group 96: marked-successors 
    -- CP-element group 96: 	94 
    -- CP-element group 96:  members (4) 
      -- CP-element group 96: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1653_sample_completed__ps
      -- CP-element group 96: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1653_sample_completed_
      -- CP-element group 96: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1653_Sample/ra
      -- CP-element group 96: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1653_Sample/$exit
      -- 
    ra_3250_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1653_inst_ack_0, ack => maxPool3D_CP_2658_elements(96)); -- 
    -- CP-element group 97:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: successors 
    -- CP-element group 97: marked-successors 
    -- CP-element group 97: 	95 
    -- CP-element group 97:  members (4) 
      -- CP-element group 97: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1653_Update/ca
      -- CP-element group 97: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1653_update_completed__ps
      -- CP-element group 97: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1653_Update/$exit
      -- CP-element group 97: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1653_update_completed_
      -- 
    ca_3255_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1653_inst_ack_1, ack => maxPool3D_CP_2658_elements(97)); -- 
    -- CP-element group 98:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: successors 
    -- CP-element group 98:  members (4) 
      -- CP-element group 98: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/R_rowx_x1_at_entry_1654_sample_start_
      -- CP-element group 98: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/R_rowx_x1_at_entry_1654_sample_start__ps
      -- CP-element group 98: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/R_rowx_x1_at_entry_1654_sample_completed__ps
      -- CP-element group 98: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/R_rowx_x1_at_entry_1654_sample_completed_
      -- 
    -- Element group maxPool3D_CP_2658_elements(98) is bound as output of CP function.
    -- CP-element group 99:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	101 
    -- CP-element group 99:  members (2) 
      -- CP-element group 99: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/R_rowx_x1_at_entry_1654_update_start__ps
      -- CP-element group 99: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/R_rowx_x1_at_entry_1654_update_start_
      -- 
    -- Element group maxPool3D_CP_2658_elements(99) is bound as output of CP function.
    -- CP-element group 100:  join  transition  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	101 
    -- CP-element group 100: successors 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/R_rowx_x1_at_entry_1654_update_completed__ps
      -- 
    maxPool3D_CP_2658_elements(100) <= maxPool3D_CP_2658_elements(101);
    -- CP-element group 101:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	99 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	100 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/R_rowx_x1_at_entry_1654_update_completed_
      -- 
    -- Element group maxPool3D_CP_2658_elements(101) is a control-delay.
    cp_element_101_delay: control_delay_element  generic map(name => " 101_delay", delay_value => 1)  port map(req => maxPool3D_CP_2658_elements(99), ack => maxPool3D_CP_2658_elements(101), clk => clk, reset =>reset);
    -- CP-element group 102:  join  transition  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	77 
    -- CP-element group 102: marked-predecessors 
    -- CP-element group 102: 	80 
    -- CP-element group 102: 	163 
    -- CP-element group 102: 	167 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	79 
    -- CP-element group 102:  members (1) 
      -- CP-element group 102: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/phi_stmt_1655_sample_start_
      -- 
    maxPool3D_cp_element_group_102: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 1,2 => 0,3 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_102"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= maxPool3D_CP_2658_elements(77) & maxPool3D_CP_2658_elements(80) & maxPool3D_CP_2658_elements(163) & maxPool3D_CP_2658_elements(167);
      gj_maxPool3D_cp_element_group_102 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2658_elements(102), clk => clk, reset => reset); --
    end block;
    -- CP-element group 103:  join  transition  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	77 
    -- CP-element group 103: marked-predecessors 
    -- CP-element group 103: 	107 
    -- CP-element group 103: 	150 
    -- CP-element group 103: 	166 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	81 
    -- CP-element group 103:  members (1) 
      -- CP-element group 103: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/phi_stmt_1655_update_start_
      -- 
    maxPool3D_cp_element_group_103: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_103"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= maxPool3D_CP_2658_elements(77) & maxPool3D_CP_2658_elements(107) & maxPool3D_CP_2658_elements(150) & maxPool3D_CP_2658_elements(166);
      gj_maxPool3D_cp_element_group_103 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2658_elements(103), clk => clk, reset => reset); --
    end block;
    -- CP-element group 104:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	79 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (1) 
      -- CP-element group 104: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/phi_stmt_1655_sample_start__ps
      -- 
    maxPool3D_CP_2658_elements(104) <= maxPool3D_CP_2658_elements(79);
    -- CP-element group 105:  join  transition  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	80 
    -- CP-element group 105:  members (1) 
      -- CP-element group 105: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/phi_stmt_1655_sample_completed__ps
      -- 
    -- Element group maxPool3D_CP_2658_elements(105) is bound as output of CP function.
    -- CP-element group 106:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	81 
    -- CP-element group 106: successors 
    -- CP-element group 106:  members (1) 
      -- CP-element group 106: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/phi_stmt_1655_update_start__ps
      -- 
    maxPool3D_CP_2658_elements(106) <= maxPool3D_CP_2658_elements(81);
    -- CP-element group 107:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	82 
    -- CP-element group 107: 	148 
    -- CP-element group 107: 	164 
    -- CP-element group 107: marked-successors 
    -- CP-element group 107: 	103 
    -- CP-element group 107:  members (2) 
      -- CP-element group 107: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/phi_stmt_1655_update_completed__ps
      -- CP-element group 107: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/phi_stmt_1655_update_completed_
      -- 
    -- Element group maxPool3D_CP_2658_elements(107) is bound as output of CP function.
    -- CP-element group 108:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	75 
    -- CP-element group 108: successors 
    -- CP-element group 108:  members (1) 
      -- CP-element group 108: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/phi_stmt_1655_loopback_trigger
      -- 
    maxPool3D_CP_2658_elements(108) <= maxPool3D_CP_2658_elements(75);
    -- CP-element group 109:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: successors 
    -- CP-element group 109:  members (2) 
      -- CP-element group 109: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/phi_stmt_1655_loopback_sample_req_ps
      -- CP-element group 109: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/phi_stmt_1655_loopback_sample_req
      -- 
    phi_stmt_1655_loopback_sample_req_3274_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1655_loopback_sample_req_3274_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(109), ack => phi_stmt_1655_req_0); -- 
    -- Element group maxPool3D_CP_2658_elements(109) is bound as output of CP function.
    -- CP-element group 110:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	76 
    -- CP-element group 110: successors 
    -- CP-element group 110:  members (1) 
      -- CP-element group 110: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/phi_stmt_1655_entry_trigger
      -- 
    maxPool3D_CP_2658_elements(110) <= maxPool3D_CP_2658_elements(76);
    -- CP-element group 111:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: successors 
    -- CP-element group 111:  members (2) 
      -- CP-element group 111: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/phi_stmt_1655_entry_sample_req_ps
      -- CP-element group 111: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/phi_stmt_1655_entry_sample_req
      -- 
    phi_stmt_1655_entry_sample_req_3277_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1655_entry_sample_req_3277_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(111), ack => phi_stmt_1655_req_1); -- 
    -- Element group maxPool3D_CP_2658_elements(111) is bound as output of CP function.
    -- CP-element group 112:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: successors 
    -- CP-element group 112:  members (2) 
      -- CP-element group 112: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/phi_stmt_1655_phi_mux_ack_ps
      -- CP-element group 112: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/phi_stmt_1655_phi_mux_ack
      -- 
    phi_stmt_1655_phi_mux_ack_3280_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1655_ack_0, ack => maxPool3D_CP_2658_elements(112)); -- 
    -- CP-element group 113:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (1) 
      -- CP-element group 113: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1658_sample_start__ps
      -- 
    -- Element group maxPool3D_CP_2658_elements(113) is bound as output of CP function.
    -- CP-element group 114:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	116 
    -- CP-element group 114:  members (1) 
      -- CP-element group 114: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1658_update_start__ps
      -- 
    -- Element group maxPool3D_CP_2658_elements(114) is bound as output of CP function.
    -- CP-element group 115:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: marked-predecessors 
    -- CP-element group 115: 	117 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	117 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1658_Sample/rr
      -- CP-element group 115: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1658_Sample/$entry
      -- CP-element group 115: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1658_sample_start_
      -- 
    rr_3293_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3293_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(115), ack => type_cast_1658_inst_req_0); -- 
    maxPool3D_cp_element_group_115: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_115"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2658_elements(113) & maxPool3D_CP_2658_elements(117);
      gj_maxPool3D_cp_element_group_115 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2658_elements(115), clk => clk, reset => reset); --
    end block;
    -- CP-element group 116:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	114 
    -- CP-element group 116: marked-predecessors 
    -- CP-element group 116: 	118 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	118 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1658_update_start_
      -- CP-element group 116: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1658_Update/$entry
      -- CP-element group 116: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1658_Update/cr
      -- 
    cr_3298_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3298_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(116), ack => type_cast_1658_inst_req_1); -- 
    maxPool3D_cp_element_group_116: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_116"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2658_elements(114) & maxPool3D_CP_2658_elements(118);
      gj_maxPool3D_cp_element_group_116 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2658_elements(116), clk => clk, reset => reset); --
    end block;
    -- CP-element group 117:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	115 
    -- CP-element group 117: successors 
    -- CP-element group 117: marked-successors 
    -- CP-element group 117: 	115 
    -- CP-element group 117:  members (4) 
      -- CP-element group 117: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1658_sample_completed__ps
      -- CP-element group 117: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1658_Sample/ra
      -- CP-element group 117: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1658_Sample/$exit
      -- CP-element group 117: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1658_sample_completed_
      -- 
    ra_3294_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1658_inst_ack_0, ack => maxPool3D_CP_2658_elements(117)); -- 
    -- CP-element group 118:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	116 
    -- CP-element group 118: successors 
    -- CP-element group 118: marked-successors 
    -- CP-element group 118: 	116 
    -- CP-element group 118:  members (4) 
      -- CP-element group 118: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1658_update_completed_
      -- CP-element group 118: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1658_update_completed__ps
      -- CP-element group 118: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1658_Update/$exit
      -- CP-element group 118: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1658_Update/ca
      -- 
    ca_3299_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1658_inst_ack_1, ack => maxPool3D_CP_2658_elements(118)); -- 
    -- CP-element group 119:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: successors 
    -- CP-element group 119:  members (4) 
      -- CP-element group 119: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/R_colx_x1_at_entry_1659_sample_completed_
      -- CP-element group 119: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/R_colx_x1_at_entry_1659_sample_start_
      -- CP-element group 119: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/R_colx_x1_at_entry_1659_sample_completed__ps
      -- CP-element group 119: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/R_colx_x1_at_entry_1659_sample_start__ps
      -- 
    -- Element group maxPool3D_CP_2658_elements(119) is bound as output of CP function.
    -- CP-element group 120:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	122 
    -- CP-element group 120:  members (2) 
      -- CP-element group 120: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/R_colx_x1_at_entry_1659_update_start_
      -- CP-element group 120: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/R_colx_x1_at_entry_1659_update_start__ps
      -- 
    -- Element group maxPool3D_CP_2658_elements(120) is bound as output of CP function.
    -- CP-element group 121:  join  transition  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	122 
    -- CP-element group 121: successors 
    -- CP-element group 121:  members (1) 
      -- CP-element group 121: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/R_colx_x1_at_entry_1659_update_completed__ps
      -- 
    maxPool3D_CP_2658_elements(121) <= maxPool3D_CP_2658_elements(122);
    -- CP-element group 122:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	120 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	121 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/R_colx_x1_at_entry_1659_update_completed_
      -- 
    -- Element group maxPool3D_CP_2658_elements(122) is a control-delay.
    cp_element_122_delay: control_delay_element  generic map(name => " 122_delay", delay_value => 1)  port map(req => maxPool3D_CP_2658_elements(120), ack => maxPool3D_CP_2658_elements(122), clk => clk, reset =>reset);
    -- CP-element group 123:  join  transition  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	77 
    -- CP-element group 123: marked-predecessors 
    -- CP-element group 123: 	80 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	79 
    -- CP-element group 123:  members (1) 
      -- CP-element group 123: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/phi_stmt_1660_sample_start_
      -- 
    maxPool3D_cp_element_group_123: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_123"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2658_elements(77) & maxPool3D_CP_2658_elements(80);
      gj_maxPool3D_cp_element_group_123 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2658_elements(123), clk => clk, reset => reset); --
    end block;
    -- CP-element group 124:  join  transition  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	77 
    -- CP-element group 124: marked-predecessors 
    -- CP-element group 124: 	128 
    -- CP-element group 124: 	146 
    -- CP-element group 124: 	162 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	81 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/phi_stmt_1660_update_start_
      -- 
    maxPool3D_cp_element_group_124: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_124"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= maxPool3D_CP_2658_elements(77) & maxPool3D_CP_2658_elements(128) & maxPool3D_CP_2658_elements(146) & maxPool3D_CP_2658_elements(162);
      gj_maxPool3D_cp_element_group_124 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2658_elements(124), clk => clk, reset => reset); --
    end block;
    -- CP-element group 125:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	79 
    -- CP-element group 125: successors 
    -- CP-element group 125:  members (1) 
      -- CP-element group 125: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/phi_stmt_1660_sample_start__ps
      -- 
    maxPool3D_CP_2658_elements(125) <= maxPool3D_CP_2658_elements(79);
    -- CP-element group 126:  join  transition  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	80 
    -- CP-element group 126:  members (1) 
      -- CP-element group 126: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/phi_stmt_1660_sample_completed__ps
      -- 
    -- Element group maxPool3D_CP_2658_elements(126) is bound as output of CP function.
    -- CP-element group 127:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	81 
    -- CP-element group 127: successors 
    -- CP-element group 127:  members (1) 
      -- CP-element group 127: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/phi_stmt_1660_update_start__ps
      -- 
    maxPool3D_CP_2658_elements(127) <= maxPool3D_CP_2658_elements(81);
    -- CP-element group 128:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	82 
    -- CP-element group 128: 	144 
    -- CP-element group 128: 	160 
    -- CP-element group 128: marked-successors 
    -- CP-element group 128: 	124 
    -- CP-element group 128:  members (2) 
      -- CP-element group 128: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/phi_stmt_1660_update_completed_
      -- CP-element group 128: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/phi_stmt_1660_update_completed__ps
      -- 
    -- Element group maxPool3D_CP_2658_elements(128) is bound as output of CP function.
    -- CP-element group 129:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	75 
    -- CP-element group 129: successors 
    -- CP-element group 129:  members (1) 
      -- CP-element group 129: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/phi_stmt_1660_loopback_trigger
      -- 
    maxPool3D_CP_2658_elements(129) <= maxPool3D_CP_2658_elements(75);
    -- CP-element group 130:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: successors 
    -- CP-element group 130:  members (2) 
      -- CP-element group 130: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/phi_stmt_1660_loopback_sample_req_ps
      -- CP-element group 130: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/phi_stmt_1660_loopback_sample_req
      -- 
    phi_stmt_1660_loopback_sample_req_3318_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1660_loopback_sample_req_3318_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(130), ack => phi_stmt_1660_req_0); -- 
    -- Element group maxPool3D_CP_2658_elements(130) is bound as output of CP function.
    -- CP-element group 131:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	76 
    -- CP-element group 131: successors 
    -- CP-element group 131:  members (1) 
      -- CP-element group 131: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/phi_stmt_1660_entry_trigger
      -- 
    maxPool3D_CP_2658_elements(131) <= maxPool3D_CP_2658_elements(76);
    -- CP-element group 132:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: successors 
    -- CP-element group 132:  members (2) 
      -- CP-element group 132: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/phi_stmt_1660_entry_sample_req_ps
      -- CP-element group 132: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/phi_stmt_1660_entry_sample_req
      -- 
    phi_stmt_1660_entry_sample_req_3321_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1660_entry_sample_req_3321_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(132), ack => phi_stmt_1660_req_1); -- 
    -- Element group maxPool3D_CP_2658_elements(132) is bound as output of CP function.
    -- CP-element group 133:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: successors 
    -- CP-element group 133:  members (2) 
      -- CP-element group 133: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/phi_stmt_1660_phi_mux_ack_ps
      -- CP-element group 133: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/phi_stmt_1660_phi_mux_ack
      -- 
    phi_stmt_1660_phi_mux_ack_3324_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1660_ack_0, ack => maxPool3D_CP_2658_elements(133)); -- 
    -- CP-element group 134:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	136 
    -- CP-element group 134:  members (1) 
      -- CP-element group 134: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1663_sample_start__ps
      -- 
    -- Element group maxPool3D_CP_2658_elements(134) is bound as output of CP function.
    -- CP-element group 135:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	137 
    -- CP-element group 135:  members (1) 
      -- CP-element group 135: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1663_update_start__ps
      -- 
    -- Element group maxPool3D_CP_2658_elements(135) is bound as output of CP function.
    -- CP-element group 136:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	134 
    -- CP-element group 136: marked-predecessors 
    -- CP-element group 136: 	138 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	138 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1663_Sample/rr
      -- CP-element group 136: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1663_Sample/$entry
      -- CP-element group 136: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1663_sample_start_
      -- 
    rr_3337_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3337_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(136), ack => type_cast_1663_inst_req_0); -- 
    maxPool3D_cp_element_group_136: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_136"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2658_elements(134) & maxPool3D_CP_2658_elements(138);
      gj_maxPool3D_cp_element_group_136 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2658_elements(136), clk => clk, reset => reset); --
    end block;
    -- CP-element group 137:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	135 
    -- CP-element group 137: marked-predecessors 
    -- CP-element group 137: 	139 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	139 
    -- CP-element group 137:  members (3) 
      -- CP-element group 137: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1663_Update/cr
      -- CP-element group 137: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1663_Update/$entry
      -- CP-element group 137: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1663_update_start_
      -- 
    cr_3342_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3342_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(137), ack => type_cast_1663_inst_req_1); -- 
    maxPool3D_cp_element_group_137: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_137"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2658_elements(135) & maxPool3D_CP_2658_elements(139);
      gj_maxPool3D_cp_element_group_137 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2658_elements(137), clk => clk, reset => reset); --
    end block;
    -- CP-element group 138:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	136 
    -- CP-element group 138: successors 
    -- CP-element group 138: marked-successors 
    -- CP-element group 138: 	136 
    -- CP-element group 138:  members (4) 
      -- CP-element group 138: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1663_Sample/ra
      -- CP-element group 138: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1663_Sample/$exit
      -- CP-element group 138: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1663_sample_completed_
      -- CP-element group 138: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1663_sample_completed__ps
      -- 
    ra_3338_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1663_inst_ack_0, ack => maxPool3D_CP_2658_elements(138)); -- 
    -- CP-element group 139:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	137 
    -- CP-element group 139: successors 
    -- CP-element group 139: marked-successors 
    -- CP-element group 139: 	137 
    -- CP-element group 139:  members (4) 
      -- CP-element group 139: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1663_Update/ca
      -- CP-element group 139: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1663_Update/$exit
      -- CP-element group 139: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1663_update_completed_
      -- CP-element group 139: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1663_update_completed__ps
      -- 
    ca_3343_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1663_inst_ack_1, ack => maxPool3D_CP_2658_elements(139)); -- 
    -- CP-element group 140:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: successors 
    -- CP-element group 140:  members (4) 
      -- CP-element group 140: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/R_chlx_x0_at_entry_1664_sample_completed_
      -- CP-element group 140: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/R_chlx_x0_at_entry_1664_sample_start_
      -- CP-element group 140: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/R_chlx_x0_at_entry_1664_sample_completed__ps
      -- CP-element group 140: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/R_chlx_x0_at_entry_1664_sample_start__ps
      -- 
    -- Element group maxPool3D_CP_2658_elements(140) is bound as output of CP function.
    -- CP-element group 141:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	143 
    -- CP-element group 141:  members (2) 
      -- CP-element group 141: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/R_chlx_x0_at_entry_1664_update_start_
      -- CP-element group 141: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/R_chlx_x0_at_entry_1664_update_start__ps
      -- 
    -- Element group maxPool3D_CP_2658_elements(141) is bound as output of CP function.
    -- CP-element group 142:  join  transition  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	143 
    -- CP-element group 142: successors 
    -- CP-element group 142:  members (1) 
      -- CP-element group 142: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/R_chlx_x0_at_entry_1664_update_completed__ps
      -- 
    maxPool3D_CP_2658_elements(142) <= maxPool3D_CP_2658_elements(143);
    -- CP-element group 143:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	141 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	142 
    -- CP-element group 143:  members (1) 
      -- CP-element group 143: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/R_chlx_x0_at_entry_1664_update_completed_
      -- 
    -- Element group maxPool3D_CP_2658_elements(143) is a control-delay.
    cp_element_143_delay: control_delay_element  generic map(name => " 143_delay", delay_value => 1)  port map(req => maxPool3D_CP_2658_elements(141), ack => maxPool3D_CP_2658_elements(143), clk => clk, reset =>reset);
    -- CP-element group 144:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	128 
    -- CP-element group 144: marked-predecessors 
    -- CP-element group 144: 	146 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	146 
    -- CP-element group 144:  members (3) 
      -- CP-element group 144: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1668_Sample/$entry
      -- CP-element group 144: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1668_Sample/rr
      -- CP-element group 144: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1668_sample_start_
      -- 
    rr_3360_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3360_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(144), ack => type_cast_1668_inst_req_0); -- 
    maxPool3D_cp_element_group_144: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_144"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2658_elements(128) & maxPool3D_CP_2658_elements(146);
      gj_maxPool3D_cp_element_group_144 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2658_elements(144), clk => clk, reset => reset); --
    end block;
    -- CP-element group 145:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: marked-predecessors 
    -- CP-element group 145: 	147 
    -- CP-element group 145: 	158 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	147 
    -- CP-element group 145:  members (3) 
      -- CP-element group 145: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1668_Update/$entry
      -- CP-element group 145: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1668_Update/cr
      -- CP-element group 145: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1668_update_start_
      -- 
    cr_3365_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3365_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(145), ack => type_cast_1668_inst_req_1); -- 
    maxPool3D_cp_element_group_145: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_145"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2658_elements(147) & maxPool3D_CP_2658_elements(158);
      gj_maxPool3D_cp_element_group_145 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2658_elements(145), clk => clk, reset => reset); --
    end block;
    -- CP-element group 146:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	144 
    -- CP-element group 146: successors 
    -- CP-element group 146: marked-successors 
    -- CP-element group 146: 	124 
    -- CP-element group 146: 	144 
    -- CP-element group 146:  members (3) 
      -- CP-element group 146: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1668_Sample/$exit
      -- CP-element group 146: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1668_Sample/ra
      -- CP-element group 146: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1668_sample_completed_
      -- 
    ra_3361_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1668_inst_ack_0, ack => maxPool3D_CP_2658_elements(146)); -- 
    -- CP-element group 147:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	145 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	156 
    -- CP-element group 147: marked-successors 
    -- CP-element group 147: 	145 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1668_update_completed_
      -- CP-element group 147: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1668_Update/$exit
      -- CP-element group 147: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1668_Update/ca
      -- 
    ca_3366_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1668_inst_ack_1, ack => maxPool3D_CP_2658_elements(147)); -- 
    -- CP-element group 148:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	107 
    -- CP-element group 148: marked-predecessors 
    -- CP-element group 148: 	150 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	150 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1672_sample_start_
      -- CP-element group 148: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1672_Sample/rr
      -- CP-element group 148: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1672_Sample/$entry
      -- 
    rr_3374_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3374_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(148), ack => type_cast_1672_inst_req_0); -- 
    maxPool3D_cp_element_group_148: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_148"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2658_elements(107) & maxPool3D_CP_2658_elements(150);
      gj_maxPool3D_cp_element_group_148 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2658_elements(148), clk => clk, reset => reset); --
    end block;
    -- CP-element group 149:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: marked-predecessors 
    -- CP-element group 149: 	151 
    -- CP-element group 149: 	158 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	151 
    -- CP-element group 149:  members (3) 
      -- CP-element group 149: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1672_update_start_
      -- CP-element group 149: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1672_Update/cr
      -- CP-element group 149: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1672_Update/$entry
      -- 
    cr_3379_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3379_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(149), ack => type_cast_1672_inst_req_1); -- 
    maxPool3D_cp_element_group_149: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_149"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2658_elements(151) & maxPool3D_CP_2658_elements(158);
      gj_maxPool3D_cp_element_group_149 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2658_elements(149), clk => clk, reset => reset); --
    end block;
    -- CP-element group 150:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	148 
    -- CP-element group 150: successors 
    -- CP-element group 150: marked-successors 
    -- CP-element group 150: 	103 
    -- CP-element group 150: 	148 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1672_sample_completed_
      -- CP-element group 150: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1672_Sample/ra
      -- CP-element group 150: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1672_Sample/$exit
      -- 
    ra_3375_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1672_inst_ack_0, ack => maxPool3D_CP_2658_elements(150)); -- 
    -- CP-element group 151:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	149 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	156 
    -- CP-element group 151: marked-successors 
    -- CP-element group 151: 	149 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1672_Update/ca
      -- CP-element group 151: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1672_Update/$exit
      -- CP-element group 151: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1672_update_completed_
      -- 
    ca_3380_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1672_inst_ack_1, ack => maxPool3D_CP_2658_elements(151)); -- 
    -- CP-element group 152:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	86 
    -- CP-element group 152: marked-predecessors 
    -- CP-element group 152: 	154 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	154 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1676_Sample/rr
      -- CP-element group 152: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1676_Sample/$entry
      -- CP-element group 152: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1676_sample_start_
      -- 
    rr_3388_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3388_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(152), ack => type_cast_1676_inst_req_0); -- 
    maxPool3D_cp_element_group_152: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_152"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2658_elements(86) & maxPool3D_CP_2658_elements(154);
      gj_maxPool3D_cp_element_group_152 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2658_elements(152), clk => clk, reset => reset); --
    end block;
    -- CP-element group 153:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: marked-predecessors 
    -- CP-element group 153: 	155 
    -- CP-element group 153: 	158 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	155 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1676_Update/cr
      -- CP-element group 153: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1676_Update/$entry
      -- CP-element group 153: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1676_update_start_
      -- 
    cr_3393_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3393_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(153), ack => type_cast_1676_inst_req_1); -- 
    maxPool3D_cp_element_group_153: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_153"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2658_elements(155) & maxPool3D_CP_2658_elements(158);
      gj_maxPool3D_cp_element_group_153 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2658_elements(153), clk => clk, reset => reset); --
    end block;
    -- CP-element group 154:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	152 
    -- CP-element group 154: successors 
    -- CP-element group 154: marked-successors 
    -- CP-element group 154: 	84 
    -- CP-element group 154: 	152 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1676_Sample/ra
      -- CP-element group 154: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1676_Sample/$exit
      -- CP-element group 154: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1676_sample_completed_
      -- 
    ra_3389_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1676_inst_ack_0, ack => maxPool3D_CP_2658_elements(154)); -- 
    -- CP-element group 155:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	153 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	156 
    -- CP-element group 155: marked-successors 
    -- CP-element group 155: 	153 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1676_Update/ca
      -- CP-element group 155: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1676_Update/$exit
      -- CP-element group 155: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1676_update_completed_
      -- 
    ca_3394_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1676_inst_ack_1, ack => maxPool3D_CP_2658_elements(155)); -- 
    -- CP-element group 156:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	147 
    -- CP-element group 156: 	151 
    -- CP-element group 156: 	155 
    -- CP-element group 156: marked-predecessors 
    -- CP-element group 156: 	158 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	158 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/call_stmt_1745_Sample/crr
      -- CP-element group 156: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/call_stmt_1745_Sample/$entry
      -- CP-element group 156: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/call_stmt_1745_sample_start_
      -- 
    crr_3402_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3402_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(156), ack => call_stmt_1745_call_req_0); -- 
    maxPool3D_cp_element_group_156: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_156"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= maxPool3D_CP_2658_elements(147) & maxPool3D_CP_2658_elements(151) & maxPool3D_CP_2658_elements(155) & maxPool3D_CP_2658_elements(158);
      gj_maxPool3D_cp_element_group_156 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2658_elements(156), clk => clk, reset => reset); --
    end block;
    -- CP-element group 157:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: marked-predecessors 
    -- CP-element group 157: 	159 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	159 
    -- CP-element group 157:  members (3) 
      -- CP-element group 157: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/call_stmt_1745_Update/ccr
      -- CP-element group 157: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/call_stmt_1745_Update/$entry
      -- CP-element group 157: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/call_stmt_1745_update_start_
      -- 
    ccr_3407_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3407_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(157), ack => call_stmt_1745_call_req_1); -- 
    maxPool3D_cp_element_group_157: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_157"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= maxPool3D_CP_2658_elements(159);
      gj_maxPool3D_cp_element_group_157 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2658_elements(157), clk => clk, reset => reset); --
    end block;
    -- CP-element group 158:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	156 
    -- CP-element group 158: successors 
    -- CP-element group 158: marked-successors 
    -- CP-element group 158: 	145 
    -- CP-element group 158: 	149 
    -- CP-element group 158: 	153 
    -- CP-element group 158: 	156 
    -- CP-element group 158:  members (3) 
      -- CP-element group 158: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/call_stmt_1745_Sample/$exit
      -- CP-element group 158: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/call_stmt_1745_Sample/cra
      -- CP-element group 158: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/call_stmt_1745_sample_completed_
      -- 
    cra_3403_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1745_call_ack_0, ack => maxPool3D_CP_2658_elements(158)); -- 
    -- CP-element group 159:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	157 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	177 
    -- CP-element group 159: marked-successors 
    -- CP-element group 159: 	157 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/call_stmt_1745_Update/cca
      -- CP-element group 159: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/call_stmt_1745_Update/$exit
      -- CP-element group 159: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/call_stmt_1745_update_completed_
      -- 
    cca_3408_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1745_call_ack_1, ack => maxPool3D_CP_2658_elements(159)); -- 
    -- CP-element group 160:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	128 
    -- CP-element group 160: marked-predecessors 
    -- CP-element group 160: 	162 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	162 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1759_sample_start_
      -- CP-element group 160: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1759_Sample/$entry
      -- CP-element group 160: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1759_Sample/rr
      -- 
    rr_3416_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3416_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(160), ack => type_cast_1759_inst_req_0); -- 
    maxPool3D_cp_element_group_160: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_160"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2658_elements(128) & maxPool3D_CP_2658_elements(162);
      gj_maxPool3D_cp_element_group_160 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2658_elements(160), clk => clk, reset => reset); --
    end block;
    -- CP-element group 161:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	80 
    -- CP-element group 161: marked-predecessors 
    -- CP-element group 161: 	163 
    -- CP-element group 161: 	170 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	163 
    -- CP-element group 161:  members (3) 
      -- CP-element group 161: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1759_update_start_
      -- CP-element group 161: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1759_Update/cr
      -- CP-element group 161: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1759_Update/$entry
      -- 
    cr_3421_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3421_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(161), ack => type_cast_1759_inst_req_1); -- 
    maxPool3D_cp_element_group_161: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_161"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool3D_CP_2658_elements(80) & maxPool3D_CP_2658_elements(163) & maxPool3D_CP_2658_elements(170);
      gj_maxPool3D_cp_element_group_161 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2658_elements(161), clk => clk, reset => reset); --
    end block;
    -- CP-element group 162:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	160 
    -- CP-element group 162: successors 
    -- CP-element group 162: marked-successors 
    -- CP-element group 162: 	124 
    -- CP-element group 162: 	160 
    -- CP-element group 162:  members (3) 
      -- CP-element group 162: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1759_sample_completed_
      -- CP-element group 162: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1759_Sample/$exit
      -- CP-element group 162: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1759_Sample/ra
      -- 
    ra_3417_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1759_inst_ack_0, ack => maxPool3D_CP_2658_elements(162)); -- 
    -- CP-element group 163:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	161 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	168 
    -- CP-element group 163: marked-successors 
    -- CP-element group 163: 	102 
    -- CP-element group 163: 	161 
    -- CP-element group 163:  members (3) 
      -- CP-element group 163: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1759_update_completed_
      -- CP-element group 163: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1759_Update/ca
      -- CP-element group 163: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1759_Update/$exit
      -- 
    ca_3422_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1759_inst_ack_1, ack => maxPool3D_CP_2658_elements(163)); -- 
    -- CP-element group 164:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	107 
    -- CP-element group 164: marked-predecessors 
    -- CP-element group 164: 	166 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	166 
    -- CP-element group 164:  members (3) 
      -- CP-element group 164: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/assign_stmt_1763_Sample/req
      -- CP-element group 164: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/assign_stmt_1763_Sample/$entry
      -- CP-element group 164: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/assign_stmt_1763_sample_start_
      -- 
    req_3430_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3430_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(164), ack => W_colx_x1_1751_delayed_1_0_1761_inst_req_0); -- 
    maxPool3D_cp_element_group_164: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_164"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2658_elements(107) & maxPool3D_CP_2658_elements(166);
      gj_maxPool3D_cp_element_group_164 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2658_elements(164), clk => clk, reset => reset); --
    end block;
    -- CP-element group 165:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	80 
    -- CP-element group 165: marked-predecessors 
    -- CP-element group 165: 	167 
    -- CP-element group 165: 	170 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	167 
    -- CP-element group 165:  members (3) 
      -- CP-element group 165: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/assign_stmt_1763_Update/req
      -- CP-element group 165: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/assign_stmt_1763_Update/$entry
      -- CP-element group 165: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/assign_stmt_1763_update_start_
      -- 
    req_3435_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3435_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(165), ack => W_colx_x1_1751_delayed_1_0_1761_inst_req_1); -- 
    maxPool3D_cp_element_group_165: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_165"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool3D_CP_2658_elements(80) & maxPool3D_CP_2658_elements(167) & maxPool3D_CP_2658_elements(170);
      gj_maxPool3D_cp_element_group_165 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2658_elements(165), clk => clk, reset => reset); --
    end block;
    -- CP-element group 166:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	164 
    -- CP-element group 166: successors 
    -- CP-element group 166: marked-successors 
    -- CP-element group 166: 	103 
    -- CP-element group 166: 	164 
    -- CP-element group 166:  members (3) 
      -- CP-element group 166: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/assign_stmt_1763_Sample/ack
      -- CP-element group 166: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/assign_stmt_1763_Sample/$exit
      -- CP-element group 166: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/assign_stmt_1763_sample_completed_
      -- 
    ack_3431_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_colx_x1_1751_delayed_1_0_1761_inst_ack_0, ack => maxPool3D_CP_2658_elements(166)); -- 
    -- CP-element group 167:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	165 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	168 
    -- CP-element group 167: marked-successors 
    -- CP-element group 167: 	102 
    -- CP-element group 167: 	165 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/assign_stmt_1763_Update/ack
      -- CP-element group 167: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/assign_stmt_1763_Update/$exit
      -- CP-element group 167: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/assign_stmt_1763_update_completed_
      -- 
    ack_3436_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_colx_x1_1751_delayed_1_0_1761_inst_ack_1, ack => maxPool3D_CP_2658_elements(167)); -- 
    -- CP-element group 168:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	163 
    -- CP-element group 168: 	167 
    -- CP-element group 168: marked-predecessors 
    -- CP-element group 168: 	170 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	170 
    -- CP-element group 168:  members (3) 
      -- CP-element group 168: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1783_Sample/$entry
      -- CP-element group 168: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1783_Sample/rr
      -- CP-element group 168: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1783_sample_start_
      -- 
    rr_3444_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3444_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(168), ack => type_cast_1783_inst_req_0); -- 
    maxPool3D_cp_element_group_168: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_168"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool3D_CP_2658_elements(163) & maxPool3D_CP_2658_elements(167) & maxPool3D_CP_2658_elements(170);
      gj_maxPool3D_cp_element_group_168 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2658_elements(168), clk => clk, reset => reset); --
    end block;
    -- CP-element group 169:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	80 
    -- CP-element group 169: marked-predecessors 
    -- CP-element group 169: 	171 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	171 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1783_update_start_
      -- CP-element group 169: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1783_Update/cr
      -- CP-element group 169: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1783_Update/$entry
      -- 
    cr_3449_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3449_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(169), ack => type_cast_1783_inst_req_1); -- 
    maxPool3D_cp_element_group_169: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_169"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2658_elements(80) & maxPool3D_CP_2658_elements(171);
      gj_maxPool3D_cp_element_group_169 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2658_elements(169), clk => clk, reset => reset); --
    end block;
    -- CP-element group 170:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	168 
    -- CP-element group 170: successors 
    -- CP-element group 170: marked-successors 
    -- CP-element group 170: 	161 
    -- CP-element group 170: 	165 
    -- CP-element group 170: 	168 
    -- CP-element group 170:  members (3) 
      -- CP-element group 170: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1783_Sample/$exit
      -- CP-element group 170: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1783_sample_completed_
      -- CP-element group 170: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1783_Sample/ra
      -- 
    ra_3445_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1783_inst_ack_0, ack => maxPool3D_CP_2658_elements(170)); -- 
    -- CP-element group 171:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	169 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	78 
    -- CP-element group 171: marked-successors 
    -- CP-element group 171: 	83 
    -- CP-element group 171: 	169 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1783_update_completed_
      -- CP-element group 171: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1783_Update/ca
      -- CP-element group 171: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/type_cast_1783_Update/$exit
      -- 
    ca_3450_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1783_inst_ack_1, ack => maxPool3D_CP_2658_elements(171)); -- 
    -- CP-element group 172:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	86 
    -- CP-element group 172: marked-predecessors 
    -- CP-element group 172: 	174 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	174 
    -- CP-element group 172:  members (3) 
      -- CP-element group 172: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/assign_stmt_1787_Sample/$entry
      -- CP-element group 172: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/assign_stmt_1787_Sample/req
      -- CP-element group 172: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/assign_stmt_1787_sample_start_
      -- 
    req_3458_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3458_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(172), ack => W_rowx_x1_1772_delayed_2_0_1785_inst_req_0); -- 
    maxPool3D_cp_element_group_172: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_172"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2658_elements(86) & maxPool3D_CP_2658_elements(174);
      gj_maxPool3D_cp_element_group_172 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2658_elements(172), clk => clk, reset => reset); --
    end block;
    -- CP-element group 173:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	80 
    -- CP-element group 173: marked-predecessors 
    -- CP-element group 173: 	175 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	175 
    -- CP-element group 173:  members (3) 
      -- CP-element group 173: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/assign_stmt_1787_Update/$entry
      -- CP-element group 173: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/assign_stmt_1787_update_start_
      -- CP-element group 173: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/assign_stmt_1787_Update/req
      -- 
    req_3463_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3463_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(173), ack => W_rowx_x1_1772_delayed_2_0_1785_inst_req_1); -- 
    maxPool3D_cp_element_group_173: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_173"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2658_elements(80) & maxPool3D_CP_2658_elements(175);
      gj_maxPool3D_cp_element_group_173 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2658_elements(173), clk => clk, reset => reset); --
    end block;
    -- CP-element group 174:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	172 
    -- CP-element group 174: successors 
    -- CP-element group 174: marked-successors 
    -- CP-element group 174: 	84 
    -- CP-element group 174: 	172 
    -- CP-element group 174:  members (3) 
      -- CP-element group 174: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/assign_stmt_1787_Sample/$exit
      -- CP-element group 174: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/assign_stmt_1787_sample_completed_
      -- CP-element group 174: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/assign_stmt_1787_Sample/ack
      -- 
    ack_3459_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rowx_x1_1772_delayed_2_0_1785_inst_ack_0, ack => maxPool3D_CP_2658_elements(174)); -- 
    -- CP-element group 175:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	173 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	78 
    -- CP-element group 175: marked-successors 
    -- CP-element group 175: 	83 
    -- CP-element group 175: 	173 
    -- CP-element group 175:  members (3) 
      -- CP-element group 175: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/assign_stmt_1787_update_completed_
      -- CP-element group 175: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/assign_stmt_1787_Update/ack
      -- CP-element group 175: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/assign_stmt_1787_Update/$exit
      -- 
    ack_3464_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rowx_x1_1772_delayed_2_0_1785_inst_ack_1, ack => maxPool3D_CP_2658_elements(175)); -- 
    -- CP-element group 176:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	77 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	78 
    -- CP-element group 176:  members (1) 
      -- CP-element group 176: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group maxPool3D_CP_2658_elements(176) is a control-delay.
    cp_element_176_delay: control_delay_element  generic map(name => " 176_delay", delay_value => 1)  port map(req => maxPool3D_CP_2658_elements(77), ack => maxPool3D_CP_2658_elements(176), clk => clk, reset =>reset);
    -- CP-element group 177:  join  transition  bypass  pipeline-parent 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	80 
    -- CP-element group 177: 	159 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	74 
    -- CP-element group 177:  members (1) 
      -- CP-element group 177: 	 branch_block_stmt_1335/do_while_stmt_1648/do_while_stmt_1648_loop_body/$exit
      -- 
    maxPool3D_cp_element_group_177: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_177"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2658_elements(80) & maxPool3D_CP_2658_elements(159);
      gj_maxPool3D_cp_element_group_177 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2658_elements(177), clk => clk, reset => reset); --
    end block;
    -- CP-element group 178:  transition  input  bypass  pipeline-parent 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	73 
    -- CP-element group 178: successors 
    -- CP-element group 178:  members (2) 
      -- CP-element group 178: 	 branch_block_stmt_1335/do_while_stmt_1648/loop_exit/ack
      -- CP-element group 178: 	 branch_block_stmt_1335/do_while_stmt_1648/loop_exit/$exit
      -- 
    ack_3469_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1648_branch_ack_0, ack => maxPool3D_CP_2658_elements(178)); -- 
    -- CP-element group 179:  transition  input  bypass  pipeline-parent 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	73 
    -- CP-element group 179: successors 
    -- CP-element group 179:  members (2) 
      -- CP-element group 179: 	 branch_block_stmt_1335/do_while_stmt_1648/loop_taken/ack
      -- CP-element group 179: 	 branch_block_stmt_1335/do_while_stmt_1648/loop_taken/$exit
      -- 
    ack_3473_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1648_branch_ack_1, ack => maxPool3D_CP_2658_elements(179)); -- 
    -- CP-element group 180:  transition  bypass  pipeline-parent 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	71 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	1 
    -- CP-element group 180:  members (1) 
      -- CP-element group 180: 	 branch_block_stmt_1335/do_while_stmt_1648/$exit
      -- 
    maxPool3D_CP_2658_elements(180) <= maxPool3D_CP_2658_elements(71);
    -- CP-element group 181:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	1 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	183 
    -- CP-element group 181: 	184 
    -- CP-element group 181:  members (18) 
      -- CP-element group 181: 	 branch_block_stmt_1335/assign_stmt_1821/$entry
      -- CP-element group 181: 	 branch_block_stmt_1335/assign_stmt_1821/type_cast_1820_update_start_
      -- CP-element group 181: 	 branch_block_stmt_1335/assign_stmt_1821__entry__
      -- CP-element group 181: 	 branch_block_stmt_1335/assign_stmt_1821/type_cast_1820_sample_start_
      -- CP-element group 181: 	 branch_block_stmt_1335/merge_stmt_1815__exit__
      -- CP-element group 181: 	 branch_block_stmt_1335/assign_stmt_1821/type_cast_1820_Sample/$entry
      -- CP-element group 181: 	 branch_block_stmt_1335/whilex_xbody_whilex_xend
      -- CP-element group 181: 	 branch_block_stmt_1335/if_stmt_1811_if_link/if_choice_transition
      -- CP-element group 181: 	 branch_block_stmt_1335/if_stmt_1811_if_link/$exit
      -- CP-element group 181: 	 branch_block_stmt_1335/assign_stmt_1821/type_cast_1820_Update/cr
      -- CP-element group 181: 	 branch_block_stmt_1335/assign_stmt_1821/type_cast_1820_Update/$entry
      -- CP-element group 181: 	 branch_block_stmt_1335/assign_stmt_1821/type_cast_1820_Sample/rr
      -- CP-element group 181: 	 branch_block_stmt_1335/whilex_xbody_whilex_xend_PhiReq/$entry
      -- CP-element group 181: 	 branch_block_stmt_1335/whilex_xbody_whilex_xend_PhiReq/$exit
      -- CP-element group 181: 	 branch_block_stmt_1335/merge_stmt_1815_PhiReqMerge
      -- CP-element group 181: 	 branch_block_stmt_1335/merge_stmt_1815_PhiAck/$entry
      -- CP-element group 181: 	 branch_block_stmt_1335/merge_stmt_1815_PhiAck/$exit
      -- CP-element group 181: 	 branch_block_stmt_1335/merge_stmt_1815_PhiAck/dummy
      -- 
    if_choice_transition_3487_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1811_branch_ack_1, ack => maxPool3D_CP_2658_elements(181)); -- 
    cr_3508_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3508_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(181), ack => type_cast_1820_inst_req_1); -- 
    rr_3503_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3503_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(181), ack => type_cast_1820_inst_req_0); -- 
    -- CP-element group 182:  merge  transition  place  input  bypass 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	1 
    -- CP-element group 182: successors 
    -- CP-element group 182:  members (5) 
      -- CP-element group 182: 	 branch_block_stmt_1335/if_stmt_1811__exit__
      -- CP-element group 182: 	 branch_block_stmt_1335/merge_stmt_1815__entry__
      -- CP-element group 182: 	 branch_block_stmt_1335/if_stmt_1811_else_link/else_choice_transition
      -- CP-element group 182: 	 branch_block_stmt_1335/if_stmt_1811_else_link/$exit
      -- CP-element group 182: 	 branch_block_stmt_1335/merge_stmt_1815_dead_link/$entry
      -- 
    else_choice_transition_3491_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1811_branch_ack_0, ack => maxPool3D_CP_2658_elements(182)); -- 
    -- CP-element group 183:  transition  input  bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	181 
    -- CP-element group 183: successors 
    -- CP-element group 183:  members (3) 
      -- CP-element group 183: 	 branch_block_stmt_1335/assign_stmt_1821/type_cast_1820_sample_completed_
      -- CP-element group 183: 	 branch_block_stmt_1335/assign_stmt_1821/type_cast_1820_Sample/ra
      -- CP-element group 183: 	 branch_block_stmt_1335/assign_stmt_1821/type_cast_1820_Sample/$exit
      -- 
    ra_3504_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1820_inst_ack_0, ack => maxPool3D_CP_2658_elements(183)); -- 
    -- CP-element group 184:  fork  transition  place  input  output  bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	181 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	185 
    -- CP-element group 184: 	186 
    -- CP-element group 184: 	188 
    -- CP-element group 184: 	190 
    -- CP-element group 184: 	192 
    -- CP-element group 184: 	194 
    -- CP-element group 184: 	196 
    -- CP-element group 184: 	198 
    -- CP-element group 184: 	200 
    -- CP-element group 184: 	202 
    -- CP-element group 184: 	204 
    -- CP-element group 184:  members (40) 
      -- CP-element group 184: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935__entry__
      -- CP-element group 184: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1828_update_start_
      -- CP-element group 184: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/call_stmt_1824_sample_start_
      -- CP-element group 184: 	 branch_block_stmt_1335/assign_stmt_1821__exit__
      -- CP-element group 184: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/call_stmt_1824_Sample/crr
      -- CP-element group 184: 	 branch_block_stmt_1335/assign_stmt_1821/$exit
      -- CP-element group 184: 	 branch_block_stmt_1335/assign_stmt_1821/type_cast_1820_update_completed_
      -- CP-element group 184: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/$entry
      -- CP-element group 184: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1847_update_start_
      -- CP-element group 184: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/call_stmt_1824_Sample/$entry
      -- CP-element group 184: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/call_stmt_1824_Update/ccr
      -- CP-element group 184: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/call_stmt_1824_update_start_
      -- CP-element group 184: 	 branch_block_stmt_1335/assign_stmt_1821/type_cast_1820_Update/ca
      -- CP-element group 184: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1837_Update/cr
      -- CP-element group 184: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/call_stmt_1824_Update/$entry
      -- CP-element group 184: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1837_Update/$entry
      -- CP-element group 184: 	 branch_block_stmt_1335/assign_stmt_1821/type_cast_1820_Update/$exit
      -- CP-element group 184: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1828_Update/cr
      -- CP-element group 184: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1837_update_start_
      -- CP-element group 184: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1828_Update/$entry
      -- CP-element group 184: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1847_Update/$entry
      -- CP-element group 184: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1847_Update/cr
      -- CP-element group 184: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1857_update_start_
      -- CP-element group 184: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1857_Update/$entry
      -- CP-element group 184: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1857_Update/cr
      -- CP-element group 184: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1867_update_start_
      -- CP-element group 184: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1867_Update/$entry
      -- CP-element group 184: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1867_Update/cr
      -- CP-element group 184: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1877_update_start_
      -- CP-element group 184: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1877_Update/$entry
      -- CP-element group 184: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1877_Update/cr
      -- CP-element group 184: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1887_update_start_
      -- CP-element group 184: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1887_Update/$entry
      -- CP-element group 184: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1887_Update/cr
      -- CP-element group 184: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1897_update_start_
      -- CP-element group 184: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1897_Update/$entry
      -- CP-element group 184: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1897_Update/cr
      -- CP-element group 184: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1907_update_start_
      -- CP-element group 184: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1907_Update/$entry
      -- CP-element group 184: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1907_Update/cr
      -- 
    ca_3509_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1820_inst_ack_1, ack => maxPool3D_CP_2658_elements(184)); -- 
    crr_3520_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3520_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(184), ack => call_stmt_1824_call_req_0); -- 
    ccr_3525_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3525_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(184), ack => call_stmt_1824_call_req_1); -- 
    cr_3553_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3553_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(184), ack => type_cast_1837_inst_req_1); -- 
    cr_3539_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3539_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(184), ack => type_cast_1828_inst_req_1); -- 
    cr_3567_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3567_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(184), ack => type_cast_1847_inst_req_1); -- 
    cr_3581_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3581_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(184), ack => type_cast_1857_inst_req_1); -- 
    cr_3595_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3595_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(184), ack => type_cast_1867_inst_req_1); -- 
    cr_3609_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3609_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(184), ack => type_cast_1877_inst_req_1); -- 
    cr_3623_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3623_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(184), ack => type_cast_1887_inst_req_1); -- 
    cr_3637_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3637_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(184), ack => type_cast_1897_inst_req_1); -- 
    cr_3651_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3651_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(184), ack => type_cast_1907_inst_req_1); -- 
    -- CP-element group 185:  transition  input  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	184 
    -- CP-element group 185: successors 
    -- CP-element group 185:  members (3) 
      -- CP-element group 185: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/call_stmt_1824_Sample/$exit
      -- CP-element group 185: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/call_stmt_1824_sample_completed_
      -- CP-element group 185: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/call_stmt_1824_Sample/cra
      -- 
    cra_3521_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1824_call_ack_0, ack => maxPool3D_CP_2658_elements(185)); -- 
    -- CP-element group 186:  transition  input  output  bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	184 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	187 
    -- CP-element group 186:  members (6) 
      -- CP-element group 186: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1828_sample_start_
      -- CP-element group 186: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/call_stmt_1824_update_completed_
      -- CP-element group 186: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1828_Sample/rr
      -- CP-element group 186: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1828_Sample/$entry
      -- CP-element group 186: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/call_stmt_1824_Update/cca
      -- CP-element group 186: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/call_stmt_1824_Update/$exit
      -- 
    cca_3526_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1824_call_ack_1, ack => maxPool3D_CP_2658_elements(186)); -- 
    rr_3534_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3534_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(186), ack => type_cast_1828_inst_req_0); -- 
    -- CP-element group 187:  transition  input  bypass 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	186 
    -- CP-element group 187: successors 
    -- CP-element group 187:  members (3) 
      -- CP-element group 187: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1828_sample_completed_
      -- CP-element group 187: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1828_Sample/ra
      -- CP-element group 187: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1828_Sample/$exit
      -- 
    ra_3535_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1828_inst_ack_0, ack => maxPool3D_CP_2658_elements(187)); -- 
    -- CP-element group 188:  fork  transition  input  output  bypass 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	184 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	189 
    -- CP-element group 188: 	191 
    -- CP-element group 188: 	193 
    -- CP-element group 188: 	195 
    -- CP-element group 188: 	197 
    -- CP-element group 188: 	199 
    -- CP-element group 188: 	201 
    -- CP-element group 188: 	203 
    -- CP-element group 188: 	228 
    -- CP-element group 188:  members (30) 
      -- CP-element group 188: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1837_sample_start_
      -- CP-element group 188: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1847_sample_start_
      -- CP-element group 188: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1837_Sample/rr
      -- CP-element group 188: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1837_Sample/$entry
      -- CP-element group 188: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1828_update_completed_
      -- CP-element group 188: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1828_Update/ca
      -- CP-element group 188: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1828_Update/$exit
      -- CP-element group 188: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1847_Sample/$entry
      -- CP-element group 188: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1847_Sample/rr
      -- CP-element group 188: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1857_sample_start_
      -- CP-element group 188: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1857_Sample/$entry
      -- CP-element group 188: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1857_Sample/rr
      -- CP-element group 188: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1867_sample_start_
      -- CP-element group 188: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1867_Sample/$entry
      -- CP-element group 188: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1867_Sample/rr
      -- CP-element group 188: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1877_sample_start_
      -- CP-element group 188: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1877_Sample/$entry
      -- CP-element group 188: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1877_Sample/rr
      -- CP-element group 188: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1887_sample_start_
      -- CP-element group 188: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1887_Sample/$entry
      -- CP-element group 188: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1887_Sample/rr
      -- CP-element group 188: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1897_sample_start_
      -- CP-element group 188: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1897_Sample/$entry
      -- CP-element group 188: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1897_Sample/rr
      -- CP-element group 188: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1907_sample_start_
      -- CP-element group 188: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1907_Sample/$entry
      -- CP-element group 188: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1907_Sample/rr
      -- CP-element group 188: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_elapsed_time_pipe_1933_sample_start_
      -- CP-element group 188: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_elapsed_time_pipe_1933_Sample/$entry
      -- CP-element group 188: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_elapsed_time_pipe_1933_Sample/req
      -- 
    ca_3540_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1828_inst_ack_1, ack => maxPool3D_CP_2658_elements(188)); -- 
    rr_3548_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3548_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(188), ack => type_cast_1837_inst_req_0); -- 
    rr_3562_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3562_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(188), ack => type_cast_1847_inst_req_0); -- 
    rr_3576_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3576_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(188), ack => type_cast_1857_inst_req_0); -- 
    rr_3590_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3590_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(188), ack => type_cast_1867_inst_req_0); -- 
    rr_3604_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3604_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(188), ack => type_cast_1877_inst_req_0); -- 
    rr_3618_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3618_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(188), ack => type_cast_1887_inst_req_0); -- 
    rr_3632_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3632_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(188), ack => type_cast_1897_inst_req_0); -- 
    rr_3646_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3646_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(188), ack => type_cast_1907_inst_req_0); -- 
    req_3772_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3772_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(188), ack => WPIPE_elapsed_time_pipe_1933_inst_req_0); -- 
    -- CP-element group 189:  transition  input  bypass 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	188 
    -- CP-element group 189: successors 
    -- CP-element group 189:  members (3) 
      -- CP-element group 189: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1837_Sample/ra
      -- CP-element group 189: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1837_Sample/$exit
      -- CP-element group 189: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1837_sample_completed_
      -- 
    ra_3549_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1837_inst_ack_0, ack => maxPool3D_CP_2658_elements(189)); -- 
    -- CP-element group 190:  transition  input  bypass 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	184 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	225 
    -- CP-element group 190:  members (3) 
      -- CP-element group 190: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1837_Update/ca
      -- CP-element group 190: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1837_update_completed_
      -- CP-element group 190: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1837_Update/$exit
      -- 
    ca_3554_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1837_inst_ack_1, ack => maxPool3D_CP_2658_elements(190)); -- 
    -- CP-element group 191:  transition  input  bypass 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	188 
    -- CP-element group 191: successors 
    -- CP-element group 191:  members (3) 
      -- CP-element group 191: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1847_sample_completed_
      -- CP-element group 191: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1847_Sample/$exit
      -- CP-element group 191: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1847_Sample/ra
      -- 
    ra_3563_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1847_inst_ack_0, ack => maxPool3D_CP_2658_elements(191)); -- 
    -- CP-element group 192:  transition  input  bypass 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	184 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	222 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1847_update_completed_
      -- CP-element group 192: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1847_Update/$exit
      -- CP-element group 192: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1847_Update/ca
      -- 
    ca_3568_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1847_inst_ack_1, ack => maxPool3D_CP_2658_elements(192)); -- 
    -- CP-element group 193:  transition  input  bypass 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	188 
    -- CP-element group 193: successors 
    -- CP-element group 193:  members (3) 
      -- CP-element group 193: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1857_sample_completed_
      -- CP-element group 193: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1857_Sample/$exit
      -- CP-element group 193: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1857_Sample/ra
      -- 
    ra_3577_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1857_inst_ack_0, ack => maxPool3D_CP_2658_elements(193)); -- 
    -- CP-element group 194:  transition  input  bypass 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	184 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	219 
    -- CP-element group 194:  members (3) 
      -- CP-element group 194: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1857_update_completed_
      -- CP-element group 194: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1857_Update/$exit
      -- CP-element group 194: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1857_Update/ca
      -- 
    ca_3582_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1857_inst_ack_1, ack => maxPool3D_CP_2658_elements(194)); -- 
    -- CP-element group 195:  transition  input  bypass 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	188 
    -- CP-element group 195: successors 
    -- CP-element group 195:  members (3) 
      -- CP-element group 195: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1867_sample_completed_
      -- CP-element group 195: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1867_Sample/$exit
      -- CP-element group 195: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1867_Sample/ra
      -- 
    ra_3591_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1867_inst_ack_0, ack => maxPool3D_CP_2658_elements(195)); -- 
    -- CP-element group 196:  transition  input  bypass 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	184 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	216 
    -- CP-element group 196:  members (3) 
      -- CP-element group 196: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1867_update_completed_
      -- CP-element group 196: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1867_Update/$exit
      -- CP-element group 196: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1867_Update/ca
      -- 
    ca_3596_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1867_inst_ack_1, ack => maxPool3D_CP_2658_elements(196)); -- 
    -- CP-element group 197:  transition  input  bypass 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	188 
    -- CP-element group 197: successors 
    -- CP-element group 197:  members (3) 
      -- CP-element group 197: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1877_sample_completed_
      -- CP-element group 197: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1877_Sample/$exit
      -- CP-element group 197: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1877_Sample/ra
      -- 
    ra_3605_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1877_inst_ack_0, ack => maxPool3D_CP_2658_elements(197)); -- 
    -- CP-element group 198:  transition  input  bypass 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	184 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	213 
    -- CP-element group 198:  members (3) 
      -- CP-element group 198: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1877_update_completed_
      -- CP-element group 198: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1877_Update/$exit
      -- CP-element group 198: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1877_Update/ca
      -- 
    ca_3610_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1877_inst_ack_1, ack => maxPool3D_CP_2658_elements(198)); -- 
    -- CP-element group 199:  transition  input  bypass 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	188 
    -- CP-element group 199: successors 
    -- CP-element group 199:  members (3) 
      -- CP-element group 199: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1887_sample_completed_
      -- CP-element group 199: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1887_Sample/$exit
      -- CP-element group 199: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1887_Sample/ra
      -- 
    ra_3619_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1887_inst_ack_0, ack => maxPool3D_CP_2658_elements(199)); -- 
    -- CP-element group 200:  transition  input  bypass 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	184 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	210 
    -- CP-element group 200:  members (3) 
      -- CP-element group 200: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1887_update_completed_
      -- CP-element group 200: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1887_Update/$exit
      -- CP-element group 200: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1887_Update/ca
      -- 
    ca_3624_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 200_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1887_inst_ack_1, ack => maxPool3D_CP_2658_elements(200)); -- 
    -- CP-element group 201:  transition  input  bypass 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	188 
    -- CP-element group 201: successors 
    -- CP-element group 201:  members (3) 
      -- CP-element group 201: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1897_sample_completed_
      -- CP-element group 201: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1897_Sample/$exit
      -- CP-element group 201: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1897_Sample/ra
      -- 
    ra_3633_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1897_inst_ack_0, ack => maxPool3D_CP_2658_elements(201)); -- 
    -- CP-element group 202:  transition  input  bypass 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	184 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	207 
    -- CP-element group 202:  members (3) 
      -- CP-element group 202: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1897_update_completed_
      -- CP-element group 202: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1897_Update/$exit
      -- CP-element group 202: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1897_Update/ca
      -- 
    ca_3638_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1897_inst_ack_1, ack => maxPool3D_CP_2658_elements(202)); -- 
    -- CP-element group 203:  transition  input  bypass 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	188 
    -- CP-element group 203: successors 
    -- CP-element group 203:  members (3) 
      -- CP-element group 203: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1907_sample_completed_
      -- CP-element group 203: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1907_Sample/$exit
      -- CP-element group 203: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1907_Sample/ra
      -- 
    ra_3647_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 203_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1907_inst_ack_0, ack => maxPool3D_CP_2658_elements(203)); -- 
    -- CP-element group 204:  transition  input  output  bypass 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	184 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	205 
    -- CP-element group 204:  members (6) 
      -- CP-element group 204: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1907_update_completed_
      -- CP-element group 204: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1907_Update/$exit
      -- CP-element group 204: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/type_cast_1907_Update/ca
      -- CP-element group 204: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1909_sample_start_
      -- CP-element group 204: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1909_Sample/$entry
      -- CP-element group 204: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1909_Sample/req
      -- 
    ca_3652_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 204_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1907_inst_ack_1, ack => maxPool3D_CP_2658_elements(204)); -- 
    req_3660_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3660_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(204), ack => WPIPE_maxpool_output_pipe_1909_inst_req_0); -- 
    -- CP-element group 205:  transition  input  output  bypass 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	204 
    -- CP-element group 205: successors 
    -- CP-element group 205: 	206 
    -- CP-element group 205:  members (6) 
      -- CP-element group 205: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1909_sample_completed_
      -- CP-element group 205: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1909_update_start_
      -- CP-element group 205: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1909_Sample/$exit
      -- CP-element group 205: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1909_Sample/ack
      -- CP-element group 205: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1909_Update/$entry
      -- CP-element group 205: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1909_Update/req
      -- 
    ack_3661_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1909_inst_ack_0, ack => maxPool3D_CP_2658_elements(205)); -- 
    req_3665_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3665_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(205), ack => WPIPE_maxpool_output_pipe_1909_inst_req_1); -- 
    -- CP-element group 206:  transition  input  bypass 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	205 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	207 
    -- CP-element group 206:  members (3) 
      -- CP-element group 206: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1909_update_completed_
      -- CP-element group 206: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1909_Update/$exit
      -- CP-element group 206: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1909_Update/ack
      -- 
    ack_3666_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 206_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1909_inst_ack_1, ack => maxPool3D_CP_2658_elements(206)); -- 
    -- CP-element group 207:  join  transition  output  bypass 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	202 
    -- CP-element group 207: 	206 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	208 
    -- CP-element group 207:  members (3) 
      -- CP-element group 207: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1912_sample_start_
      -- CP-element group 207: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1912_Sample/$entry
      -- CP-element group 207: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1912_Sample/req
      -- 
    req_3674_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3674_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(207), ack => WPIPE_maxpool_output_pipe_1912_inst_req_0); -- 
    maxPool3D_cp_element_group_207: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_207"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2658_elements(202) & maxPool3D_CP_2658_elements(206);
      gj_maxPool3D_cp_element_group_207 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2658_elements(207), clk => clk, reset => reset); --
    end block;
    -- CP-element group 208:  transition  input  output  bypass 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	207 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	209 
    -- CP-element group 208:  members (6) 
      -- CP-element group 208: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1912_sample_completed_
      -- CP-element group 208: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1912_update_start_
      -- CP-element group 208: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1912_Sample/$exit
      -- CP-element group 208: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1912_Sample/ack
      -- CP-element group 208: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1912_Update/$entry
      -- CP-element group 208: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1912_Update/req
      -- 
    ack_3675_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 208_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1912_inst_ack_0, ack => maxPool3D_CP_2658_elements(208)); -- 
    req_3679_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3679_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(208), ack => WPIPE_maxpool_output_pipe_1912_inst_req_1); -- 
    -- CP-element group 209:  transition  input  bypass 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	208 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	210 
    -- CP-element group 209:  members (3) 
      -- CP-element group 209: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1912_update_completed_
      -- CP-element group 209: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1912_Update/$exit
      -- CP-element group 209: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1912_Update/ack
      -- 
    ack_3680_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1912_inst_ack_1, ack => maxPool3D_CP_2658_elements(209)); -- 
    -- CP-element group 210:  join  transition  output  bypass 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	200 
    -- CP-element group 210: 	209 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	211 
    -- CP-element group 210:  members (3) 
      -- CP-element group 210: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1915_sample_start_
      -- CP-element group 210: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1915_Sample/$entry
      -- CP-element group 210: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1915_Sample/req
      -- 
    req_3688_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3688_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(210), ack => WPIPE_maxpool_output_pipe_1915_inst_req_0); -- 
    maxPool3D_cp_element_group_210: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_210"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2658_elements(200) & maxPool3D_CP_2658_elements(209);
      gj_maxPool3D_cp_element_group_210 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2658_elements(210), clk => clk, reset => reset); --
    end block;
    -- CP-element group 211:  transition  input  output  bypass 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	210 
    -- CP-element group 211: successors 
    -- CP-element group 211: 	212 
    -- CP-element group 211:  members (6) 
      -- CP-element group 211: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1915_sample_completed_
      -- CP-element group 211: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1915_update_start_
      -- CP-element group 211: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1915_Sample/$exit
      -- CP-element group 211: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1915_Sample/ack
      -- CP-element group 211: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1915_Update/$entry
      -- CP-element group 211: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1915_Update/req
      -- 
    ack_3689_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 211_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1915_inst_ack_0, ack => maxPool3D_CP_2658_elements(211)); -- 
    req_3693_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3693_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(211), ack => WPIPE_maxpool_output_pipe_1915_inst_req_1); -- 
    -- CP-element group 212:  transition  input  bypass 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	211 
    -- CP-element group 212: successors 
    -- CP-element group 212: 	213 
    -- CP-element group 212:  members (3) 
      -- CP-element group 212: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1915_update_completed_
      -- CP-element group 212: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1915_Update/$exit
      -- CP-element group 212: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1915_Update/ack
      -- 
    ack_3694_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 212_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1915_inst_ack_1, ack => maxPool3D_CP_2658_elements(212)); -- 
    -- CP-element group 213:  join  transition  output  bypass 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	198 
    -- CP-element group 213: 	212 
    -- CP-element group 213: successors 
    -- CP-element group 213: 	214 
    -- CP-element group 213:  members (3) 
      -- CP-element group 213: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1918_sample_start_
      -- CP-element group 213: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1918_Sample/$entry
      -- CP-element group 213: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1918_Sample/req
      -- 
    req_3702_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3702_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(213), ack => WPIPE_maxpool_output_pipe_1918_inst_req_0); -- 
    maxPool3D_cp_element_group_213: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_213"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2658_elements(198) & maxPool3D_CP_2658_elements(212);
      gj_maxPool3D_cp_element_group_213 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2658_elements(213), clk => clk, reset => reset); --
    end block;
    -- CP-element group 214:  transition  input  output  bypass 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	213 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	215 
    -- CP-element group 214:  members (6) 
      -- CP-element group 214: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1918_sample_completed_
      -- CP-element group 214: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1918_update_start_
      -- CP-element group 214: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1918_Sample/$exit
      -- CP-element group 214: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1918_Sample/ack
      -- CP-element group 214: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1918_Update/$entry
      -- CP-element group 214: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1918_Update/req
      -- 
    ack_3703_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 214_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1918_inst_ack_0, ack => maxPool3D_CP_2658_elements(214)); -- 
    req_3707_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3707_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(214), ack => WPIPE_maxpool_output_pipe_1918_inst_req_1); -- 
    -- CP-element group 215:  transition  input  bypass 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	214 
    -- CP-element group 215: successors 
    -- CP-element group 215: 	216 
    -- CP-element group 215:  members (3) 
      -- CP-element group 215: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1918_update_completed_
      -- CP-element group 215: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1918_Update/$exit
      -- CP-element group 215: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1918_Update/ack
      -- 
    ack_3708_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 215_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1918_inst_ack_1, ack => maxPool3D_CP_2658_elements(215)); -- 
    -- CP-element group 216:  join  transition  output  bypass 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	196 
    -- CP-element group 216: 	215 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	217 
    -- CP-element group 216:  members (3) 
      -- CP-element group 216: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1921_sample_start_
      -- CP-element group 216: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1921_Sample/$entry
      -- CP-element group 216: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1921_Sample/req
      -- 
    req_3716_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3716_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(216), ack => WPIPE_maxpool_output_pipe_1921_inst_req_0); -- 
    maxPool3D_cp_element_group_216: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_216"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2658_elements(196) & maxPool3D_CP_2658_elements(215);
      gj_maxPool3D_cp_element_group_216 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2658_elements(216), clk => clk, reset => reset); --
    end block;
    -- CP-element group 217:  transition  input  output  bypass 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	216 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	218 
    -- CP-element group 217:  members (6) 
      -- CP-element group 217: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1921_sample_completed_
      -- CP-element group 217: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1921_update_start_
      -- CP-element group 217: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1921_Sample/$exit
      -- CP-element group 217: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1921_Sample/ack
      -- CP-element group 217: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1921_Update/$entry
      -- CP-element group 217: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1921_Update/req
      -- 
    ack_3717_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 217_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1921_inst_ack_0, ack => maxPool3D_CP_2658_elements(217)); -- 
    req_3721_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3721_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(217), ack => WPIPE_maxpool_output_pipe_1921_inst_req_1); -- 
    -- CP-element group 218:  transition  input  bypass 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	217 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	219 
    -- CP-element group 218:  members (3) 
      -- CP-element group 218: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1921_update_completed_
      -- CP-element group 218: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1921_Update/$exit
      -- CP-element group 218: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1921_Update/ack
      -- 
    ack_3722_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 218_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1921_inst_ack_1, ack => maxPool3D_CP_2658_elements(218)); -- 
    -- CP-element group 219:  join  transition  output  bypass 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	194 
    -- CP-element group 219: 	218 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	220 
    -- CP-element group 219:  members (3) 
      -- CP-element group 219: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1924_sample_start_
      -- CP-element group 219: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1924_Sample/$entry
      -- CP-element group 219: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1924_Sample/req
      -- 
    req_3730_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3730_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(219), ack => WPIPE_maxpool_output_pipe_1924_inst_req_0); -- 
    maxPool3D_cp_element_group_219: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_219"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2658_elements(194) & maxPool3D_CP_2658_elements(218);
      gj_maxPool3D_cp_element_group_219 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2658_elements(219), clk => clk, reset => reset); --
    end block;
    -- CP-element group 220:  transition  input  output  bypass 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	219 
    -- CP-element group 220: successors 
    -- CP-element group 220: 	221 
    -- CP-element group 220:  members (6) 
      -- CP-element group 220: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1924_sample_completed_
      -- CP-element group 220: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1924_update_start_
      -- CP-element group 220: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1924_Sample/$exit
      -- CP-element group 220: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1924_Sample/ack
      -- CP-element group 220: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1924_Update/$entry
      -- CP-element group 220: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1924_Update/req
      -- 
    ack_3731_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1924_inst_ack_0, ack => maxPool3D_CP_2658_elements(220)); -- 
    req_3735_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3735_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(220), ack => WPIPE_maxpool_output_pipe_1924_inst_req_1); -- 
    -- CP-element group 221:  transition  input  bypass 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	220 
    -- CP-element group 221: successors 
    -- CP-element group 221: 	222 
    -- CP-element group 221:  members (3) 
      -- CP-element group 221: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1924_update_completed_
      -- CP-element group 221: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1924_Update/$exit
      -- CP-element group 221: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1924_Update/ack
      -- 
    ack_3736_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1924_inst_ack_1, ack => maxPool3D_CP_2658_elements(221)); -- 
    -- CP-element group 222:  join  transition  output  bypass 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	192 
    -- CP-element group 222: 	221 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	223 
    -- CP-element group 222:  members (3) 
      -- CP-element group 222: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1927_sample_start_
      -- CP-element group 222: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1927_Sample/$entry
      -- CP-element group 222: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1927_Sample/req
      -- 
    req_3744_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3744_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(222), ack => WPIPE_maxpool_output_pipe_1927_inst_req_0); -- 
    maxPool3D_cp_element_group_222: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_222"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2658_elements(192) & maxPool3D_CP_2658_elements(221);
      gj_maxPool3D_cp_element_group_222 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2658_elements(222), clk => clk, reset => reset); --
    end block;
    -- CP-element group 223:  transition  input  output  bypass 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	222 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	224 
    -- CP-element group 223:  members (6) 
      -- CP-element group 223: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1927_sample_completed_
      -- CP-element group 223: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1927_update_start_
      -- CP-element group 223: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1927_Sample/$exit
      -- CP-element group 223: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1927_Sample/ack
      -- CP-element group 223: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1927_Update/$entry
      -- CP-element group 223: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1927_Update/req
      -- 
    ack_3745_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 223_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1927_inst_ack_0, ack => maxPool3D_CP_2658_elements(223)); -- 
    req_3749_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3749_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(223), ack => WPIPE_maxpool_output_pipe_1927_inst_req_1); -- 
    -- CP-element group 224:  transition  input  bypass 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	223 
    -- CP-element group 224: successors 
    -- CP-element group 224: 	225 
    -- CP-element group 224:  members (3) 
      -- CP-element group 224: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1927_update_completed_
      -- CP-element group 224: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1927_Update/$exit
      -- CP-element group 224: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1927_Update/ack
      -- 
    ack_3750_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1927_inst_ack_1, ack => maxPool3D_CP_2658_elements(224)); -- 
    -- CP-element group 225:  join  transition  output  bypass 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	190 
    -- CP-element group 225: 	224 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	226 
    -- CP-element group 225:  members (3) 
      -- CP-element group 225: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1930_sample_start_
      -- CP-element group 225: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1930_Sample/$entry
      -- CP-element group 225: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1930_Sample/req
      -- 
    req_3758_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3758_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(225), ack => WPIPE_maxpool_output_pipe_1930_inst_req_0); -- 
    maxPool3D_cp_element_group_225: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_225"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2658_elements(190) & maxPool3D_CP_2658_elements(224);
      gj_maxPool3D_cp_element_group_225 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2658_elements(225), clk => clk, reset => reset); --
    end block;
    -- CP-element group 226:  transition  input  output  bypass 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	225 
    -- CP-element group 226: successors 
    -- CP-element group 226: 	227 
    -- CP-element group 226:  members (6) 
      -- CP-element group 226: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1930_sample_completed_
      -- CP-element group 226: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1930_update_start_
      -- CP-element group 226: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1930_Sample/$exit
      -- CP-element group 226: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1930_Sample/ack
      -- CP-element group 226: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1930_Update/$entry
      -- CP-element group 226: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1930_Update/req
      -- 
    ack_3759_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 226_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1930_inst_ack_0, ack => maxPool3D_CP_2658_elements(226)); -- 
    req_3763_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3763_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(226), ack => WPIPE_maxpool_output_pipe_1930_inst_req_1); -- 
    -- CP-element group 227:  transition  input  bypass 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	226 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	230 
    -- CP-element group 227:  members (3) 
      -- CP-element group 227: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1930_update_completed_
      -- CP-element group 227: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1930_Update/$exit
      -- CP-element group 227: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_maxpool_output_pipe_1930_Update/ack
      -- 
    ack_3764_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 227_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1930_inst_ack_1, ack => maxPool3D_CP_2658_elements(227)); -- 
    -- CP-element group 228:  transition  input  output  bypass 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	188 
    -- CP-element group 228: successors 
    -- CP-element group 228: 	229 
    -- CP-element group 228:  members (6) 
      -- CP-element group 228: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_elapsed_time_pipe_1933_sample_completed_
      -- CP-element group 228: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_elapsed_time_pipe_1933_update_start_
      -- CP-element group 228: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_elapsed_time_pipe_1933_Sample/$exit
      -- CP-element group 228: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_elapsed_time_pipe_1933_Sample/ack
      -- CP-element group 228: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_elapsed_time_pipe_1933_Update/$entry
      -- CP-element group 228: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_elapsed_time_pipe_1933_Update/req
      -- 
    ack_3773_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 228_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_elapsed_time_pipe_1933_inst_ack_0, ack => maxPool3D_CP_2658_elements(228)); -- 
    req_3777_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3777_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(228), ack => WPIPE_elapsed_time_pipe_1933_inst_req_1); -- 
    -- CP-element group 229:  transition  input  bypass 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	228 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	230 
    -- CP-element group 229:  members (3) 
      -- CP-element group 229: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_elapsed_time_pipe_1933_update_completed_
      -- CP-element group 229: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_elapsed_time_pipe_1933_Update/$exit
      -- CP-element group 229: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/WPIPE_elapsed_time_pipe_1933_Update/ack
      -- 
    ack_3778_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 229_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_elapsed_time_pipe_1933_inst_ack_1, ack => maxPool3D_CP_2658_elements(229)); -- 
    -- CP-element group 230:  join  fork  transition  place  output  bypass 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	227 
    -- CP-element group 230: 	229 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	231 
    -- CP-element group 230: 	232 
    -- CP-element group 230: 	233 
    -- CP-element group 230: 	234 
    -- CP-element group 230: 	237 
    -- CP-element group 230:  members (19) 
      -- CP-element group 230: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935__exit__
      -- CP-element group 230: 	 branch_block_stmt_1335/assign_stmt_1940_to_call_stmt_1956__entry__
      -- CP-element group 230: 	 branch_block_stmt_1335/call_stmt_1824_to_assign_stmt_1935/$exit
      -- CP-element group 230: 	 branch_block_stmt_1335/assign_stmt_1940_to_call_stmt_1956/$entry
      -- CP-element group 230: 	 branch_block_stmt_1335/assign_stmt_1940_to_call_stmt_1956/type_cast_1939_sample_start_
      -- CP-element group 230: 	 branch_block_stmt_1335/assign_stmt_1940_to_call_stmt_1956/type_cast_1939_update_start_
      -- CP-element group 230: 	 branch_block_stmt_1335/assign_stmt_1940_to_call_stmt_1956/type_cast_1939_Sample/$entry
      -- CP-element group 230: 	 branch_block_stmt_1335/assign_stmt_1940_to_call_stmt_1956/type_cast_1939_Sample/rr
      -- CP-element group 230: 	 branch_block_stmt_1335/assign_stmt_1940_to_call_stmt_1956/type_cast_1939_Update/$entry
      -- CP-element group 230: 	 branch_block_stmt_1335/assign_stmt_1940_to_call_stmt_1956/type_cast_1939_Update/cr
      -- CP-element group 230: 	 branch_block_stmt_1335/assign_stmt_1940_to_call_stmt_1956/type_cast_1943_sample_start_
      -- CP-element group 230: 	 branch_block_stmt_1335/assign_stmt_1940_to_call_stmt_1956/type_cast_1943_update_start_
      -- CP-element group 230: 	 branch_block_stmt_1335/assign_stmt_1940_to_call_stmt_1956/type_cast_1943_Sample/$entry
      -- CP-element group 230: 	 branch_block_stmt_1335/assign_stmt_1940_to_call_stmt_1956/type_cast_1943_Sample/rr
      -- CP-element group 230: 	 branch_block_stmt_1335/assign_stmt_1940_to_call_stmt_1956/type_cast_1943_Update/$entry
      -- CP-element group 230: 	 branch_block_stmt_1335/assign_stmt_1940_to_call_stmt_1956/type_cast_1943_Update/cr
      -- CP-element group 230: 	 branch_block_stmt_1335/assign_stmt_1940_to_call_stmt_1956/call_stmt_1956_update_start_
      -- CP-element group 230: 	 branch_block_stmt_1335/assign_stmt_1940_to_call_stmt_1956/call_stmt_1956_Update/$entry
      -- CP-element group 230: 	 branch_block_stmt_1335/assign_stmt_1940_to_call_stmt_1956/call_stmt_1956_Update/ccr
      -- 
    rr_3789_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3789_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(230), ack => type_cast_1939_inst_req_0); -- 
    cr_3794_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3794_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(230), ack => type_cast_1939_inst_req_1); -- 
    rr_3803_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3803_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(230), ack => type_cast_1943_inst_req_0); -- 
    cr_3808_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3808_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(230), ack => type_cast_1943_inst_req_1); -- 
    ccr_3822_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3822_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(230), ack => call_stmt_1956_call_req_1); -- 
    maxPool3D_cp_element_group_230: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_230"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2658_elements(227) & maxPool3D_CP_2658_elements(229);
      gj_maxPool3D_cp_element_group_230 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2658_elements(230), clk => clk, reset => reset); --
    end block;
    -- CP-element group 231:  transition  input  bypass 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	230 
    -- CP-element group 231: successors 
    -- CP-element group 231:  members (3) 
      -- CP-element group 231: 	 branch_block_stmt_1335/assign_stmt_1940_to_call_stmt_1956/type_cast_1939_sample_completed_
      -- CP-element group 231: 	 branch_block_stmt_1335/assign_stmt_1940_to_call_stmt_1956/type_cast_1939_Sample/$exit
      -- CP-element group 231: 	 branch_block_stmt_1335/assign_stmt_1940_to_call_stmt_1956/type_cast_1939_Sample/ra
      -- 
    ra_3790_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 231_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1939_inst_ack_0, ack => maxPool3D_CP_2658_elements(231)); -- 
    -- CP-element group 232:  transition  input  bypass 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	230 
    -- CP-element group 232: successors 
    -- CP-element group 232: 	235 
    -- CP-element group 232:  members (3) 
      -- CP-element group 232: 	 branch_block_stmt_1335/assign_stmt_1940_to_call_stmt_1956/type_cast_1939_update_completed_
      -- CP-element group 232: 	 branch_block_stmt_1335/assign_stmt_1940_to_call_stmt_1956/type_cast_1939_Update/$exit
      -- CP-element group 232: 	 branch_block_stmt_1335/assign_stmt_1940_to_call_stmt_1956/type_cast_1939_Update/ca
      -- 
    ca_3795_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 232_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1939_inst_ack_1, ack => maxPool3D_CP_2658_elements(232)); -- 
    -- CP-element group 233:  transition  input  bypass 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	230 
    -- CP-element group 233: successors 
    -- CP-element group 233:  members (3) 
      -- CP-element group 233: 	 branch_block_stmt_1335/assign_stmt_1940_to_call_stmt_1956/type_cast_1943_sample_completed_
      -- CP-element group 233: 	 branch_block_stmt_1335/assign_stmt_1940_to_call_stmt_1956/type_cast_1943_Sample/$exit
      -- CP-element group 233: 	 branch_block_stmt_1335/assign_stmt_1940_to_call_stmt_1956/type_cast_1943_Sample/ra
      -- 
    ra_3804_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 233_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1943_inst_ack_0, ack => maxPool3D_CP_2658_elements(233)); -- 
    -- CP-element group 234:  transition  input  bypass 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	230 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	235 
    -- CP-element group 234:  members (3) 
      -- CP-element group 234: 	 branch_block_stmt_1335/assign_stmt_1940_to_call_stmt_1956/type_cast_1943_update_completed_
      -- CP-element group 234: 	 branch_block_stmt_1335/assign_stmt_1940_to_call_stmt_1956/type_cast_1943_Update/$exit
      -- CP-element group 234: 	 branch_block_stmt_1335/assign_stmt_1940_to_call_stmt_1956/type_cast_1943_Update/ca
      -- 
    ca_3809_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 234_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1943_inst_ack_1, ack => maxPool3D_CP_2658_elements(234)); -- 
    -- CP-element group 235:  join  transition  output  bypass 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	232 
    -- CP-element group 235: 	234 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	236 
    -- CP-element group 235:  members (3) 
      -- CP-element group 235: 	 branch_block_stmt_1335/assign_stmt_1940_to_call_stmt_1956/call_stmt_1956_sample_start_
      -- CP-element group 235: 	 branch_block_stmt_1335/assign_stmt_1940_to_call_stmt_1956/call_stmt_1956_Sample/$entry
      -- CP-element group 235: 	 branch_block_stmt_1335/assign_stmt_1940_to_call_stmt_1956/call_stmt_1956_Sample/crr
      -- 
    crr_3817_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3817_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(235), ack => call_stmt_1956_call_req_0); -- 
    maxPool3D_cp_element_group_235: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_235"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2658_elements(232) & maxPool3D_CP_2658_elements(234);
      gj_maxPool3D_cp_element_group_235 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2658_elements(235), clk => clk, reset => reset); --
    end block;
    -- CP-element group 236:  transition  input  bypass 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	235 
    -- CP-element group 236: successors 
    -- CP-element group 236:  members (3) 
      -- CP-element group 236: 	 branch_block_stmt_1335/assign_stmt_1940_to_call_stmt_1956/call_stmt_1956_sample_completed_
      -- CP-element group 236: 	 branch_block_stmt_1335/assign_stmt_1940_to_call_stmt_1956/call_stmt_1956_Sample/$exit
      -- CP-element group 236: 	 branch_block_stmt_1335/assign_stmt_1940_to_call_stmt_1956/call_stmt_1956_Sample/cra
      -- 
    cra_3818_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 236_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1956_call_ack_0, ack => maxPool3D_CP_2658_elements(236)); -- 
    -- CP-element group 237:  transition  place  input  bypass 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	230 
    -- CP-element group 237: successors 
    -- CP-element group 237:  members (16) 
      -- CP-element group 237: 	 branch_block_stmt_1335/branch_block_stmt_1335__exit__
      -- CP-element group 237: 	 branch_block_stmt_1335/assign_stmt_1940_to_call_stmt_1956__exit__
      -- CP-element group 237: 	 branch_block_stmt_1335/return__
      -- CP-element group 237: 	 branch_block_stmt_1335/$exit
      -- CP-element group 237: 	 branch_block_stmt_1335/merge_stmt_1958__exit__
      -- CP-element group 237: 	 $exit
      -- CP-element group 237: 	 branch_block_stmt_1335/assign_stmt_1940_to_call_stmt_1956/$exit
      -- CP-element group 237: 	 branch_block_stmt_1335/assign_stmt_1940_to_call_stmt_1956/call_stmt_1956_update_completed_
      -- CP-element group 237: 	 branch_block_stmt_1335/assign_stmt_1940_to_call_stmt_1956/call_stmt_1956_Update/$exit
      -- CP-element group 237: 	 branch_block_stmt_1335/assign_stmt_1940_to_call_stmt_1956/call_stmt_1956_Update/cca
      -- CP-element group 237: 	 branch_block_stmt_1335/return___PhiReq/$entry
      -- CP-element group 237: 	 branch_block_stmt_1335/return___PhiReq/$exit
      -- CP-element group 237: 	 branch_block_stmt_1335/merge_stmt_1958_PhiReqMerge
      -- CP-element group 237: 	 branch_block_stmt_1335/merge_stmt_1958_PhiAck/$entry
      -- CP-element group 237: 	 branch_block_stmt_1335/merge_stmt_1958_PhiAck/$exit
      -- CP-element group 237: 	 branch_block_stmt_1335/merge_stmt_1958_PhiAck/dummy
      -- 
    cca_3823_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 237_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1956_call_ack_1, ack => maxPool3D_CP_2658_elements(237)); -- 
    -- CP-element group 238:  transition  output  delay-element  bypass 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	56 
    -- CP-element group 238: successors 
    -- CP-element group 238: 	242 
    -- CP-element group 238:  members (5) 
      -- CP-element group 238: 	 branch_block_stmt_1335/bbx_xnph_forx_xbody_PhiReq/$exit
      -- CP-element group 238: 	 branch_block_stmt_1335/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1561/$exit
      -- CP-element group 238: 	 branch_block_stmt_1335/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1561/phi_stmt_1561_sources/$exit
      -- CP-element group 238: 	 branch_block_stmt_1335/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1561/phi_stmt_1561_sources/type_cast_1565_konst_delay_trans
      -- CP-element group 238: 	 branch_block_stmt_1335/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1561/phi_stmt_1561_req
      -- 
    phi_stmt_1561_req_3846_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1561_req_3846_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(238), ack => phi_stmt_1561_req_0); -- 
    -- Element group maxPool3D_CP_2658_elements(238) is a control-delay.
    cp_element_238_delay: control_delay_element  generic map(name => " 238_delay", delay_value => 1)  port map(req => maxPool3D_CP_2658_elements(56), ack => maxPool3D_CP_2658_elements(238), clk => clk, reset =>reset);
    -- CP-element group 239:  transition  input  bypass 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	60 
    -- CP-element group 239: successors 
    -- CP-element group 239: 	241 
    -- CP-element group 239:  members (2) 
      -- CP-element group 239: 	 branch_block_stmt_1335/forx_xbody_forx_xbody_PhiReq/phi_stmt_1561/phi_stmt_1561_sources/type_cast_1567/SplitProtocol/Sample/$exit
      -- CP-element group 239: 	 branch_block_stmt_1335/forx_xbody_forx_xbody_PhiReq/phi_stmt_1561/phi_stmt_1561_sources/type_cast_1567/SplitProtocol/Sample/ra
      -- 
    ra_3866_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 239_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1567_inst_ack_0, ack => maxPool3D_CP_2658_elements(239)); -- 
    -- CP-element group 240:  transition  input  bypass 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	60 
    -- CP-element group 240: successors 
    -- CP-element group 240: 	241 
    -- CP-element group 240:  members (2) 
      -- CP-element group 240: 	 branch_block_stmt_1335/forx_xbody_forx_xbody_PhiReq/phi_stmt_1561/phi_stmt_1561_sources/type_cast_1567/SplitProtocol/Update/$exit
      -- CP-element group 240: 	 branch_block_stmt_1335/forx_xbody_forx_xbody_PhiReq/phi_stmt_1561/phi_stmt_1561_sources/type_cast_1567/SplitProtocol/Update/ca
      -- 
    ca_3871_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 240_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1567_inst_ack_1, ack => maxPool3D_CP_2658_elements(240)); -- 
    -- CP-element group 241:  join  transition  output  bypass 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	239 
    -- CP-element group 241: 	240 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	242 
    -- CP-element group 241:  members (6) 
      -- CP-element group 241: 	 branch_block_stmt_1335/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 241: 	 branch_block_stmt_1335/forx_xbody_forx_xbody_PhiReq/phi_stmt_1561/$exit
      -- CP-element group 241: 	 branch_block_stmt_1335/forx_xbody_forx_xbody_PhiReq/phi_stmt_1561/phi_stmt_1561_sources/$exit
      -- CP-element group 241: 	 branch_block_stmt_1335/forx_xbody_forx_xbody_PhiReq/phi_stmt_1561/phi_stmt_1561_sources/type_cast_1567/$exit
      -- CP-element group 241: 	 branch_block_stmt_1335/forx_xbody_forx_xbody_PhiReq/phi_stmt_1561/phi_stmt_1561_sources/type_cast_1567/SplitProtocol/$exit
      -- CP-element group 241: 	 branch_block_stmt_1335/forx_xbody_forx_xbody_PhiReq/phi_stmt_1561/phi_stmt_1561_req
      -- 
    phi_stmt_1561_req_3872_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1561_req_3872_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(241), ack => phi_stmt_1561_req_1); -- 
    maxPool3D_cp_element_group_241: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "maxPool3D_cp_element_group_241"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool3D_CP_2658_elements(239) & maxPool3D_CP_2658_elements(240);
      gj_maxPool3D_cp_element_group_241 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool3D_CP_2658_elements(241), clk => clk, reset => reset); --
    end block;
    -- CP-element group 242:  merge  transition  place  bypass 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	238 
    -- CP-element group 242: 	241 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	243 
    -- CP-element group 242:  members (2) 
      -- CP-element group 242: 	 branch_block_stmt_1335/merge_stmt_1560_PhiReqMerge
      -- CP-element group 242: 	 branch_block_stmt_1335/merge_stmt_1560_PhiAck/$entry
      -- 
    maxPool3D_CP_2658_elements(242) <= OrReduce(maxPool3D_CP_2658_elements(238) & maxPool3D_CP_2658_elements(241));
    -- CP-element group 243:  fork  transition  place  input  output  bypass 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	242 
    -- CP-element group 243: successors 
    -- CP-element group 243: 	57 
    -- CP-element group 243: 	58 
    -- CP-element group 243:  members (11) 
      -- CP-element group 243: 	 branch_block_stmt_1335/call_stmt_1570_to_assign_stmt_1581__entry__
      -- CP-element group 243: 	 branch_block_stmt_1335/merge_stmt_1560__exit__
      -- CP-element group 243: 	 branch_block_stmt_1335/call_stmt_1570_to_assign_stmt_1581/$entry
      -- CP-element group 243: 	 branch_block_stmt_1335/call_stmt_1570_to_assign_stmt_1581/call_stmt_1570_sample_start_
      -- CP-element group 243: 	 branch_block_stmt_1335/call_stmt_1570_to_assign_stmt_1581/call_stmt_1570_update_start_
      -- CP-element group 243: 	 branch_block_stmt_1335/call_stmt_1570_to_assign_stmt_1581/call_stmt_1570_Sample/$entry
      -- CP-element group 243: 	 branch_block_stmt_1335/call_stmt_1570_to_assign_stmt_1581/call_stmt_1570_Sample/crr
      -- CP-element group 243: 	 branch_block_stmt_1335/call_stmt_1570_to_assign_stmt_1581/call_stmt_1570_Update/$entry
      -- CP-element group 243: 	 branch_block_stmt_1335/call_stmt_1570_to_assign_stmt_1581/call_stmt_1570_Update/ccr
      -- CP-element group 243: 	 branch_block_stmt_1335/merge_stmt_1560_PhiAck/$exit
      -- CP-element group 243: 	 branch_block_stmt_1335/merge_stmt_1560_PhiAck/phi_stmt_1561_ack
      -- 
    phi_stmt_1561_ack_3877_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 243_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1561_ack_0, ack => maxPool3D_CP_2658_elements(243)); -- 
    crr_3110_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3110_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(243), ack => call_stmt_1570_call_req_0); -- 
    ccr_3115_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3115_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(243), ack => call_stmt_1570_call_req_1); -- 
    -- CP-element group 244:  merge  fork  transition  place  output  bypass 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	54 
    -- CP-element group 244: 	59 
    -- CP-element group 244: successors 
    -- CP-element group 244: 	61 
    -- CP-element group 244: 	62 
    -- CP-element group 244:  members (17) 
      -- CP-element group 244: 	 branch_block_stmt_1335/call_stmt_1605__entry__
      -- CP-element group 244: 	 branch_block_stmt_1335/assign_stmt_1597_to_assign_stmt_1602__entry__
      -- CP-element group 244: 	 branch_block_stmt_1335/merge_stmt_1590__exit__
      -- CP-element group 244: 	 branch_block_stmt_1335/assign_stmt_1597_to_assign_stmt_1602__exit__
      -- CP-element group 244: 	 branch_block_stmt_1335/assign_stmt_1597_to_assign_stmt_1602/$entry
      -- CP-element group 244: 	 branch_block_stmt_1335/assign_stmt_1597_to_assign_stmt_1602/$exit
      -- CP-element group 244: 	 branch_block_stmt_1335/call_stmt_1605/$entry
      -- CP-element group 244: 	 branch_block_stmt_1335/call_stmt_1605/call_stmt_1605_sample_start_
      -- CP-element group 244: 	 branch_block_stmt_1335/call_stmt_1605/call_stmt_1605_update_start_
      -- CP-element group 244: 	 branch_block_stmt_1335/call_stmt_1605/call_stmt_1605_Sample/$entry
      -- CP-element group 244: 	 branch_block_stmt_1335/call_stmt_1605/call_stmt_1605_Sample/crr
      -- CP-element group 244: 	 branch_block_stmt_1335/call_stmt_1605/call_stmt_1605_Update/$entry
      -- CP-element group 244: 	 branch_block_stmt_1335/call_stmt_1605/call_stmt_1605_Update/ccr
      -- CP-element group 244: 	 branch_block_stmt_1335/merge_stmt_1590_PhiReqMerge
      -- CP-element group 244: 	 branch_block_stmt_1335/merge_stmt_1590_PhiAck/$entry
      -- CP-element group 244: 	 branch_block_stmt_1335/merge_stmt_1590_PhiAck/$exit
      -- CP-element group 244: 	 branch_block_stmt_1335/merge_stmt_1590_PhiAck/dummy
      -- 
    crr_3149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(244), ack => call_stmt_1605_call_req_0); -- 
    ccr_3154_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3154_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool3D_CP_2658_elements(244), ack => call_stmt_1605_call_req_1); -- 
    maxPool3D_CP_2658_elements(244) <= OrReduce(maxPool3D_CP_2658_elements(54) & maxPool3D_CP_2658_elements(59));
    maxPool3D_do_while_stmt_1648_terminator_3474: loop_terminator -- 
      generic map (name => " maxPool3D_do_while_stmt_1648_terminator_3474", max_iterations_in_flight =>15) 
      port map(loop_body_exit => maxPool3D_CP_2658_elements(74),loop_continue => maxPool3D_CP_2658_elements(179),loop_terminate => maxPool3D_CP_2658_elements(178),loop_back => maxPool3D_CP_2658_elements(72),loop_exit => maxPool3D_CP_2658_elements(71),clk => clk, reset => reset); -- 
    phi_stmt_1650_phi_seq_3264_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= maxPool3D_CP_2658_elements(87);
      maxPool3D_CP_2658_elements(92)<= src_sample_reqs(0);
      src_sample_acks(0)  <= maxPool3D_CP_2658_elements(96);
      maxPool3D_CP_2658_elements(93)<= src_update_reqs(0);
      src_update_acks(0)  <= maxPool3D_CP_2658_elements(97);
      maxPool3D_CP_2658_elements(88) <= phi_mux_reqs(0);
      triggers(1)  <= maxPool3D_CP_2658_elements(89);
      maxPool3D_CP_2658_elements(98)<= src_sample_reqs(1);
      src_sample_acks(1)  <= maxPool3D_CP_2658_elements(98);
      maxPool3D_CP_2658_elements(99)<= src_update_reqs(1);
      src_update_acks(1)  <= maxPool3D_CP_2658_elements(100);
      maxPool3D_CP_2658_elements(90) <= phi_mux_reqs(1);
      phi_stmt_1650_phi_seq_3264 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1650_phi_seq_3264") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => maxPool3D_CP_2658_elements(79), 
          phi_sample_ack => maxPool3D_CP_2658_elements(85), 
          phi_update_req => maxPool3D_CP_2658_elements(81), 
          phi_update_ack => maxPool3D_CP_2658_elements(86), 
          phi_mux_ack => maxPool3D_CP_2658_elements(91), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1655_phi_seq_3308_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= maxPool3D_CP_2658_elements(108);
      maxPool3D_CP_2658_elements(113)<= src_sample_reqs(0);
      src_sample_acks(0)  <= maxPool3D_CP_2658_elements(117);
      maxPool3D_CP_2658_elements(114)<= src_update_reqs(0);
      src_update_acks(0)  <= maxPool3D_CP_2658_elements(118);
      maxPool3D_CP_2658_elements(109) <= phi_mux_reqs(0);
      triggers(1)  <= maxPool3D_CP_2658_elements(110);
      maxPool3D_CP_2658_elements(119)<= src_sample_reqs(1);
      src_sample_acks(1)  <= maxPool3D_CP_2658_elements(119);
      maxPool3D_CP_2658_elements(120)<= src_update_reqs(1);
      src_update_acks(1)  <= maxPool3D_CP_2658_elements(121);
      maxPool3D_CP_2658_elements(111) <= phi_mux_reqs(1);
      phi_stmt_1655_phi_seq_3308 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1655_phi_seq_3308") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => maxPool3D_CP_2658_elements(104), 
          phi_sample_ack => maxPool3D_CP_2658_elements(105), 
          phi_update_req => maxPool3D_CP_2658_elements(106), 
          phi_update_ack => maxPool3D_CP_2658_elements(107), 
          phi_mux_ack => maxPool3D_CP_2658_elements(112), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1660_phi_seq_3352_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= maxPool3D_CP_2658_elements(129);
      maxPool3D_CP_2658_elements(134)<= src_sample_reqs(0);
      src_sample_acks(0)  <= maxPool3D_CP_2658_elements(138);
      maxPool3D_CP_2658_elements(135)<= src_update_reqs(0);
      src_update_acks(0)  <= maxPool3D_CP_2658_elements(139);
      maxPool3D_CP_2658_elements(130) <= phi_mux_reqs(0);
      triggers(1)  <= maxPool3D_CP_2658_elements(131);
      maxPool3D_CP_2658_elements(140)<= src_sample_reqs(1);
      src_sample_acks(1)  <= maxPool3D_CP_2658_elements(140);
      maxPool3D_CP_2658_elements(141)<= src_update_reqs(1);
      src_update_acks(1)  <= maxPool3D_CP_2658_elements(142);
      maxPool3D_CP_2658_elements(132) <= phi_mux_reqs(1);
      phi_stmt_1660_phi_seq_3352 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1660_phi_seq_3352") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => maxPool3D_CP_2658_elements(125), 
          phi_sample_ack => maxPool3D_CP_2658_elements(126), 
          phi_update_req => maxPool3D_CP_2658_elements(127), 
          phi_update_ack => maxPool3D_CP_2658_elements(128), 
          phi_mux_ack => maxPool3D_CP_2658_elements(133), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_3216_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= maxPool3D_CP_2658_elements(75);
        preds(1)  <= maxPool3D_CP_2658_elements(76);
        entry_tmerge_3216 : transition_merge -- 
          generic map(name => " entry_tmerge_3216")
          port map (preds => preds, symbol_out => maxPool3D_CP_2658_elements(77));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal NOT_u1_u1_1810_wire : std_logic_vector(0 downto 0);
    signal add101_1629 : std_logic_vector(31 downto 0);
    signal add117_1687 : std_logic_vector(31 downto 0);
    signal add119_1697 : std_logic_vector(31 downto 0);
    signal add132_1713 : std_logic_vector(31 downto 0);
    signal add135_1723 : std_logic_vector(31 downto 0);
    signal add13_1385 : std_logic_vector(15 downto 0);
    signal add142_1728 : std_logic_vector(31 downto 0);
    signal add146_1733 : std_logic_vector(31 downto 0);
    signal add149_1738 : std_logic_vector(31 downto 0);
    signal add23_1410 : std_logic_vector(15 downto 0);
    signal add33_1435 : std_logic_vector(15 downto 0);
    signal add43_1460 : std_logic_vector(31 downto 0);
    signal add53_1485 : std_logic_vector(15 downto 0);
    signal add_1360 : std_logic_vector(31 downto 0);
    signal call11_1376 : std_logic_vector(7 downto 0);
    signal call150_1745 : std_logic_vector(7 downto 0);
    signal call16_1388 : std_logic_vector(7 downto 0);
    signal call180_1824 : std_logic_vector(63 downto 0);
    signal call21_1401 : std_logic_vector(7 downto 0);
    signal call26_1413 : std_logic_vector(7 downto 0);
    signal call2_1351 : std_logic_vector(7 downto 0);
    signal call31_1426 : std_logic_vector(7 downto 0);
    signal call36_1438 : std_logic_vector(7 downto 0);
    signal call41_1451 : std_logic_vector(7 downto 0);
    signal call46_1463 : std_logic_vector(7 downto 0);
    signal call51_1476 : std_logic_vector(7 downto 0);
    signal call6_1363 : std_logic_vector(7 downto 0);
    signal call89_1605 : std_logic_vector(63 downto 0);
    signal call_1338 : std_logic_vector(7 downto 0);
    signal chlx_x0_1660 : std_logic_vector(15 downto 0);
    signal chlx_x0_at_entry_1642 : std_logic_vector(15 downto 0);
    signal chlx_x1_1775 : std_logic_vector(15 downto 0);
    signal cmp157_1756 : std_logic_vector(0 downto 0);
    signal cmp165_1780 : std_logic_vector(0 downto 0);
    signal cmp175_1804 : std_logic_vector(0 downto 0);
    signal cmp257_1506 : std_logic_vector(0 downto 0);
    signal colx_x1_1655 : std_logic_vector(15 downto 0);
    signal colx_x1_1751_delayed_1_0_1763 : std_logic_vector(15 downto 0);
    signal colx_x1_at_entry_1637 : std_logic_vector(15 downto 0);
    signal colx_x2_1799 : std_logic_vector(15 downto 0);
    signal conv100_1614 : std_logic_vector(31 downto 0);
    signal conv107_1669 : std_logic_vector(31 downto 0);
    signal conv111_1673 : std_logic_vector(31 downto 0);
    signal conv113_1618 : std_logic_vector(31 downto 0);
    signal conv115_1677 : std_logic_vector(31 downto 0);
    signal conv12_1380 : std_logic_vector(15 downto 0);
    signal conv181_1829 : std_logic_vector(63 downto 0);
    signal conv187_1838 : std_logic_vector(7 downto 0);
    signal conv192_1848 : std_logic_vector(7 downto 0);
    signal conv198_1858 : std_logic_vector(7 downto 0);
    signal conv19_1392 : std_logic_vector(15 downto 0);
    signal conv1_1342 : std_logic_vector(31 downto 0);
    signal conv204_1868 : std_logic_vector(7 downto 0);
    signal conv210_1878 : std_logic_vector(7 downto 0);
    signal conv216_1888 : std_logic_vector(7 downto 0);
    signal conv222_1898 : std_logic_vector(7 downto 0);
    signal conv228_1908 : std_logic_vector(7 downto 0);
    signal conv22_1405 : std_logic_vector(15 downto 0);
    signal conv250_1940 : std_logic_vector(31 downto 0);
    signal conv253_1944 : std_logic_vector(31 downto 0);
    signal conv29_1417 : std_logic_vector(15 downto 0);
    signal conv32_1430 : std_logic_vector(15 downto 0);
    signal conv39_1442 : std_logic_vector(31 downto 0);
    signal conv3_1355 : std_logic_vector(31 downto 0);
    signal conv42_1455 : std_logic_vector(31 downto 0);
    signal conv49_1467 : std_logic_vector(15 downto 0);
    signal conv52_1480 : std_logic_vector(15 downto 0);
    signal conv59_1490 : std_logic_vector(31 downto 0);
    signal conv90_1821 : std_logic_vector(63 downto 0);
    signal conv98_1610 : std_logic_vector(31 downto 0);
    signal conv9_1367 : std_logic_vector(15 downto 0);
    signal exitcond1_1581 : std_logic_vector(0 downto 0);
    signal iNsTr_14_1545 : std_logic_vector(63 downto 0);
    signal iNsTr_20_1561 : std_logic_vector(63 downto 0);
    signal inc152_1751 : std_logic_vector(15 downto 0);
    signal inc160_1760 : std_logic_vector(15 downto 0);
    signal inc160x_xcolx_x1_1768 : std_logic_vector(15 downto 0);
    signal inc169_1784 : std_logic_vector(15 downto 0);
    signal inc169x_xrowx_x1_1792 : std_logic_vector(15 downto 0);
    signal indvarx_xnext_1576 : std_logic_vector(63 downto 0);
    signal mul116_1682 : std_logic_vector(31 downto 0);
    signal mul118_1692 : std_logic_vector(31 downto 0);
    signal mul131_1708 : std_logic_vector(31 downto 0);
    signal mul133_1624 : std_logic_vector(31 downto 0);
    signal mul251_1949 : std_logic_vector(31 downto 0);
    signal mul254_1954 : std_logic_vector(31 downto 0);
    signal mul62_1500 : std_logic_vector(31 downto 0);
    signal mul86_1602 : std_logic_vector(15 downto 0);
    signal mul_1495 : std_logic_vector(31 downto 0);
    signal rowx_x1_1650 : std_logic_vector(15 downto 0);
    signal rowx_x1_1772_delayed_2_0_1787 : std_logic_vector(15 downto 0);
    signal rowx_x1_at_entry_1632 : std_logic_vector(15 downto 0);
    signal shl10_1373 : std_logic_vector(15 downto 0);
    signal shl120_1703 : std_logic_vector(31 downto 0);
    signal shl134_1718 : std_logic_vector(31 downto 0);
    signal shl20_1398 : std_logic_vector(15 downto 0);
    signal shl30_1423 : std_logic_vector(15 downto 0);
    signal shl40_1448 : std_logic_vector(31 downto 0);
    signal shl50_1473 : std_logic_vector(15 downto 0);
    signal shl_1348 : std_logic_vector(31 downto 0);
    signal shr189_1844 : std_logic_vector(63 downto 0);
    signal shr195_1854 : std_logic_vector(63 downto 0);
    signal shr201_1864 : std_logic_vector(63 downto 0);
    signal shr207_1874 : std_logic_vector(63 downto 0);
    signal shr213_1884 : std_logic_vector(63 downto 0);
    signal shr219_1894 : std_logic_vector(63 downto 0);
    signal shr225_1904 : std_logic_vector(63 downto 0);
    signal shr79255_1597 : std_logic_vector(15 downto 0);
    signal sub_1834 : std_logic_vector(63 downto 0);
    signal tmp260_1523 : std_logic_vector(31 downto 0);
    signal tmp261_1529 : std_logic_vector(31 downto 0);
    signal tmp261x_xop_1541 : std_logic_vector(31 downto 0);
    signal tmp262_1535 : std_logic_vector(0 downto 0);
    signal tmp265_1558 : std_logic_vector(63 downto 0);
    signal tmp_1518 : std_logic_vector(31 downto 0);
    signal type_cast_1346_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1371_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1396_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1421_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1446_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1471_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1504_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1527_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1533_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1539_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1549_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1556_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1565_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1567_wire : std_logic_vector(63 downto 0);
    signal type_cast_1574_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1595_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1622_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1653_wire : std_logic_vector(15 downto 0);
    signal type_cast_1658_wire : std_logic_vector(15 downto 0);
    signal type_cast_1663_wire : std_logic_vector(15 downto 0);
    signal type_cast_1701_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1749_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1772_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1796_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1819_wire : std_logic_vector(63 downto 0);
    signal type_cast_1827_wire : std_logic_vector(63 downto 0);
    signal type_cast_1842_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1852_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1862_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1872_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1882_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1892_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1902_wire_constant : std_logic_vector(63 downto 0);
    signal whilex_xbody_whilex_xend_taken_1807 : std_logic_vector(0 downto 0);
    signal xx_xop_1551 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    chlx_x0_at_entry_1642 <= "0000000000000000";
    colx_x1_at_entry_1637 <= "0000000000000000";
    rowx_x1_at_entry_1632 <= "0000000000000000";
    type_cast_1346_wire_constant <= "00000000000000000000000000001000";
    type_cast_1371_wire_constant <= "0000000000001000";
    type_cast_1396_wire_constant <= "0000000000001000";
    type_cast_1421_wire_constant <= "0000000000001000";
    type_cast_1446_wire_constant <= "00000000000000000000000000001000";
    type_cast_1471_wire_constant <= "0000000000001000";
    type_cast_1504_wire_constant <= "00000000000000000000000000001111";
    type_cast_1527_wire_constant <= "00000000000000000000000000000100";
    type_cast_1533_wire_constant <= "00000000000000000000000000000001";
    type_cast_1539_wire_constant <= "11111111111111111111111111111111";
    type_cast_1549_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1556_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1565_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1574_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1595_wire_constant <= "0000000000000100";
    type_cast_1622_wire_constant <= "00000000000000000000000000000001";
    type_cast_1701_wire_constant <= "00000000000000000000000000000010";
    type_cast_1749_wire_constant <= "0000000000000001";
    type_cast_1772_wire_constant <= "0000000000000000";
    type_cast_1796_wire_constant <= "0000000000000000";
    type_cast_1842_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1852_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1862_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1872_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1882_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1892_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1902_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    phi_stmt_1561: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1565_wire_constant & type_cast_1567_wire;
      req <= phi_stmt_1561_req_0 & phi_stmt_1561_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1561",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1561_ack_0,
          idata => idata,
          odata => iNsTr_20_1561,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1561
    phi_stmt_1650: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1653_wire & rowx_x1_at_entry_1632;
      req <= phi_stmt_1650_req_0 & phi_stmt_1650_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1650",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1650_ack_0,
          idata => idata,
          odata => rowx_x1_1650,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1650
    phi_stmt_1655: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1658_wire & colx_x1_at_entry_1637;
      req <= phi_stmt_1655_req_0 & phi_stmt_1655_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1655",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1655_ack_0,
          idata => idata,
          odata => colx_x1_1655,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1655
    phi_stmt_1660: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1663_wire & chlx_x0_at_entry_1642;
      req <= phi_stmt_1660_req_0 & phi_stmt_1660_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1660",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1660_ack_0,
          idata => idata,
          odata => chlx_x0_1660,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1660
    -- flow-through select operator MUX_1557_inst
    tmp265_1558 <= xx_xop_1551 when (tmp262_1535(0) /=  '0') else type_cast_1556_wire_constant;
    -- flow-through select operator MUX_1774_inst
    chlx_x1_1775 <= type_cast_1772_wire_constant when (cmp157_1756(0) /=  '0') else inc152_1751;
    -- flow-through select operator MUX_1798_inst
    colx_x2_1799 <= type_cast_1796_wire_constant when (cmp165_1780(0) /=  '0') else inc160x_xcolx_x1_1768;
    W_colx_x1_1751_delayed_1_0_1761_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_colx_x1_1751_delayed_1_0_1761_inst_req_0;
      W_colx_x1_1751_delayed_1_0_1761_inst_ack_0<= wack(0);
      rreq(0) <= W_colx_x1_1751_delayed_1_0_1761_inst_req_1;
      W_colx_x1_1751_delayed_1_0_1761_inst_ack_1<= rack(0);
      W_colx_x1_1751_delayed_1_0_1761_inst : InterlockBuffer generic map ( -- 
        name => "W_colx_x1_1751_delayed_1_0_1761_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => colx_x1_1655,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => colx_x1_1751_delayed_1_0_1763,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_rowx_x1_1772_delayed_2_0_1785_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_rowx_x1_1772_delayed_2_0_1785_inst_req_0;
      W_rowx_x1_1772_delayed_2_0_1785_inst_ack_0<= wack(0);
      rreq(0) <= W_rowx_x1_1772_delayed_2_0_1785_inst_req_1;
      W_rowx_x1_1772_delayed_2_0_1785_inst_ack_1<= rack(0);
      W_rowx_x1_1772_delayed_2_0_1785_inst : InterlockBuffer generic map ( -- 
        name => "W_rowx_x1_1772_delayed_2_0_1785_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rowx_x1_1650,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => rowx_x1_1772_delayed_2_0_1787,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock W_whilex_xbody_whilex_xend_taken_1805_inst
    process(cmp175_1804) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := cmp175_1804(0 downto 0);
      whilex_xbody_whilex_xend_taken_1807 <= tmp_var; -- 
    end process;
    type_cast_1341_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1341_inst_req_0;
      type_cast_1341_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1341_inst_req_1;
      type_cast_1341_inst_ack_1<= rack(0);
      type_cast_1341_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1341_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_1338,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1_1342,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1354_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1354_inst_req_0;
      type_cast_1354_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1354_inst_req_1;
      type_cast_1354_inst_ack_1<= rack(0);
      type_cast_1354_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1354_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_1351,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv3_1355,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1366_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1366_inst_req_0;
      type_cast_1366_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1366_inst_req_1;
      type_cast_1366_inst_ack_1<= rack(0);
      type_cast_1366_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1366_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call6_1363,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv9_1367,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1379_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1379_inst_req_0;
      type_cast_1379_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1379_inst_req_1;
      type_cast_1379_inst_ack_1<= rack(0);
      type_cast_1379_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1379_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call11_1376,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv12_1380,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1391_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1391_inst_req_0;
      type_cast_1391_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1391_inst_req_1;
      type_cast_1391_inst_ack_1<= rack(0);
      type_cast_1391_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1391_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call16_1388,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv19_1392,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1404_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1404_inst_req_0;
      type_cast_1404_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1404_inst_req_1;
      type_cast_1404_inst_ack_1<= rack(0);
      type_cast_1404_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1404_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call21_1401,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv22_1405,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1416_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1416_inst_req_0;
      type_cast_1416_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1416_inst_req_1;
      type_cast_1416_inst_ack_1<= rack(0);
      type_cast_1416_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1416_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call26_1413,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv29_1417,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1429_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1429_inst_req_0;
      type_cast_1429_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1429_inst_req_1;
      type_cast_1429_inst_ack_1<= rack(0);
      type_cast_1429_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1429_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call31_1426,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv32_1430,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1441_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1441_inst_req_0;
      type_cast_1441_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1441_inst_req_1;
      type_cast_1441_inst_ack_1<= rack(0);
      type_cast_1441_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1441_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call36_1438,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv39_1442,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1454_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1454_inst_req_0;
      type_cast_1454_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1454_inst_req_1;
      type_cast_1454_inst_ack_1<= rack(0);
      type_cast_1454_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1454_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call41_1451,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv42_1455,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1466_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1466_inst_req_0;
      type_cast_1466_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1466_inst_req_1;
      type_cast_1466_inst_ack_1<= rack(0);
      type_cast_1466_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1466_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call46_1463,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv49_1467,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1479_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1479_inst_req_0;
      type_cast_1479_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1479_inst_req_1;
      type_cast_1479_inst_ack_1<= rack(0);
      type_cast_1479_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1479_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call51_1476,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv52_1480,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1489_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1489_inst_req_0;
      type_cast_1489_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1489_inst_req_1;
      type_cast_1489_inst_ack_1<= rack(0);
      type_cast_1489_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1489_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add23_1410,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv59_1490,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1544_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1544_inst_req_0;
      type_cast_1544_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1544_inst_req_1;
      type_cast_1544_inst_ack_1<= rack(0);
      type_cast_1544_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1544_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp261x_xop_1541,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_14_1545,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1567_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1567_inst_req_0;
      type_cast_1567_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1567_inst_req_1;
      type_cast_1567_inst_ack_1<= rack(0);
      type_cast_1567_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1567_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1576,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1567_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1609_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1609_inst_req_0;
      type_cast_1609_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1609_inst_req_1;
      type_cast_1609_inst_ack_1<= rack(0);
      type_cast_1609_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1609_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr79255_1597,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv98_1610,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1613_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1613_inst_req_0;
      type_cast_1613_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1613_inst_req_1;
      type_cast_1613_inst_ack_1<= rack(0);
      type_cast_1613_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1613_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => mul86_1602,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv100_1614,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1617_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1617_inst_req_0;
      type_cast_1617_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1617_inst_req_1;
      type_cast_1617_inst_ack_1<= rack(0);
      type_cast_1617_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1617_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add33_1435,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv113_1618,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1653_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1653_inst_req_0;
      type_cast_1653_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1653_inst_req_1;
      type_cast_1653_inst_ack_1<= rack(0);
      type_cast_1653_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1653_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc169x_xrowx_x1_1792,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1653_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1658_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1658_inst_req_0;
      type_cast_1658_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1658_inst_req_1;
      type_cast_1658_inst_ack_1<= rack(0);
      type_cast_1658_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1658_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => colx_x2_1799,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1658_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1663_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1663_inst_req_0;
      type_cast_1663_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1663_inst_req_1;
      type_cast_1663_inst_ack_1<= rack(0);
      type_cast_1663_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1663_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => chlx_x1_1775,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1663_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1668_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1668_inst_req_0;
      type_cast_1668_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1668_inst_req_1;
      type_cast_1668_inst_ack_1<= rack(0);
      type_cast_1668_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1668_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => chlx_x0_1660,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv107_1669,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1672_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1672_inst_req_0;
      type_cast_1672_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1672_inst_req_1;
      type_cast_1672_inst_ack_1<= rack(0);
      type_cast_1672_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1672_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => colx_x1_1655,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv111_1673,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1676_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1676_inst_req_0;
      type_cast_1676_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1676_inst_req_1;
      type_cast_1676_inst_ack_1<= rack(0);
      type_cast_1676_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1676_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rowx_x1_1650,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv115_1677,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1759_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1759_inst_req_0;
      type_cast_1759_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1759_inst_req_1;
      type_cast_1759_inst_ack_1<= rack(0);
      type_cast_1759_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1759_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp157_1756,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc160_1760,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1783_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1783_inst_req_0;
      type_cast_1783_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1783_inst_req_1;
      type_cast_1783_inst_ack_1<= rack(0);
      type_cast_1783_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1783_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp165_1780,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc169_1784,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1820_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1820_inst_req_0;
      type_cast_1820_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1820_inst_req_1;
      type_cast_1820_inst_ack_1<= rack(0);
      type_cast_1820_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1820_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1819_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv90_1821,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1828_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1828_inst_req_0;
      type_cast_1828_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1828_inst_req_1;
      type_cast_1828_inst_ack_1<= rack(0);
      type_cast_1828_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1828_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1827_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv181_1829,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1837_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1837_inst_req_0;
      type_cast_1837_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1837_inst_req_1;
      type_cast_1837_inst_ack_1<= rack(0);
      type_cast_1837_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1837_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub_1834,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv187_1838,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1847_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1847_inst_req_0;
      type_cast_1847_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1847_inst_req_1;
      type_cast_1847_inst_ack_1<= rack(0);
      type_cast_1847_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1847_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr189_1844,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv192_1848,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1857_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1857_inst_req_0;
      type_cast_1857_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1857_inst_req_1;
      type_cast_1857_inst_ack_1<= rack(0);
      type_cast_1857_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1857_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr195_1854,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv198_1858,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1867_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1867_inst_req_0;
      type_cast_1867_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1867_inst_req_1;
      type_cast_1867_inst_ack_1<= rack(0);
      type_cast_1867_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1867_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr201_1864,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv204_1868,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1877_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1877_inst_req_0;
      type_cast_1877_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1877_inst_req_1;
      type_cast_1877_inst_ack_1<= rack(0);
      type_cast_1877_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1877_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr207_1874,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv210_1878,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1887_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1887_inst_req_0;
      type_cast_1887_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1887_inst_req_1;
      type_cast_1887_inst_ack_1<= rack(0);
      type_cast_1887_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1887_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr213_1884,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv216_1888,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1897_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1897_inst_req_0;
      type_cast_1897_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1897_inst_req_1;
      type_cast_1897_inst_ack_1<= rack(0);
      type_cast_1897_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1897_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr219_1894,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv222_1898,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1907_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1907_inst_req_0;
      type_cast_1907_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1907_inst_req_1;
      type_cast_1907_inst_ack_1<= rack(0);
      type_cast_1907_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1907_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr225_1904,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv228_1908,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1939_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1939_inst_req_0;
      type_cast_1939_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1939_inst_req_1;
      type_cast_1939_inst_ack_1<= rack(0);
      type_cast_1939_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1939_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add13_1385,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv250_1940,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1943_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1943_inst_req_0;
      type_cast_1943_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1943_inst_req_1;
      type_cast_1943_inst_ack_1<= rack(0);
      type_cast_1943_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1943_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add53_1485,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv253_1944,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    do_while_stmt_1648_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NOT_u1_u1_1810_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1648_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1648_branch_req_0,
          ack0 => do_while_stmt_1648_branch_ack_0,
          ack1 => do_while_stmt_1648_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1507_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp257_1506;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1507_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1507_branch_req_0,
          ack0 => if_stmt_1507_branch_ack_0,
          ack1 => if_stmt_1507_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1582_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond1_1581;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1582_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1582_branch_req_0,
          ack0 => if_stmt_1582_branch_ack_0,
          ack1 => if_stmt_1582_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1811_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= whilex_xbody_whilex_xend_taken_1807;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1811_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1811_branch_req_0,
          ack0 => if_stmt_1811_branch_ack_0,
          ack1 => if_stmt_1811_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1750_inst
    process(chlx_x0_1660) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(chlx_x0_1660, type_cast_1749_wire_constant, tmp_var);
      inc152_1751 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1767_inst
    process(inc160_1760, colx_x1_1751_delayed_1_0_1763) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc160_1760, colx_x1_1751_delayed_1_0_1763, tmp_var);
      inc160x_xcolx_x1_1768 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1791_inst
    process(inc169_1784, rowx_x1_1772_delayed_2_0_1787) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc169_1784, rowx_x1_1772_delayed_2_0_1787, tmp_var);
      inc169x_xrowx_x1_1792 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1540_inst
    process(tmp261_1529) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp261_1529, type_cast_1539_wire_constant, tmp_var);
      tmp261x_xop_1541 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1628_inst
    process(conv100_1614, conv98_1610) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv100_1614, conv98_1610, tmp_var);
      add101_1629 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1686_inst
    process(conv111_1673, mul116_1682) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv111_1673, mul116_1682, tmp_var);
      add117_1687 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1696_inst
    process(mul118_1692, conv107_1669) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul118_1692, conv107_1669, tmp_var);
      add119_1697 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1712_inst
    process(conv111_1673, mul131_1708) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv111_1673, mul131_1708, tmp_var);
      add132_1713 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1722_inst
    process(shl134_1718, conv107_1669) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shl134_1718, conv107_1669, tmp_var);
      add135_1723 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1727_inst
    process(add135_1723, conv98_1610) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add135_1723, conv98_1610, tmp_var);
      add142_1728 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1732_inst
    process(add135_1723, conv100_1614) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add135_1723, conv100_1614, tmp_var);
      add146_1733 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1737_inst
    process(add101_1629, add135_1723) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add101_1629, add135_1723, tmp_var);
      add149_1738 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1550_inst
    process(iNsTr_14_1545) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_14_1545, type_cast_1549_wire_constant, tmp_var);
      xx_xop_1551 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1575_inst
    process(iNsTr_20_1561) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_20_1561, type_cast_1574_wire_constant, tmp_var);
      indvarx_xnext_1576 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_1755_inst
    process(inc152_1751, shr79255_1597) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc152_1751, shr79255_1597, tmp_var);
      cmp157_1756 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_1779_inst
    process(inc160x_xcolx_x1_1768, add33_1435) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc160x_xcolx_x1_1768, add33_1435, tmp_var);
      cmp165_1780 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_1803_inst
    process(inc169x_xrowx_x1_1792, add13_1385) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(inc169x_xrowx_x1_1792, add13_1385, tmp_var);
      cmp175_1804 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1580_inst
    process(indvarx_xnext_1576, tmp265_1558) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_1576, tmp265_1558, tmp_var);
      exitcond1_1581 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_1596_inst
    process(add53_1485) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add53_1485, type_cast_1595_wire_constant, tmp_var);
      shr79255_1597 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1528_inst
    process(tmp260_1523) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp260_1523, type_cast_1527_wire_constant, tmp_var);
      tmp261_1529 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1843_inst
    process(sub_1834) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1834, type_cast_1842_wire_constant, tmp_var);
      shr189_1844 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1853_inst
    process(sub_1834) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1834, type_cast_1852_wire_constant, tmp_var);
      shr195_1854 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1863_inst
    process(sub_1834) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1834, type_cast_1862_wire_constant, tmp_var);
      shr201_1864 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1873_inst
    process(sub_1834) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1834, type_cast_1872_wire_constant, tmp_var);
      shr207_1874 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1883_inst
    process(sub_1834) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1834, type_cast_1882_wire_constant, tmp_var);
      shr213_1884 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1893_inst
    process(sub_1834) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1834, type_cast_1892_wire_constant, tmp_var);
      shr219_1894 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1903_inst
    process(sub_1834) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1834, type_cast_1902_wire_constant, tmp_var);
      shr225_1904 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1601_inst
    process(shr79255_1597, add23_1410) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(shr79255_1597, add23_1410, tmp_var);
      mul86_1602 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1494_inst
    process(conv59_1490, add_1360) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv59_1490, add_1360, tmp_var);
      mul_1495 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1499_inst
    process(mul_1495, add43_1460) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_1495, add43_1460, tmp_var);
      mul62_1500 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1517_inst
    process(add_1360, add43_1460) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add_1360, add43_1460, tmp_var);
      tmp_1518 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1522_inst
    process(tmp_1518, conv59_1490) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp_1518, conv59_1490, tmp_var);
      tmp260_1523 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1681_inst
    process(conv115_1677, conv113_1618) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv115_1677, conv113_1618, tmp_var);
      mul116_1682 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1691_inst
    process(add117_1687, conv98_1610) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add117_1687, conv98_1610, tmp_var);
      mul118_1692 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1707_inst
    process(conv115_1677, conv59_1490) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv115_1677, conv59_1490, tmp_var);
      mul131_1708 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1717_inst
    process(mul133_1624, add132_1713) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul133_1624, add132_1713, tmp_var);
      shl134_1718 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1948_inst
    process(conv113_1618, conv250_1940) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv113_1618, conv250_1940, tmp_var);
      mul251_1949 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1953_inst
    process(mul251_1949, conv253_1944) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul251_1949, conv253_1944, tmp_var);
      mul254_1954 <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_1810_inst
    process(cmp175_1804) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", cmp175_1804, tmp_var);
      NOT_u1_u1_1810_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u16_u16_1384_inst
    process(shl10_1373, conv12_1380) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl10_1373, conv12_1380, tmp_var);
      add13_1385 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_1409_inst
    process(shl20_1398, conv22_1405) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl20_1398, conv22_1405, tmp_var);
      add23_1410 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_1434_inst
    process(shl30_1423, conv32_1430) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl30_1423, conv32_1430, tmp_var);
      add33_1435 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_1484_inst
    process(shl50_1473, conv52_1480) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl50_1473, conv52_1480, tmp_var);
      add53_1485 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_1359_inst
    process(shl_1348, conv3_1355) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_1348, conv3_1355, tmp_var);
      add_1360 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_1459_inst
    process(shl40_1448, conv42_1455) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl40_1448, conv42_1455, tmp_var);
      add43_1460 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_1372_inst
    process(conv9_1367) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv9_1367, type_cast_1371_wire_constant, tmp_var);
      shl10_1373 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_1397_inst
    process(conv19_1392) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv19_1392, type_cast_1396_wire_constant, tmp_var);
      shl20_1398 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_1422_inst
    process(conv29_1417) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv29_1417, type_cast_1421_wire_constant, tmp_var);
      shl30_1423 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_1472_inst
    process(conv49_1467) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv49_1467, type_cast_1471_wire_constant, tmp_var);
      shl50_1473 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1347_inst
    process(conv1_1342) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv1_1342, type_cast_1346_wire_constant, tmp_var);
      shl_1348 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1447_inst
    process(conv39_1442) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv39_1442, type_cast_1446_wire_constant, tmp_var);
      shl40_1448 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1623_inst
    process(conv98_1610) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv98_1610, type_cast_1622_wire_constant, tmp_var);
      mul133_1624 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1702_inst
    process(add119_1697) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add119_1697, type_cast_1701_wire_constant, tmp_var);
      shl120_1703 <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_1833_inst
    process(conv181_1829, conv90_1821) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv181_1829, conv90_1821, tmp_var);
      sub_1834 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1505_inst
    process(mul62_1500) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul62_1500, type_cast_1504_wire_constant, tmp_var);
      cmp257_1506 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1534_inst
    process(tmp261_1529) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp261_1529, type_cast_1533_wire_constant, tmp_var);
      tmp262_1535 <= tmp_var; --
    end process;
    -- unary operator type_cast_1819_inst
    process(call89_1605) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call89_1605, tmp_var);
      type_cast_1819_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1827_inst
    process(call180_1824) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call180_1824, tmp_var);
      type_cast_1827_wire <= tmp_var; -- 
    end process;
    -- shared inport operator group (0) : RPIPE_maxpool_input_pipe_1450_inst RPIPE_maxpool_input_pipe_1412_inst RPIPE_maxpool_input_pipe_1400_inst RPIPE_maxpool_input_pipe_1437_inst RPIPE_maxpool_input_pipe_1475_inst RPIPE_maxpool_input_pipe_1387_inst RPIPE_maxpool_input_pipe_1425_inst RPIPE_maxpool_input_pipe_1462_inst RPIPE_maxpool_input_pipe_1375_inst RPIPE_maxpool_input_pipe_1362_inst RPIPE_maxpool_input_pipe_1350_inst RPIPE_maxpool_input_pipe_1337_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(95 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 11 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 11 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 11 downto 0);
      signal guard_vector : std_logic_vector( 11 downto 0);
      constant outBUFs : IntegerArray(11 downto 0) := (11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(11 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false);
      constant guardBuffering: IntegerArray(11 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2);
      -- 
    begin -- 
      reqL_unguarded(11) <= RPIPE_maxpool_input_pipe_1450_inst_req_0;
      reqL_unguarded(10) <= RPIPE_maxpool_input_pipe_1412_inst_req_0;
      reqL_unguarded(9) <= RPIPE_maxpool_input_pipe_1400_inst_req_0;
      reqL_unguarded(8) <= RPIPE_maxpool_input_pipe_1437_inst_req_0;
      reqL_unguarded(7) <= RPIPE_maxpool_input_pipe_1475_inst_req_0;
      reqL_unguarded(6) <= RPIPE_maxpool_input_pipe_1387_inst_req_0;
      reqL_unguarded(5) <= RPIPE_maxpool_input_pipe_1425_inst_req_0;
      reqL_unguarded(4) <= RPIPE_maxpool_input_pipe_1462_inst_req_0;
      reqL_unguarded(3) <= RPIPE_maxpool_input_pipe_1375_inst_req_0;
      reqL_unguarded(2) <= RPIPE_maxpool_input_pipe_1362_inst_req_0;
      reqL_unguarded(1) <= RPIPE_maxpool_input_pipe_1350_inst_req_0;
      reqL_unguarded(0) <= RPIPE_maxpool_input_pipe_1337_inst_req_0;
      RPIPE_maxpool_input_pipe_1450_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_maxpool_input_pipe_1412_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_maxpool_input_pipe_1400_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_maxpool_input_pipe_1437_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_maxpool_input_pipe_1475_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_maxpool_input_pipe_1387_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_maxpool_input_pipe_1425_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_maxpool_input_pipe_1462_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_maxpool_input_pipe_1375_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_maxpool_input_pipe_1362_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_maxpool_input_pipe_1350_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_maxpool_input_pipe_1337_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(11) <= RPIPE_maxpool_input_pipe_1450_inst_req_1;
      reqR_unguarded(10) <= RPIPE_maxpool_input_pipe_1412_inst_req_1;
      reqR_unguarded(9) <= RPIPE_maxpool_input_pipe_1400_inst_req_1;
      reqR_unguarded(8) <= RPIPE_maxpool_input_pipe_1437_inst_req_1;
      reqR_unguarded(7) <= RPIPE_maxpool_input_pipe_1475_inst_req_1;
      reqR_unguarded(6) <= RPIPE_maxpool_input_pipe_1387_inst_req_1;
      reqR_unguarded(5) <= RPIPE_maxpool_input_pipe_1425_inst_req_1;
      reqR_unguarded(4) <= RPIPE_maxpool_input_pipe_1462_inst_req_1;
      reqR_unguarded(3) <= RPIPE_maxpool_input_pipe_1375_inst_req_1;
      reqR_unguarded(2) <= RPIPE_maxpool_input_pipe_1362_inst_req_1;
      reqR_unguarded(1) <= RPIPE_maxpool_input_pipe_1350_inst_req_1;
      reqR_unguarded(0) <= RPIPE_maxpool_input_pipe_1337_inst_req_1;
      RPIPE_maxpool_input_pipe_1450_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_maxpool_input_pipe_1412_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_maxpool_input_pipe_1400_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_maxpool_input_pipe_1437_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_maxpool_input_pipe_1475_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_maxpool_input_pipe_1387_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_maxpool_input_pipe_1425_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_maxpool_input_pipe_1462_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_maxpool_input_pipe_1375_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_maxpool_input_pipe_1362_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_maxpool_input_pipe_1350_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_maxpool_input_pipe_1337_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      call41_1451 <= data_out(95 downto 88);
      call26_1413 <= data_out(87 downto 80);
      call21_1401 <= data_out(79 downto 72);
      call36_1438 <= data_out(71 downto 64);
      call51_1476 <= data_out(63 downto 56);
      call16_1388 <= data_out(55 downto 48);
      call31_1426 <= data_out(47 downto 40);
      call46_1463 <= data_out(39 downto 32);
      call11_1376 <= data_out(31 downto 24);
      call6_1363 <= data_out(23 downto 16);
      call2_1351 <= data_out(15 downto 8);
      call_1338 <= data_out(7 downto 0);
      maxpool_input_pipe_read_0_gI: SplitGuardInterface generic map(name => "maxpool_input_pipe_read_0_gI", nreqs => 12, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      maxpool_input_pipe_read_0: InputPortRevised -- 
        generic map ( name => "maxpool_input_pipe_read_0", data_width => 8,  num_reqs => 12,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => maxpool_input_pipe_pipe_read_req(0),
          oack => maxpool_input_pipe_pipe_read_ack(0),
          odata => maxpool_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_elapsed_time_pipe_1933_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_elapsed_time_pipe_1933_inst_req_0;
      WPIPE_elapsed_time_pipe_1933_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_elapsed_time_pipe_1933_inst_req_1;
      WPIPE_elapsed_time_pipe_1933_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= shr225_1904;
      elapsed_time_pipe_write_0_gI: SplitGuardInterface generic map(name => "elapsed_time_pipe_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      elapsed_time_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "elapsed_time_pipe", data_width => 64, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => elapsed_time_pipe_pipe_write_req(0),
          oack => elapsed_time_pipe_pipe_write_ack(0),
          odata => elapsed_time_pipe_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_maxpool_output_pipe_1918_inst WPIPE_maxpool_output_pipe_1930_inst WPIPE_maxpool_output_pipe_1927_inst WPIPE_maxpool_output_pipe_1924_inst WPIPE_maxpool_output_pipe_1921_inst WPIPE_maxpool_output_pipe_1915_inst WPIPE_maxpool_output_pipe_1912_inst WPIPE_maxpool_output_pipe_1909_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 7 downto 0);
      signal update_req, update_ack : BooleanArray( 7 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 7 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 7 downto 0);
      signal guard_vector : std_logic_vector( 7 downto 0);
      constant inBUFs : IntegerArray(7 downto 0) := (7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(7 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false);
      constant guardBuffering: IntegerArray(7 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2);
      -- 
    begin -- 
      sample_req_unguarded(7) <= WPIPE_maxpool_output_pipe_1918_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_maxpool_output_pipe_1930_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_maxpool_output_pipe_1927_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_maxpool_output_pipe_1924_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_maxpool_output_pipe_1921_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_maxpool_output_pipe_1915_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_maxpool_output_pipe_1912_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_maxpool_output_pipe_1909_inst_req_0;
      WPIPE_maxpool_output_pipe_1918_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_maxpool_output_pipe_1930_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_maxpool_output_pipe_1927_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_maxpool_output_pipe_1924_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_maxpool_output_pipe_1921_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_maxpool_output_pipe_1915_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_maxpool_output_pipe_1912_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_maxpool_output_pipe_1909_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(7) <= WPIPE_maxpool_output_pipe_1918_inst_req_1;
      update_req_unguarded(6) <= WPIPE_maxpool_output_pipe_1930_inst_req_1;
      update_req_unguarded(5) <= WPIPE_maxpool_output_pipe_1927_inst_req_1;
      update_req_unguarded(4) <= WPIPE_maxpool_output_pipe_1924_inst_req_1;
      update_req_unguarded(3) <= WPIPE_maxpool_output_pipe_1921_inst_req_1;
      update_req_unguarded(2) <= WPIPE_maxpool_output_pipe_1915_inst_req_1;
      update_req_unguarded(1) <= WPIPE_maxpool_output_pipe_1912_inst_req_1;
      update_req_unguarded(0) <= WPIPE_maxpool_output_pipe_1909_inst_req_1;
      WPIPE_maxpool_output_pipe_1918_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_maxpool_output_pipe_1930_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_maxpool_output_pipe_1927_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_maxpool_output_pipe_1924_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_maxpool_output_pipe_1921_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_maxpool_output_pipe_1915_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_maxpool_output_pipe_1912_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_maxpool_output_pipe_1909_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      data_in <= conv210_1878 & conv187_1838 & conv192_1848 & conv198_1858 & conv204_1868 & conv216_1888 & conv222_1898 & conv228_1908;
      maxpool_output_pipe_write_1_gI: SplitGuardInterface generic map(name => "maxpool_output_pipe_write_1_gI", nreqs => 8, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      maxpool_output_pipe_write_1: OutputPortRevised -- 
        generic map ( name => "maxpool_output_pipe", data_width => 8, num_reqs => 8, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => maxpool_output_pipe_pipe_write_req(0),
          oack => maxpool_output_pipe_pipe_write_ack(0),
          odata => maxpool_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared call operator group (0) : call_stmt_1570_call 
    fill_T_call_group_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1570_call_req_0;
      call_stmt_1570_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1570_call_req_1;
      call_stmt_1570_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      fill_T_call_group_0_gI: SplitGuardInterface generic map(name => "fill_T_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= iNsTr_20_1561;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 64,
        owidth => 64,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => fill_T_call_reqs(0),
          ackR => fill_T_call_acks(0),
          dataR => fill_T_call_data(63 downto 0),
          tagR => fill_T_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => fill_T_return_acks(0), -- cross-over
          ackL => fill_T_return_reqs(0), -- cross-over
          tagL => fill_T_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_1605_call call_stmt_1824_call 
    timer_call_group_1: Block -- 
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_1605_call_req_0;
      reqL_unguarded(0) <= call_stmt_1824_call_req_0;
      call_stmt_1605_call_ack_0 <= ackL_unguarded(1);
      call_stmt_1824_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_1605_call_req_1;
      reqR_unguarded(0) <= call_stmt_1824_call_req_1;
      call_stmt_1605_call_ack_1 <= ackR_unguarded(1);
      call_stmt_1824_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      timer_call_group_1_accessRegulator_0: access_regulator_base generic map (name => "timer_call_group_1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      timer_call_group_1_accessRegulator_1: access_regulator_base generic map (name => "timer_call_group_1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      timer_call_group_1_gI: SplitGuardInterface generic map(name => "timer_call_group_1_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      call89_1605 <= data_out(127 downto 64);
      call180_1824 <= data_out(63 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 2,
        nreqs => 2,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => timer_call_reqs(0),
          ackR => timer_call_acks(0),
          tagR => timer_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => timer_return_acks(0), -- cross-over
          ackL => timer_return_reqs(0), -- cross-over
          dataL => timer_return_data(63 downto 0),
          tagL => timer_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- shared call operator group (2) : call_stmt_1745_call 
    maxPool4_call_group_2: Block -- 
      signal data_in: std_logic_vector(159 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 17);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1745_call_req_0;
      call_stmt_1745_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1745_call_req_1;
      call_stmt_1745_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      maxPool4_call_group_2_gI: SplitGuardInterface generic map(name => "maxPool4_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= shl120_1703 & add135_1723 & add142_1728 & add146_1733 & add149_1738;
      call150_1745 <= data_out(7 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 160,
        owidth => 160,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => maxPool4_call_reqs(0),
          ackR => maxPool4_call_acks(0),
          dataR => maxPool4_call_data(159 downto 0),
          tagR => maxPool4_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 8,
          owidth => 8,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => maxPool4_return_acks(0), -- cross-over
          ackL => maxPool4_return_reqs(0), -- cross-over
          dataL => maxPool4_return_data(7 downto 0),
          tagL => maxPool4_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- shared call operator group (3) : call_stmt_1956_call 
    sendB_call_group_3: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1956_call_req_0;
      call_stmt_1956_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1956_call_req_1;
      call_stmt_1956_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      sendB_call_group_3_gI: SplitGuardInterface generic map(name => "sendB_call_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= mul254_1954;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 32,
        owidth => 32,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => sendB_call_reqs(0),
          ackR => sendB_call_acks(0),
          dataR => sendB_call_data(31 downto 0),
          tagR => sendB_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => sendB_return_acks(0), -- cross-over
          ackL => sendB_return_reqs(0), -- cross-over
          tagL => sendB_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 3
    -- 
  end Block; -- data_path
  -- 
end maxPool3D_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity maxPool4 is -- 
  generic (tag_length : integer); 
  port ( -- 
    addr : in  std_logic_vector(31 downto 0);
    addr1 : in  std_logic_vector(31 downto 0);
    addr2 : in  std_logic_vector(31 downto 0);
    addr3 : in  std_logic_vector(31 downto 0);
    addr4 : in  std_logic_vector(31 downto 0);
    output : out  std_logic_vector(7 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(255 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(2 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity maxPool4;
architecture maxPool4_arch of maxPool4 is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 160)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 8)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal addr_buffer :  std_logic_vector(31 downto 0);
  signal addr_update_enable: Boolean;
  signal addr1_buffer :  std_logic_vector(31 downto 0);
  signal addr1_update_enable: Boolean;
  signal addr2_buffer :  std_logic_vector(31 downto 0);
  signal addr2_update_enable: Boolean;
  signal addr3_buffer :  std_logic_vector(31 downto 0);
  signal addr3_update_enable: Boolean;
  signal addr4_buffer :  std_logic_vector(31 downto 0);
  signal addr4_update_enable: Boolean;
  -- output port buffer signals
  signal output_buffer :  std_logic_vector(7 downto 0);
  signal output_update_enable: Boolean;
  signal maxPool4_CP_346_start: Boolean;
  signal maxPool4_CP_346_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal slice_246_inst_ack_0 : boolean;
  signal slice_266_inst_ack_0 : boolean;
  signal slice_270_inst_ack_1 : boolean;
  signal slice_246_inst_req_0 : boolean;
  signal slice_242_inst_ack_1 : boolean;
  signal slice_238_inst_req_1 : boolean;
  signal slice_242_inst_req_1 : boolean;
  signal slice_234_inst_ack_1 : boolean;
  signal slice_246_inst_ack_1 : boolean;
  signal slice_266_inst_ack_1 : boolean;
  signal slice_238_inst_ack_0 : boolean;
  signal slice_242_inst_ack_0 : boolean;
  signal slice_230_inst_ack_1 : boolean;
  signal slice_222_inst_ack_0 : boolean;
  signal slice_234_inst_req_1 : boolean;
  signal slice_234_inst_ack_0 : boolean;
  signal slice_226_inst_req_1 : boolean;
  signal slice_222_inst_req_0 : boolean;
  signal slice_230_inst_req_1 : boolean;
  signal slice_214_inst_ack_0 : boolean;
  signal slice_378_inst_req_1 : boolean;
  signal slice_214_inst_req_0 : boolean;
  signal slice_242_inst_req_0 : boolean;
  signal slice_238_inst_req_0 : boolean;
  signal slice_246_inst_req_1 : boolean;
  signal W_myptr5_1040_delayed_8_0_1040_inst_ack_0 : boolean;
  signal slice_370_inst_req_0 : boolean;
  signal slice_230_inst_ack_0 : boolean;
  signal slice_226_inst_ack_0 : boolean;
  signal W_myptr5_1040_delayed_8_0_1040_inst_req_1 : boolean;
  signal slice_230_inst_req_0 : boolean;
  signal slice_254_inst_ack_0 : boolean;
  signal slice_250_inst_ack_1 : boolean;
  signal slice_258_inst_ack_1 : boolean;
  signal slice_258_inst_req_1 : boolean;
  signal slice_378_inst_ack_1 : boolean;
  signal slice_234_inst_req_0 : boolean;
  signal slice_266_inst_req_1 : boolean;
  signal slice_250_inst_req_1 : boolean;
  signal W_myptr5_1040_delayed_8_0_1040_inst_req_0 : boolean;
  signal slice_226_inst_req_0 : boolean;
  signal slice_210_inst_ack_0 : boolean;
  signal slice_250_inst_ack_0 : boolean;
  signal slice_270_inst_req_1 : boolean;
  signal slice_210_inst_req_0 : boolean;
  signal slice_218_inst_ack_1 : boolean;
  signal slice_262_inst_ack_1 : boolean;
  signal slice_218_inst_req_1 : boolean;
  signal slice_390_inst_req_1 : boolean;
  signal addr_of_1064_final_reg_req_0 : boolean;
  signal slice_266_inst_req_0 : boolean;
  signal slice_218_inst_ack_0 : boolean;
  signal slice_218_inst_req_0 : boolean;
  signal slice_262_inst_ack_0 : boolean;
  signal CONCAT_u32_u64_1081_inst_req_0 : boolean;
  signal slice_254_inst_ack_1 : boolean;
  signal slice_258_inst_ack_0 : boolean;
  signal slice_210_inst_ack_1 : boolean;
  signal slice_210_inst_req_1 : boolean;
  signal slice_270_inst_req_0 : boolean;
  signal slice_270_inst_ack_0 : boolean;
  signal slice_254_inst_req_0 : boolean;
  signal slice_250_inst_req_0 : boolean;
  signal ptr_deref_121_load_0_req_0 : boolean;
  signal ptr_deref_121_load_0_ack_0 : boolean;
  signal slice_262_inst_req_0 : boolean;
  signal slice_366_inst_ack_1 : boolean;
  signal slice_262_inst_req_1 : boolean;
  signal slice_238_inst_ack_1 : boolean;
  signal W_myptr5_1040_delayed_8_0_1040_inst_ack_1 : boolean;
  signal slice_206_inst_ack_1 : boolean;
  signal slice_222_inst_ack_1 : boolean;
  signal slice_206_inst_req_1 : boolean;
  signal slice_222_inst_req_1 : boolean;
  signal slice_370_inst_ack_0 : boolean;
  signal slice_214_inst_ack_1 : boolean;
  signal slice_214_inst_req_1 : boolean;
  signal slice_258_inst_req_0 : boolean;
  signal slice_366_inst_req_1 : boolean;
  signal slice_390_inst_ack_1 : boolean;
  signal addr_of_1064_final_reg_ack_0 : boolean;
  signal slice_254_inst_req_1 : boolean;
  signal slice_226_inst_ack_1 : boolean;
  signal slice_382_inst_req_0 : boolean;
  signal slice_370_inst_req_1 : boolean;
  signal array_obj_ref_95_index_offset_req_0 : boolean;
  signal array_obj_ref_95_index_offset_ack_0 : boolean;
  signal array_obj_ref_95_index_offset_req_1 : boolean;
  signal array_obj_ref_95_index_offset_ack_1 : boolean;
  signal addr_of_96_final_reg_req_0 : boolean;
  signal addr_of_96_final_reg_ack_0 : boolean;
  signal slice_370_inst_ack_1 : boolean;
  signal addr_of_96_final_reg_req_1 : boolean;
  signal addr_of_96_final_reg_ack_1 : boolean;
  signal array_obj_ref_102_index_offset_req_0 : boolean;
  signal array_obj_ref_102_index_offset_ack_0 : boolean;
  signal array_obj_ref_102_index_offset_req_1 : boolean;
  signal array_obj_ref_102_index_offset_ack_1 : boolean;
  signal addr_of_103_final_reg_req_0 : boolean;
  signal addr_of_103_final_reg_ack_0 : boolean;
  signal addr_of_103_final_reg_req_1 : boolean;
  signal addr_of_103_final_reg_ack_1 : boolean;
  signal array_obj_ref_109_index_offset_req_0 : boolean;
  signal array_obj_ref_109_index_offset_ack_0 : boolean;
  signal ptr_deref_1044_store_0_req_0 : boolean;
  signal array_obj_ref_109_index_offset_req_1 : boolean;
  signal array_obj_ref_109_index_offset_ack_1 : boolean;
  signal CONCAT_u32_u64_1081_inst_ack_0 : boolean;
  signal slice_374_inst_req_0 : boolean;
  signal addr_of_110_final_reg_req_0 : boolean;
  signal addr_of_110_final_reg_ack_0 : boolean;
  signal addr_of_110_final_reg_req_1 : boolean;
  signal addr_of_110_final_reg_ack_1 : boolean;
  signal slice_374_inst_ack_0 : boolean;
  signal array_obj_ref_1037_index_offset_req_0 : boolean;
  signal array_obj_ref_1037_index_offset_ack_0 : boolean;
  signal array_obj_ref_1063_index_offset_req_0 : boolean;
  signal ptr_deref_1044_store_0_ack_0 : boolean;
  signal array_obj_ref_116_index_offset_req_0 : boolean;
  signal array_obj_ref_116_index_offset_ack_0 : boolean;
  signal array_obj_ref_1037_index_offset_req_1 : boolean;
  signal array_obj_ref_116_index_offset_req_1 : boolean;
  signal array_obj_ref_116_index_offset_ack_1 : boolean;
  signal W_myptr6_1063_delayed_8_0_1066_inst_req_0 : boolean;
  signal array_obj_ref_1037_index_offset_ack_1 : boolean;
  signal addr_of_117_final_reg_req_0 : boolean;
  signal array_obj_ref_1063_index_offset_ack_0 : boolean;
  signal addr_of_117_final_reg_ack_0 : boolean;
  signal addr_of_1064_final_reg_req_1 : boolean;
  signal addr_of_117_final_reg_req_1 : boolean;
  signal addr_of_117_final_reg_ack_1 : boolean;
  signal ptr_deref_121_load_0_req_1 : boolean;
  signal ptr_deref_121_load_0_ack_1 : boolean;
  signal CONCAT_u32_u64_1055_inst_req_0 : boolean;
  signal ptr_deref_125_load_0_req_0 : boolean;
  signal ptr_deref_125_load_0_ack_0 : boolean;
  signal slice_374_inst_req_1 : boolean;
  signal CONCAT_u32_u64_1055_inst_ack_0 : boolean;
  signal ptr_deref_125_load_0_req_1 : boolean;
  signal ptr_deref_125_load_0_ack_1 : boolean;
  signal addr_of_1038_final_reg_req_0 : boolean;
  signal slice_374_inst_ack_1 : boolean;
  signal addr_of_1038_final_reg_ack_0 : boolean;
  signal ptr_deref_1044_store_0_req_1 : boolean;
  signal ptr_deref_129_load_0_req_0 : boolean;
  signal ptr_deref_129_load_0_ack_0 : boolean;
  signal CONCAT_u32_u64_1055_inst_req_1 : boolean;
  signal ptr_deref_129_load_0_req_1 : boolean;
  signal ptr_deref_129_load_0_ack_1 : boolean;
  signal W_myptr6_1063_delayed_8_0_1066_inst_ack_0 : boolean;
  signal slice_378_inst_req_0 : boolean;
  signal addr_of_1038_final_reg_req_1 : boolean;
  signal addr_of_1038_final_reg_ack_1 : boolean;
  signal array_obj_ref_1063_index_offset_req_1 : boolean;
  signal CONCAT_u32_u64_1055_inst_ack_1 : boolean;
  signal ptr_deref_1044_store_0_ack_1 : boolean;
  signal ptr_deref_133_load_0_req_0 : boolean;
  signal ptr_deref_133_load_0_ack_0 : boolean;
  signal array_obj_ref_1063_index_offset_ack_1 : boolean;
  signal ptr_deref_133_load_0_req_1 : boolean;
  signal ptr_deref_133_load_0_ack_1 : boolean;
  signal slice_138_inst_req_0 : boolean;
  signal slice_138_inst_ack_0 : boolean;
  signal slice_138_inst_req_1 : boolean;
  signal slice_138_inst_ack_1 : boolean;
  signal slice_142_inst_req_0 : boolean;
  signal slice_142_inst_ack_0 : boolean;
  signal slice_142_inst_req_1 : boolean;
  signal slice_142_inst_ack_1 : boolean;
  signal slice_146_inst_req_0 : boolean;
  signal slice_146_inst_ack_0 : boolean;
  signal slice_146_inst_req_1 : boolean;
  signal slice_146_inst_ack_1 : boolean;
  signal slice_150_inst_req_0 : boolean;
  signal slice_150_inst_ack_0 : boolean;
  signal slice_150_inst_req_1 : boolean;
  signal slice_150_inst_ack_1 : boolean;
  signal slice_154_inst_req_0 : boolean;
  signal slice_154_inst_ack_0 : boolean;
  signal slice_154_inst_req_1 : boolean;
  signal slice_154_inst_ack_1 : boolean;
  signal slice_158_inst_req_0 : boolean;
  signal slice_158_inst_ack_0 : boolean;
  signal slice_158_inst_req_1 : boolean;
  signal slice_158_inst_ack_1 : boolean;
  signal slice_162_inst_req_0 : boolean;
  signal slice_162_inst_ack_0 : boolean;
  signal slice_162_inst_req_1 : boolean;
  signal slice_162_inst_ack_1 : boolean;
  signal slice_166_inst_req_0 : boolean;
  signal slice_166_inst_ack_0 : boolean;
  signal slice_166_inst_req_1 : boolean;
  signal slice_166_inst_ack_1 : boolean;
  signal slice_170_inst_req_0 : boolean;
  signal slice_170_inst_ack_0 : boolean;
  signal slice_170_inst_req_1 : boolean;
  signal slice_170_inst_ack_1 : boolean;
  signal slice_174_inst_req_0 : boolean;
  signal slice_174_inst_ack_0 : boolean;
  signal slice_174_inst_req_1 : boolean;
  signal slice_174_inst_ack_1 : boolean;
  signal slice_178_inst_req_0 : boolean;
  signal slice_178_inst_ack_0 : boolean;
  signal slice_178_inst_req_1 : boolean;
  signal slice_178_inst_ack_1 : boolean;
  signal slice_182_inst_req_0 : boolean;
  signal slice_182_inst_ack_0 : boolean;
  signal slice_182_inst_req_1 : boolean;
  signal slice_182_inst_ack_1 : boolean;
  signal slice_186_inst_req_0 : boolean;
  signal slice_186_inst_ack_0 : boolean;
  signal slice_186_inst_req_1 : boolean;
  signal slice_186_inst_ack_1 : boolean;
  signal slice_190_inst_req_0 : boolean;
  signal slice_190_inst_ack_0 : boolean;
  signal slice_190_inst_req_1 : boolean;
  signal slice_190_inst_ack_1 : boolean;
  signal slice_194_inst_req_0 : boolean;
  signal slice_194_inst_ack_0 : boolean;
  signal slice_194_inst_req_1 : boolean;
  signal slice_194_inst_ack_1 : boolean;
  signal slice_198_inst_req_0 : boolean;
  signal slice_198_inst_ack_0 : boolean;
  signal slice_198_inst_req_1 : boolean;
  signal slice_198_inst_ack_1 : boolean;
  signal slice_202_inst_req_0 : boolean;
  signal slice_202_inst_ack_0 : boolean;
  signal slice_202_inst_req_1 : boolean;
  signal slice_202_inst_ack_1 : boolean;
  signal slice_206_inst_req_0 : boolean;
  signal slice_206_inst_ack_0 : boolean;
  signal ptr_deref_1070_store_0_req_1 : boolean;
  signal ptr_deref_1070_store_0_ack_1 : boolean;
  signal slice_274_inst_req_0 : boolean;
  signal slice_274_inst_ack_0 : boolean;
  signal slice_274_inst_req_1 : boolean;
  signal slice_274_inst_ack_1 : boolean;
  signal slice_390_inst_ack_0 : boolean;
  signal slice_366_inst_ack_0 : boolean;
  signal slice_390_inst_req_0 : boolean;
  signal slice_278_inst_req_0 : boolean;
  signal slice_278_inst_ack_0 : boolean;
  signal slice_278_inst_req_1 : boolean;
  signal slice_278_inst_ack_1 : boolean;
  signal ptr_deref_1070_store_0_ack_0 : boolean;
  signal slice_366_inst_req_0 : boolean;
  signal slice_282_inst_req_0 : boolean;
  signal slice_282_inst_ack_0 : boolean;
  signal slice_282_inst_req_1 : boolean;
  signal slice_282_inst_ack_1 : boolean;
  signal ptr_deref_1070_store_0_req_0 : boolean;
  signal slice_286_inst_req_0 : boolean;
  signal slice_286_inst_ack_0 : boolean;
  signal slice_286_inst_req_1 : boolean;
  signal slice_286_inst_ack_1 : boolean;
  signal slice_290_inst_req_0 : boolean;
  signal slice_290_inst_ack_0 : boolean;
  signal slice_290_inst_req_1 : boolean;
  signal slice_290_inst_ack_1 : boolean;
  signal slice_386_inst_ack_1 : boolean;
  signal CONCAT_u32_u64_1081_inst_ack_1 : boolean;
  signal slice_386_inst_req_1 : boolean;
  signal slice_294_inst_req_0 : boolean;
  signal slice_294_inst_ack_0 : boolean;
  signal slice_294_inst_req_1 : boolean;
  signal slice_294_inst_ack_1 : boolean;
  signal slice_298_inst_req_0 : boolean;
  signal slice_298_inst_ack_0 : boolean;
  signal slice_298_inst_req_1 : boolean;
  signal slice_298_inst_ack_1 : boolean;
  signal slice_386_inst_ack_0 : boolean;
  signal slice_386_inst_req_0 : boolean;
  signal slice_302_inst_req_0 : boolean;
  signal slice_302_inst_ack_0 : boolean;
  signal slice_302_inst_req_1 : boolean;
  signal slice_302_inst_ack_1 : boolean;
  signal CONCAT_u32_u64_1081_inst_req_1 : boolean;
  signal slice_306_inst_req_0 : boolean;
  signal slice_306_inst_ack_0 : boolean;
  signal W_myptr6_1063_delayed_8_0_1066_inst_ack_1 : boolean;
  signal slice_306_inst_req_1 : boolean;
  signal slice_306_inst_ack_1 : boolean;
  signal slice_362_inst_ack_1 : boolean;
  signal slice_362_inst_req_1 : boolean;
  signal W_myptr6_1063_delayed_8_0_1066_inst_req_1 : boolean;
  signal slice_310_inst_req_0 : boolean;
  signal slice_310_inst_ack_0 : boolean;
  signal slice_310_inst_req_1 : boolean;
  signal slice_310_inst_ack_1 : boolean;
  signal slice_382_inst_ack_1 : boolean;
  signal slice_362_inst_ack_0 : boolean;
  signal slice_382_inst_req_1 : boolean;
  signal slice_314_inst_req_0 : boolean;
  signal slice_314_inst_ack_0 : boolean;
  signal slice_362_inst_req_0 : boolean;
  signal slice_314_inst_req_1 : boolean;
  signal slice_314_inst_ack_1 : boolean;
  signal addr_of_1064_final_reg_ack_1 : boolean;
  signal slice_382_inst_ack_0 : boolean;
  signal slice_318_inst_req_0 : boolean;
  signal slice_318_inst_ack_0 : boolean;
  signal slice_378_inst_ack_0 : boolean;
  signal slice_318_inst_req_1 : boolean;
  signal slice_318_inst_ack_1 : boolean;
  signal slice_322_inst_req_0 : boolean;
  signal slice_322_inst_ack_0 : boolean;
  signal slice_322_inst_req_1 : boolean;
  signal slice_322_inst_ack_1 : boolean;
  signal slice_326_inst_req_0 : boolean;
  signal slice_326_inst_ack_0 : boolean;
  signal slice_326_inst_req_1 : boolean;
  signal slice_326_inst_ack_1 : boolean;
  signal slice_330_inst_req_0 : boolean;
  signal slice_330_inst_ack_0 : boolean;
  signal slice_330_inst_req_1 : boolean;
  signal slice_330_inst_ack_1 : boolean;
  signal slice_334_inst_req_0 : boolean;
  signal slice_334_inst_ack_0 : boolean;
  signal slice_334_inst_req_1 : boolean;
  signal slice_334_inst_ack_1 : boolean;
  signal slice_338_inst_req_0 : boolean;
  signal slice_338_inst_ack_0 : boolean;
  signal slice_338_inst_req_1 : boolean;
  signal slice_338_inst_ack_1 : boolean;
  signal slice_342_inst_req_0 : boolean;
  signal slice_342_inst_ack_0 : boolean;
  signal slice_342_inst_req_1 : boolean;
  signal slice_342_inst_ack_1 : boolean;
  signal slice_346_inst_req_0 : boolean;
  signal slice_346_inst_ack_0 : boolean;
  signal slice_346_inst_req_1 : boolean;
  signal slice_346_inst_ack_1 : boolean;
  signal slice_350_inst_req_0 : boolean;
  signal slice_350_inst_ack_0 : boolean;
  signal slice_350_inst_req_1 : boolean;
  signal slice_350_inst_ack_1 : boolean;
  signal slice_354_inst_req_0 : boolean;
  signal slice_354_inst_ack_0 : boolean;
  signal slice_354_inst_req_1 : boolean;
  signal slice_354_inst_ack_1 : boolean;
  signal slice_358_inst_req_0 : boolean;
  signal slice_358_inst_ack_0 : boolean;
  signal slice_358_inst_req_1 : boolean;
  signal slice_358_inst_ack_1 : boolean;
  signal array_obj_ref_1089_index_offset_req_0 : boolean;
  signal array_obj_ref_1089_index_offset_ack_0 : boolean;
  signal array_obj_ref_1089_index_offset_req_1 : boolean;
  signal array_obj_ref_1089_index_offset_ack_1 : boolean;
  signal addr_of_1090_final_reg_req_0 : boolean;
  signal addr_of_1090_final_reg_ack_0 : boolean;
  signal addr_of_1090_final_reg_req_1 : boolean;
  signal addr_of_1090_final_reg_ack_1 : boolean;
  signal W_myptr7_1086_delayed_8_0_1092_inst_req_0 : boolean;
  signal W_myptr7_1086_delayed_8_0_1092_inst_ack_0 : boolean;
  signal W_myptr7_1086_delayed_8_0_1092_inst_req_1 : boolean;
  signal W_myptr7_1086_delayed_8_0_1092_inst_ack_1 : boolean;
  signal CONCAT_u32_u64_1107_inst_req_0 : boolean;
  signal CONCAT_u32_u64_1107_inst_ack_0 : boolean;
  signal CONCAT_u32_u64_1107_inst_req_1 : boolean;
  signal CONCAT_u32_u64_1107_inst_ack_1 : boolean;
  signal ptr_deref_1096_store_0_req_0 : boolean;
  signal ptr_deref_1096_store_0_ack_0 : boolean;
  signal ptr_deref_1096_store_0_req_1 : boolean;
  signal ptr_deref_1096_store_0_ack_1 : boolean;
  signal array_obj_ref_1115_index_offset_req_0 : boolean;
  signal array_obj_ref_1115_index_offset_ack_0 : boolean;
  signal array_obj_ref_1115_index_offset_req_1 : boolean;
  signal array_obj_ref_1115_index_offset_ack_1 : boolean;
  signal addr_of_1116_final_reg_req_0 : boolean;
  signal addr_of_1116_final_reg_ack_0 : boolean;
  signal addr_of_1116_final_reg_req_1 : boolean;
  signal addr_of_1116_final_reg_ack_1 : boolean;
  signal W_myptr8_1109_delayed_8_0_1118_inst_req_0 : boolean;
  signal W_myptr8_1109_delayed_8_0_1118_inst_ack_0 : boolean;
  signal W_myptr8_1109_delayed_8_0_1118_inst_req_1 : boolean;
  signal W_myptr8_1109_delayed_8_0_1118_inst_ack_1 : boolean;
  signal CONCAT_u32_u64_1133_inst_req_0 : boolean;
  signal CONCAT_u32_u64_1133_inst_ack_0 : boolean;
  signal CONCAT_u32_u64_1133_inst_req_1 : boolean;
  signal CONCAT_u32_u64_1133_inst_ack_1 : boolean;
  signal ptr_deref_1122_store_0_req_0 : boolean;
  signal ptr_deref_1122_store_0_ack_0 : boolean;
  signal ptr_deref_1122_store_0_req_1 : boolean;
  signal ptr_deref_1122_store_0_ack_1 : boolean;
  signal type_cast_1137_inst_req_0 : boolean;
  signal type_cast_1137_inst_ack_0 : boolean;
  signal type_cast_1137_inst_req_1 : boolean;
  signal type_cast_1137_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "maxPool4_input_buffer", -- 
      buffer_size => 2,
      bypass_flag => false,
      data_width => tag_length + 160) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(31 downto 0) <= addr;
  addr_buffer <= in_buffer_data_out(31 downto 0);
  in_buffer_data_in(63 downto 32) <= addr1;
  addr1_buffer <= in_buffer_data_out(63 downto 32);
  in_buffer_data_in(95 downto 64) <= addr2;
  addr2_buffer <= in_buffer_data_out(95 downto 64);
  in_buffer_data_in(127 downto 96) <= addr3;
  addr3_buffer <= in_buffer_data_out(127 downto 96);
  in_buffer_data_in(159 downto 128) <= addr4;
  addr4_buffer <= in_buffer_data_out(159 downto 128);
  in_buffer_data_in(tag_length + 159 downto 160) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 159 downto 160);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 1,6 => 15);
    constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1,6 => 15);
    constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 7); -- 
  begin -- 
    preds <= addr_update_enable & addr1_update_enable & addr2_update_enable & addr3_update_enable & addr4_update_enable & in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  maxPool4_CP_346_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "maxPool4_out_buffer", -- 
      buffer_size => 2,
      full_rate => false,
      data_width => tag_length + 8) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(7 downto 0) <= output_buffer;
  output <= out_buffer_data_out(7 downto 0);
  out_buffer_data_in(tag_length + 7 downto 8) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 7 downto 8);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 15);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= maxPool4_CP_346_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  output_update_enable_join: block -- 
    constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
    constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
    constant place_delays: IntegerArray(0 to 0) := (0 => 0);
    constant joinName: string(1 to 25) := "output_update_enable_join"; 
    signal preds: BooleanArray(1 to 1); -- 
  begin -- 
    preds(1) <= out_buffer_write_ack_symbol;
    gj_output_update_enable_join : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => output_update_enable, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 15,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= maxPool4_CP_346_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= maxPool4_CP_346_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  maxPool4_CP_346: Block -- control-path 
    signal maxPool4_CP_346_elements: BooleanArray(398 downto 0);
    -- 
  begin -- 
    maxPool4_CP_346_elements(0) <= maxPool4_CP_346_start;
    maxPool4_CP_346_symbol <= maxPool4_CP_346_elements(398);
    -- CP-element group 0:  transition  bypass  pipeline-parent 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (1) 
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	10 
    -- CP-element group 1: 	11 
    -- CP-element group 1: 	9 
    -- CP-element group 1: 	16 
    -- CP-element group 1: 	17 
    -- CP-element group 1: 	18 
    -- CP-element group 1: 	23 
    -- CP-element group 1: 	24 
    -- CP-element group 1: 	25 
    -- CP-element group 1: 	30 
    -- CP-element group 1: 	31 
    -- CP-element group 1: 	32 
    -- CP-element group 1: 	309 
    -- CP-element group 1: 	310 
    -- CP-element group 1: 	311 
    -- CP-element group 1: 	328 
    -- CP-element group 1: 	329 
    -- CP-element group 1: 	330 
    -- CP-element group 1: 	347 
    -- CP-element group 1: 	348 
    -- CP-element group 1: 	349 
    -- CP-element group 1: 	366 
    -- CP-element group 1: 	367 
    -- CP-element group 1: 	368 
    -- CP-element group 1:  members (105) 
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1063_index_scale_1/scale_rename_req
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1063_index_scale_1/scale_rename_ack
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1037_index_resize_1/$entry
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1063_index_scale_1/$exit
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1037_index_resize_1/$exit
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1037_index_resized_1
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1037_index_scaled_1
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1037_index_computed_1
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1037_index_resize_1/index_resize_req
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1063_index_scale_1/$entry
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/$entry
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_95_index_resized_1
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_95_index_scaled_1
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_95_index_computed_1
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_95_index_resize_1/$entry
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_95_index_resize_1/$exit
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_95_index_resize_1/index_resize_req
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_95_index_resize_1/index_resize_ack
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1037_index_resize_1/index_resize_ack
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_95_index_scale_1/$entry
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_95_index_scale_1/$exit
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_95_index_scale_1/scale_rename_req
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_95_index_scale_1/scale_rename_ack
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_95_final_index_sum_regn_Sample/$entry
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_95_final_index_sum_regn_Sample/req
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1037_index_scale_1/$entry
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1037_index_scale_1/$exit
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1037_index_scale_1/scale_rename_req
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_102_index_resized_1
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_102_index_scaled_1
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_102_index_computed_1
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_102_index_resize_1/$entry
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_102_index_resize_1/$exit
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_102_index_resize_1/index_resize_req
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_102_index_resize_1/index_resize_ack
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_102_index_scale_1/$entry
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_102_index_scale_1/$exit
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_102_index_scale_1/scale_rename_req
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_102_index_scale_1/scale_rename_ack
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_102_final_index_sum_regn_Sample/$entry
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_102_final_index_sum_regn_Sample/req
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1063_final_index_sum_regn_Sample/$entry
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1037_index_scale_1/scale_rename_ack
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_109_index_resized_1
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_109_index_scaled_1
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_109_index_computed_1
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_109_index_resize_1/$entry
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_109_index_resize_1/$exit
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_109_index_resize_1/index_resize_req
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_109_index_resize_1/index_resize_ack
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_109_index_scale_1/$entry
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_109_index_scale_1/$exit
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_109_index_scale_1/scale_rename_req
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_109_index_scale_1/scale_rename_ack
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_109_final_index_sum_regn_Sample/$entry
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_109_final_index_sum_regn_Sample/req
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1037_final_index_sum_regn_Sample/$entry
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1037_final_index_sum_regn_Sample/req
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_116_index_resized_1
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_116_index_scaled_1
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_116_index_computed_1
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_116_index_resize_1/$entry
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_116_index_resize_1/$exit
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_116_index_resize_1/index_resize_req
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_116_index_resize_1/index_resize_ack
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1063_final_index_sum_regn_Sample/req
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_116_index_scale_1/$entry
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_116_index_scale_1/$exit
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_116_index_scale_1/scale_rename_req
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_116_index_scale_1/scale_rename_ack
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_116_final_index_sum_regn_Sample/$entry
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_116_final_index_sum_regn_Sample/req
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1063_index_resize_1/index_resize_ack
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1063_index_resize_1/index_resize_req
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1063_index_resize_1/$exit
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1063_index_resize_1/$entry
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1063_index_computed_1
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1063_index_scaled_1
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1063_index_resized_1
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1089_index_resized_1
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1089_index_scaled_1
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1089_index_computed_1
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1089_index_resize_1/$entry
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1089_index_resize_1/$exit
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1089_index_resize_1/index_resize_req
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1089_index_resize_1/index_resize_ack
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1089_index_scale_1/$entry
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1089_index_scale_1/$exit
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1089_index_scale_1/scale_rename_req
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1089_index_scale_1/scale_rename_ack
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1089_final_index_sum_regn_Sample/$entry
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1089_final_index_sum_regn_Sample/req
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1115_index_resized_1
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1115_index_scaled_1
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1115_index_computed_1
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1115_index_resize_1/$entry
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1115_index_resize_1/$exit
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1115_index_resize_1/index_resize_req
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1115_index_resize_1/index_resize_ack
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1115_index_scale_1/$entry
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1115_index_scale_1/$exit
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1115_index_scale_1/scale_rename_req
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1115_index_scale_1/scale_rename_ack
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1115_final_index_sum_regn_Sample/$entry
      -- CP-element group 1: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1115_final_index_sum_regn_Sample/req
      -- 
    req_388_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_388_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(1), ack => array_obj_ref_95_index_offset_req_0); -- 
    req_434_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_434_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(1), ack => array_obj_ref_102_index_offset_req_0); -- 
    req_480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(1), ack => array_obj_ref_109_index_offset_req_0); -- 
    req_526_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_526_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(1), ack => array_obj_ref_116_index_offset_req_0); -- 
    req_1668_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1668_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(1), ack => array_obj_ref_1037_index_offset_req_0); -- 
    req_1792_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1792_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(1), ack => array_obj_ref_1063_index_offset_req_0); -- 
    req_1916_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1916_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(1), ack => array_obj_ref_1089_index_offset_req_0); -- 
    req_2040_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2040_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(1), ack => array_obj_ref_1115_index_offset_req_0); -- 
    maxPool4_CP_346_elements(1) <= maxPool4_CP_346_elements(0);
    -- CP-element group 2:  join  transition  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: marked-predecessors 
    -- CP-element group 2: 	311 
    -- CP-element group 2: 	330 
    -- CP-element group 2: 	349 
    -- CP-element group 2: 	368 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	392 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 assign_stmt_97_to_assign_stmt_1138/addr_update_enable
      -- CP-element group 2: 	 assign_stmt_97_to_assign_stmt_1138/addr_update_enable_out
      -- 
    maxPool4_cp_element_group_2: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant joinName: string(1 to 27) := "maxPool4_cp_element_group_2"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(311) & maxPool4_CP_346_elements(330) & maxPool4_CP_346_elements(349) & maxPool4_CP_346_elements(368);
      gj_maxPool4_cp_element_group_2 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(2), clk => clk, reset => reset); --
    end block;
    -- CP-element group 3:  join  transition  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: marked-predecessors 
    -- CP-element group 3: 	11 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	393 
    -- CP-element group 3:  members (2) 
      -- CP-element group 3: 	 assign_stmt_97_to_assign_stmt_1138/addr1_update_enable
      -- CP-element group 3: 	 assign_stmt_97_to_assign_stmt_1138/addr1_update_enable_out
      -- 
    maxPool4_cp_element_group_3: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 1);
      constant joinName: string(1 to 27) := "maxPool4_cp_element_group_3"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= maxPool4_CP_346_elements(11);
      gj_maxPool4_cp_element_group_3 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(3), clk => clk, reset => reset); --
    end block;
    -- CP-element group 4:  join  transition  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: marked-predecessors 
    -- CP-element group 4: 	18 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	394 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 assign_stmt_97_to_assign_stmt_1138/addr2_update_enable
      -- CP-element group 4: 	 assign_stmt_97_to_assign_stmt_1138/addr2_update_enable_out
      -- 
    maxPool4_cp_element_group_4: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 1);
      constant joinName: string(1 to 27) := "maxPool4_cp_element_group_4"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= maxPool4_CP_346_elements(18);
      gj_maxPool4_cp_element_group_4 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(4), clk => clk, reset => reset); --
    end block;
    -- CP-element group 5:  join  transition  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: marked-predecessors 
    -- CP-element group 5: 	25 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	395 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 assign_stmt_97_to_assign_stmt_1138/addr3_update_enable
      -- CP-element group 5: 	 assign_stmt_97_to_assign_stmt_1138/addr3_update_enable_out
      -- 
    maxPool4_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 1);
      constant joinName: string(1 to 27) := "maxPool4_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= maxPool4_CP_346_elements(25);
      gj_maxPool4_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(5), clk => clk, reset => reset); --
    end block;
    -- CP-element group 6:  join  transition  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: marked-predecessors 
    -- CP-element group 6: 	32 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	396 
    -- CP-element group 6:  members (2) 
      -- CP-element group 6: 	 assign_stmt_97_to_assign_stmt_1138/addr4_update_enable
      -- CP-element group 6: 	 assign_stmt_97_to_assign_stmt_1138/addr4_update_enable_out
      -- 
    maxPool4_cp_element_group_6: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 1);
      constant joinName: string(1 to 27) := "maxPool4_cp_element_group_6"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= maxPool4_CP_346_elements(32);
      gj_maxPool4_cp_element_group_6 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(6), clk => clk, reset => reset); --
    end block;
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	397 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	385 
    -- CP-element group 7:  members (2) 
      -- CP-element group 7: 	 assign_stmt_97_to_assign_stmt_1138/output_update_enable
      -- CP-element group 7: 	 assign_stmt_97_to_assign_stmt_1138/output_update_enable_in
      -- 
    maxPool4_CP_346_elements(7) <= maxPool4_CP_346_elements(397);
    -- CP-element group 8:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	12 
    -- CP-element group 8: marked-predecessors 
    -- CP-element group 8: 	13 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	13 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_96_sample_start_
      -- CP-element group 8: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_96_request/$entry
      -- CP-element group 8: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_96_request/req
      -- 
    req_403_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_403_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(8), ack => addr_of_96_final_reg_req_0); -- 
    maxPool4_cp_element_group_8: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 27) := "maxPool4_cp_element_group_8"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(12) & maxPool4_CP_346_elements(13);
      gj_maxPool4_cp_element_group_8 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(8), clk => clk, reset => reset); --
    end block;
    -- CP-element group 9:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	1 
    -- CP-element group 9: marked-predecessors 
    -- CP-element group 9: 	38 
    -- CP-element group 9: 	14 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	14 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_96_update_start_
      -- CP-element group 9: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_96_complete/$entry
      -- CP-element group 9: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_96_complete/req
      -- 
    req_408_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_408_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(9), ack => addr_of_96_final_reg_req_1); -- 
    maxPool4_cp_element_group_9: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 27) := "maxPool4_cp_element_group_9"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(1) & maxPool4_CP_346_elements(38) & maxPool4_CP_346_elements(14);
      gj_maxPool4_cp_element_group_9 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(9), clk => clk, reset => reset); --
    end block;
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	1 
    -- CP-element group 10: marked-predecessors 
    -- CP-element group 10: 	12 
    -- CP-element group 10: 	13 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	12 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_95_final_index_sum_regn_update_start
      -- CP-element group 10: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_95_final_index_sum_regn_Update/$entry
      -- CP-element group 10: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_95_final_index_sum_regn_Update/req
      -- 
    req_393_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_393_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(10), ack => array_obj_ref_95_index_offset_req_1); -- 
    maxPool4_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(1) & maxPool4_CP_346_elements(12) & maxPool4_CP_346_elements(13);
      gj_maxPool4_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	1 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	391 
    -- CP-element group 11: marked-successors 
    -- CP-element group 11: 	3 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_95_final_index_sum_regn_sample_complete
      -- CP-element group 11: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_95_final_index_sum_regn_Sample/$exit
      -- CP-element group 11: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_95_final_index_sum_regn_Sample/ack
      -- 
    ack_389_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_95_index_offset_ack_0, ack => maxPool4_CP_346_elements(11)); -- 
    -- CP-element group 12:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	10 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	8 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	10 
    -- CP-element group 12:  members (8) 
      -- CP-element group 12: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_95_root_address_calculated
      -- CP-element group 12: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_95_offset_calculated
      -- CP-element group 12: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_95_final_index_sum_regn_Update/$exit
      -- CP-element group 12: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_95_final_index_sum_regn_Update/ack
      -- CP-element group 12: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_95_base_plus_offset/$entry
      -- CP-element group 12: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_95_base_plus_offset/$exit
      -- CP-element group 12: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_95_base_plus_offset/sum_rename_req
      -- CP-element group 12: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_95_base_plus_offset/sum_rename_ack
      -- 
    ack_394_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_95_index_offset_ack_1, ack => maxPool4_CP_346_elements(12)); -- 
    -- CP-element group 13:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	8 
    -- CP-element group 13: successors 
    -- CP-element group 13: marked-successors 
    -- CP-element group 13: 	10 
    -- CP-element group 13: 	8 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_96_sample_completed_
      -- CP-element group 13: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_96_request/$exit
      -- CP-element group 13: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_96_request/ack
      -- 
    ack_404_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_96_final_reg_ack_0, ack => maxPool4_CP_346_elements(13)); -- 
    -- CP-element group 14:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	9 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	36 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	9 
    -- CP-element group 14:  members (19) 
      -- CP-element group 14: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_121_word_address_calculated
      -- CP-element group 14: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_121_root_address_calculated
      -- CP-element group 14: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_121_base_address_resized
      -- CP-element group 14: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_121_base_addr_resize/$entry
      -- CP-element group 14: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_121_base_addr_resize/$exit
      -- CP-element group 14: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_121_base_addr_resize/base_resize_req
      -- CP-element group 14: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_121_base_addr_resize/base_resize_ack
      -- CP-element group 14: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_121_base_plus_offset/$entry
      -- CP-element group 14: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_121_base_plus_offset/$exit
      -- CP-element group 14: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_121_base_plus_offset/sum_rename_req
      -- CP-element group 14: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_121_base_plus_offset/sum_rename_ack
      -- CP-element group 14: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_121_word_addrgen/$entry
      -- CP-element group 14: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_121_word_addrgen/$exit
      -- CP-element group 14: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_121_word_addrgen/root_register_req
      -- CP-element group 14: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_121_word_addrgen/root_register_ack
      -- CP-element group 14: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_96_update_completed_
      -- CP-element group 14: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_96_complete/$exit
      -- CP-element group 14: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_96_complete/ack
      -- CP-element group 14: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_121_base_address_calculated
      -- 
    ack_409_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_96_final_reg_ack_1, ack => maxPool4_CP_346_elements(14)); -- 
    -- CP-element group 15:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	19 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	20 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	20 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_103_sample_start_
      -- CP-element group 15: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_103_request/$entry
      -- CP-element group 15: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_103_request/req
      -- 
    req_449_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_449_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(15), ack => addr_of_103_final_reg_req_0); -- 
    maxPool4_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(19) & maxPool4_CP_346_elements(20);
      gj_maxPool4_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	1 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	42 
    -- CP-element group 16: 	21 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	21 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_103_update_start_
      -- CP-element group 16: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_103_complete/$entry
      -- CP-element group 16: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_103_complete/req
      -- 
    req_454_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_454_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(16), ack => addr_of_103_final_reg_req_1); -- 
    maxPool4_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(1) & maxPool4_CP_346_elements(42) & maxPool4_CP_346_elements(21);
      gj_maxPool4_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	1 
    -- CP-element group 17: marked-predecessors 
    -- CP-element group 17: 	19 
    -- CP-element group 17: 	20 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	19 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_102_final_index_sum_regn_update_start
      -- CP-element group 17: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_102_final_index_sum_regn_Update/$entry
      -- CP-element group 17: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_102_final_index_sum_regn_Update/req
      -- 
    req_439_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_439_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(17), ack => array_obj_ref_102_index_offset_req_1); -- 
    maxPool4_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(1) & maxPool4_CP_346_elements(19) & maxPool4_CP_346_elements(20);
      gj_maxPool4_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	1 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	391 
    -- CP-element group 18: marked-successors 
    -- CP-element group 18: 	4 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_102_final_index_sum_regn_sample_complete
      -- CP-element group 18: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_102_final_index_sum_regn_Sample/$exit
      -- CP-element group 18: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_102_final_index_sum_regn_Sample/ack
      -- 
    ack_435_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_102_index_offset_ack_0, ack => maxPool4_CP_346_elements(18)); -- 
    -- CP-element group 19:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	17 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	15 
    -- CP-element group 19: marked-successors 
    -- CP-element group 19: 	17 
    -- CP-element group 19:  members (8) 
      -- CP-element group 19: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_102_root_address_calculated
      -- CP-element group 19: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_102_offset_calculated
      -- CP-element group 19: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_102_final_index_sum_regn_Update/$exit
      -- CP-element group 19: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_102_final_index_sum_regn_Update/ack
      -- CP-element group 19: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_102_base_plus_offset/$entry
      -- CP-element group 19: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_102_base_plus_offset/$exit
      -- CP-element group 19: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_102_base_plus_offset/sum_rename_req
      -- CP-element group 19: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_102_base_plus_offset/sum_rename_ack
      -- 
    ack_440_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_102_index_offset_ack_1, ack => maxPool4_CP_346_elements(19)); -- 
    -- CP-element group 20:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	15 
    -- CP-element group 20: successors 
    -- CP-element group 20: marked-successors 
    -- CP-element group 20: 	15 
    -- CP-element group 20: 	17 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_103_sample_completed_
      -- CP-element group 20: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_103_request/$exit
      -- CP-element group 20: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_103_request/ack
      -- 
    ack_450_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_103_final_reg_ack_0, ack => maxPool4_CP_346_elements(20)); -- 
    -- CP-element group 21:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	16 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	40 
    -- CP-element group 21: marked-successors 
    -- CP-element group 21: 	16 
    -- CP-element group 21:  members (19) 
      -- CP-element group 21: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_103_update_completed_
      -- CP-element group 21: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_103_complete/$exit
      -- CP-element group 21: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_103_complete/ack
      -- CP-element group 21: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_125_base_address_calculated
      -- CP-element group 21: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_125_word_address_calculated
      -- CP-element group 21: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_125_root_address_calculated
      -- CP-element group 21: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_125_base_address_resized
      -- CP-element group 21: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_125_base_addr_resize/$entry
      -- CP-element group 21: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_125_base_addr_resize/$exit
      -- CP-element group 21: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_125_base_addr_resize/base_resize_req
      -- CP-element group 21: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_125_base_addr_resize/base_resize_ack
      -- CP-element group 21: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_125_base_plus_offset/$entry
      -- CP-element group 21: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_125_base_plus_offset/$exit
      -- CP-element group 21: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_125_base_plus_offset/sum_rename_req
      -- CP-element group 21: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_125_base_plus_offset/sum_rename_ack
      -- CP-element group 21: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_125_word_addrgen/$entry
      -- CP-element group 21: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_125_word_addrgen/$exit
      -- CP-element group 21: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_125_word_addrgen/root_register_req
      -- CP-element group 21: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_125_word_addrgen/root_register_ack
      -- 
    ack_455_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_103_final_reg_ack_1, ack => maxPool4_CP_346_elements(21)); -- 
    -- CP-element group 22:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	26 
    -- CP-element group 22: marked-predecessors 
    -- CP-element group 22: 	27 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	27 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_110_sample_start_
      -- CP-element group 22: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_110_request/$entry
      -- CP-element group 22: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_110_request/req
      -- 
    req_495_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_495_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(22), ack => addr_of_110_final_reg_req_0); -- 
    maxPool4_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(26) & maxPool4_CP_346_elements(27);
      gj_maxPool4_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	1 
    -- CP-element group 23: marked-predecessors 
    -- CP-element group 23: 	46 
    -- CP-element group 23: 	28 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	28 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_110_update_start_
      -- CP-element group 23: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_110_complete/$entry
      -- CP-element group 23: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_110_complete/req
      -- 
    req_500_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_500_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(23), ack => addr_of_110_final_reg_req_1); -- 
    maxPool4_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(1) & maxPool4_CP_346_elements(46) & maxPool4_CP_346_elements(28);
      gj_maxPool4_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	1 
    -- CP-element group 24: marked-predecessors 
    -- CP-element group 24: 	26 
    -- CP-element group 24: 	27 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	26 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_109_final_index_sum_regn_update_start
      -- CP-element group 24: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_109_final_index_sum_regn_Update/$entry
      -- CP-element group 24: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_109_final_index_sum_regn_Update/req
      -- 
    req_485_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_485_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(24), ack => array_obj_ref_109_index_offset_req_1); -- 
    maxPool4_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(1) & maxPool4_CP_346_elements(26) & maxPool4_CP_346_elements(27);
      gj_maxPool4_cp_element_group_24 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(24), clk => clk, reset => reset); --
    end block;
    -- CP-element group 25:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	1 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	391 
    -- CP-element group 25: marked-successors 
    -- CP-element group 25: 	5 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_109_final_index_sum_regn_sample_complete
      -- CP-element group 25: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_109_final_index_sum_regn_Sample/$exit
      -- CP-element group 25: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_109_final_index_sum_regn_Sample/ack
      -- 
    ack_481_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_109_index_offset_ack_0, ack => maxPool4_CP_346_elements(25)); -- 
    -- CP-element group 26:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	22 
    -- CP-element group 26: marked-successors 
    -- CP-element group 26: 	24 
    -- CP-element group 26:  members (8) 
      -- CP-element group 26: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_109_root_address_calculated
      -- CP-element group 26: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_109_offset_calculated
      -- CP-element group 26: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_109_final_index_sum_regn_Update/$exit
      -- CP-element group 26: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_109_final_index_sum_regn_Update/ack
      -- CP-element group 26: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_109_base_plus_offset/$entry
      -- CP-element group 26: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_109_base_plus_offset/$exit
      -- CP-element group 26: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_109_base_plus_offset/sum_rename_req
      -- CP-element group 26: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_109_base_plus_offset/sum_rename_ack
      -- 
    ack_486_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_109_index_offset_ack_1, ack => maxPool4_CP_346_elements(26)); -- 
    -- CP-element group 27:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	22 
    -- CP-element group 27: successors 
    -- CP-element group 27: marked-successors 
    -- CP-element group 27: 	22 
    -- CP-element group 27: 	24 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_110_sample_completed_
      -- CP-element group 27: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_110_request/$exit
      -- CP-element group 27: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_110_request/ack
      -- 
    ack_496_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_110_final_reg_ack_0, ack => maxPool4_CP_346_elements(27)); -- 
    -- CP-element group 28:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	23 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	44 
    -- CP-element group 28: marked-successors 
    -- CP-element group 28: 	23 
    -- CP-element group 28:  members (19) 
      -- CP-element group 28: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_110_update_completed_
      -- CP-element group 28: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_110_complete/$exit
      -- CP-element group 28: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_110_complete/ack
      -- CP-element group 28: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_129_base_address_calculated
      -- CP-element group 28: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_129_word_address_calculated
      -- CP-element group 28: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_129_root_address_calculated
      -- CP-element group 28: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_129_base_address_resized
      -- CP-element group 28: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_129_base_addr_resize/$entry
      -- CP-element group 28: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_129_base_addr_resize/$exit
      -- CP-element group 28: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_129_base_addr_resize/base_resize_req
      -- CP-element group 28: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_129_base_addr_resize/base_resize_ack
      -- CP-element group 28: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_129_base_plus_offset/$entry
      -- CP-element group 28: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_129_base_plus_offset/$exit
      -- CP-element group 28: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_129_base_plus_offset/sum_rename_req
      -- CP-element group 28: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_129_base_plus_offset/sum_rename_ack
      -- CP-element group 28: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_129_word_addrgen/$entry
      -- CP-element group 28: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_129_word_addrgen/$exit
      -- CP-element group 28: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_129_word_addrgen/root_register_req
      -- CP-element group 28: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_129_word_addrgen/root_register_ack
      -- 
    ack_501_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_110_final_reg_ack_1, ack => maxPool4_CP_346_elements(28)); -- 
    -- CP-element group 29:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	33 
    -- CP-element group 29: marked-predecessors 
    -- CP-element group 29: 	34 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	34 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_117_sample_start_
      -- CP-element group 29: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_117_request/$entry
      -- CP-element group 29: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_117_request/req
      -- 
    req_541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(29), ack => addr_of_117_final_reg_req_0); -- 
    maxPool4_cp_element_group_29: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_29"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(33) & maxPool4_CP_346_elements(34);
      gj_maxPool4_cp_element_group_29 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(29), clk => clk, reset => reset); --
    end block;
    -- CP-element group 30:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	1 
    -- CP-element group 30: marked-predecessors 
    -- CP-element group 30: 	35 
    -- CP-element group 30: 	50 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	35 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_117_update_start_
      -- CP-element group 30: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_117_complete/$entry
      -- CP-element group 30: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_117_complete/req
      -- 
    req_546_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_546_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(30), ack => addr_of_117_final_reg_req_1); -- 
    maxPool4_cp_element_group_30: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_30"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(1) & maxPool4_CP_346_elements(35) & maxPool4_CP_346_elements(50);
      gj_maxPool4_cp_element_group_30 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(30), clk => clk, reset => reset); --
    end block;
    -- CP-element group 31:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	1 
    -- CP-element group 31: marked-predecessors 
    -- CP-element group 31: 	34 
    -- CP-element group 31: 	33 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_116_final_index_sum_regn_update_start
      -- CP-element group 31: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_116_final_index_sum_regn_Update/$entry
      -- CP-element group 31: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_116_final_index_sum_regn_Update/req
      -- 
    req_531_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_531_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(31), ack => array_obj_ref_116_index_offset_req_1); -- 
    maxPool4_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(1) & maxPool4_CP_346_elements(34) & maxPool4_CP_346_elements(33);
      gj_maxPool4_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	1 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	391 
    -- CP-element group 32: marked-successors 
    -- CP-element group 32: 	6 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_116_final_index_sum_regn_sample_complete
      -- CP-element group 32: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_116_final_index_sum_regn_Sample/$exit
      -- CP-element group 32: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_116_final_index_sum_regn_Sample/ack
      -- 
    ack_527_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_116_index_offset_ack_0, ack => maxPool4_CP_346_elements(32)); -- 
    -- CP-element group 33:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	29 
    -- CP-element group 33: marked-successors 
    -- CP-element group 33: 	31 
    -- CP-element group 33:  members (8) 
      -- CP-element group 33: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_116_root_address_calculated
      -- CP-element group 33: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_116_offset_calculated
      -- CP-element group 33: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_116_final_index_sum_regn_Update/$exit
      -- CP-element group 33: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_116_final_index_sum_regn_Update/ack
      -- CP-element group 33: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_116_base_plus_offset/$entry
      -- CP-element group 33: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_116_base_plus_offset/$exit
      -- CP-element group 33: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_116_base_plus_offset/sum_rename_req
      -- CP-element group 33: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_116_base_plus_offset/sum_rename_ack
      -- 
    ack_532_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_116_index_offset_ack_1, ack => maxPool4_CP_346_elements(33)); -- 
    -- CP-element group 34:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	29 
    -- CP-element group 34: successors 
    -- CP-element group 34: marked-successors 
    -- CP-element group 34: 	29 
    -- CP-element group 34: 	31 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_117_sample_completed_
      -- CP-element group 34: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_117_request/$exit
      -- CP-element group 34: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_117_request/ack
      -- 
    ack_542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_117_final_reg_ack_0, ack => maxPool4_CP_346_elements(34)); -- 
    -- CP-element group 35:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	30 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	48 
    -- CP-element group 35: marked-successors 
    -- CP-element group 35: 	30 
    -- CP-element group 35:  members (19) 
      -- CP-element group 35: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_133_root_address_calculated
      -- CP-element group 35: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_117_update_completed_
      -- CP-element group 35: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_117_complete/$exit
      -- CP-element group 35: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_117_complete/ack
      -- CP-element group 35: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_133_base_address_calculated
      -- CP-element group 35: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_133_word_address_calculated
      -- CP-element group 35: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_133_base_address_resized
      -- CP-element group 35: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_133_base_addr_resize/$entry
      -- CP-element group 35: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_133_base_addr_resize/$exit
      -- CP-element group 35: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_133_base_addr_resize/base_resize_req
      -- CP-element group 35: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_133_base_addr_resize/base_resize_ack
      -- CP-element group 35: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_133_base_plus_offset/$entry
      -- CP-element group 35: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_133_base_plus_offset/$exit
      -- CP-element group 35: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_133_base_plus_offset/sum_rename_req
      -- CP-element group 35: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_133_base_plus_offset/sum_rename_ack
      -- CP-element group 35: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_133_word_addrgen/$entry
      -- CP-element group 35: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_133_word_addrgen/$exit
      -- CP-element group 35: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_133_word_addrgen/root_register_req
      -- CP-element group 35: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_133_word_addrgen/root_register_ack
      -- 
    ack_547_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_117_final_reg_ack_1, ack => maxPool4_CP_346_elements(35)); -- 
    -- CP-element group 36:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	14 
    -- CP-element group 36: marked-predecessors 
    -- CP-element group 36: 	38 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	38 
    -- CP-element group 36:  members (5) 
      -- CP-element group 36: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_121_Sample/$entry
      -- CP-element group 36: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_121_Sample/word_access_start/$entry
      -- CP-element group 36: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_121_Sample/word_access_start/word_0/$entry
      -- CP-element group 36: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_121_Sample/word_access_start/word_0/rr
      -- CP-element group 36: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_121_sample_start_
      -- 
    rr_580_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_580_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(36), ack => ptr_deref_121_load_0_req_0); -- 
    maxPool4_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(14) & maxPool4_CP_346_elements(38);
      gj_maxPool4_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	39 
    -- CP-element group 37: 	54 
    -- CP-element group 37: 	58 
    -- CP-element group 37: 	62 
    -- CP-element group 37: 	66 
    -- CP-element group 37: 	70 
    -- CP-element group 37: 	74 
    -- CP-element group 37: 	78 
    -- CP-element group 37: 	82 
    -- CP-element group 37: 	86 
    -- CP-element group 37: 	90 
    -- CP-element group 37: 	94 
    -- CP-element group 37: 	98 
    -- CP-element group 37: 	102 
    -- CP-element group 37: 	106 
    -- CP-element group 37: 	110 
    -- CP-element group 37: 	114 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	39 
    -- CP-element group 37:  members (5) 
      -- CP-element group 37: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_121_Update/$entry
      -- CP-element group 37: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_121_update_start_
      -- CP-element group 37: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_121_Update/word_access_complete/$entry
      -- CP-element group 37: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_121_Update/word_access_complete/word_0/$entry
      -- CP-element group 37: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_121_Update/word_access_complete/word_0/cr
      -- 
    cr_591_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_591_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(37), ack => ptr_deref_121_load_0_req_1); -- 
    maxPool4_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 16) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_markings: IntegerArray(0 to 16)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_delays: IntegerArray(0 to 16) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 17); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(39) & maxPool4_CP_346_elements(54) & maxPool4_CP_346_elements(58) & maxPool4_CP_346_elements(62) & maxPool4_CP_346_elements(66) & maxPool4_CP_346_elements(70) & maxPool4_CP_346_elements(74) & maxPool4_CP_346_elements(78) & maxPool4_CP_346_elements(82) & maxPool4_CP_346_elements(86) & maxPool4_CP_346_elements(90) & maxPool4_CP_346_elements(94) & maxPool4_CP_346_elements(98) & maxPool4_CP_346_elements(102) & maxPool4_CP_346_elements(106) & maxPool4_CP_346_elements(110) & maxPool4_CP_346_elements(114);
      gj_maxPool4_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 17, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	36 
    -- CP-element group 38: successors 
    -- CP-element group 38: marked-successors 
    -- CP-element group 38: 	36 
    -- CP-element group 38: 	9 
    -- CP-element group 38:  members (5) 
      -- CP-element group 38: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_121_Sample/$exit
      -- CP-element group 38: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_121_Sample/word_access_start/$exit
      -- CP-element group 38: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_121_Sample/word_access_start/word_0/$exit
      -- CP-element group 38: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_121_Sample/word_access_start/word_0/ra
      -- CP-element group 38: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_121_sample_completed_
      -- 
    ra_581_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_121_load_0_ack_0, ack => maxPool4_CP_346_elements(38)); -- 
    -- CP-element group 39:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	37 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	52 
    -- CP-element group 39: 	56 
    -- CP-element group 39: 	60 
    -- CP-element group 39: 	64 
    -- CP-element group 39: 	68 
    -- CP-element group 39: 	72 
    -- CP-element group 39: 	76 
    -- CP-element group 39: 	80 
    -- CP-element group 39: 	84 
    -- CP-element group 39: 	88 
    -- CP-element group 39: 	92 
    -- CP-element group 39: 	96 
    -- CP-element group 39: 	100 
    -- CP-element group 39: 	104 
    -- CP-element group 39: 	108 
    -- CP-element group 39: 	112 
    -- CP-element group 39: marked-successors 
    -- CP-element group 39: 	37 
    -- CP-element group 39:  members (9) 
      -- CP-element group 39: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_121_Update/$exit
      -- CP-element group 39: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_121_update_completed_
      -- CP-element group 39: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_121_Update/word_access_complete/$exit
      -- CP-element group 39: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_121_Update/word_access_complete/word_0/$exit
      -- CP-element group 39: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_121_Update/word_access_complete/word_0/ca
      -- CP-element group 39: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_121_Update/ptr_deref_121_Merge/$entry
      -- CP-element group 39: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_121_Update/ptr_deref_121_Merge/$exit
      -- CP-element group 39: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_121_Update/ptr_deref_121_Merge/merge_req
      -- CP-element group 39: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_121_Update/ptr_deref_121_Merge/merge_ack
      -- 
    ca_592_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_121_load_0_ack_1, ack => maxPool4_CP_346_elements(39)); -- 
    -- CP-element group 40:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	21 
    -- CP-element group 40: marked-predecessors 
    -- CP-element group 40: 	42 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	42 
    -- CP-element group 40:  members (5) 
      -- CP-element group 40: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_125_sample_start_
      -- CP-element group 40: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_125_Sample/$entry
      -- CP-element group 40: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_125_Sample/word_access_start/$entry
      -- CP-element group 40: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_125_Sample/word_access_start/word_0/$entry
      -- CP-element group 40: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_125_Sample/word_access_start/word_0/rr
      -- 
    rr_630_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_630_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(40), ack => ptr_deref_125_load_0_req_0); -- 
    maxPool4_cp_element_group_40: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_40"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(21) & maxPool4_CP_346_elements(42);
      gj_maxPool4_cp_element_group_40 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(40), clk => clk, reset => reset); --
    end block;
    -- CP-element group 41:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: marked-predecessors 
    -- CP-element group 41: 	43 
    -- CP-element group 41: 	118 
    -- CP-element group 41: 	122 
    -- CP-element group 41: 	126 
    -- CP-element group 41: 	130 
    -- CP-element group 41: 	134 
    -- CP-element group 41: 	138 
    -- CP-element group 41: 	142 
    -- CP-element group 41: 	146 
    -- CP-element group 41: 	150 
    -- CP-element group 41: 	154 
    -- CP-element group 41: 	158 
    -- CP-element group 41: 	162 
    -- CP-element group 41: 	166 
    -- CP-element group 41: 	170 
    -- CP-element group 41: 	174 
    -- CP-element group 41: 	178 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	43 
    -- CP-element group 41:  members (5) 
      -- CP-element group 41: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_125_update_start_
      -- CP-element group 41: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_125_Update/$entry
      -- CP-element group 41: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_125_Update/word_access_complete/$entry
      -- CP-element group 41: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_125_Update/word_access_complete/word_0/$entry
      -- CP-element group 41: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_125_Update/word_access_complete/word_0/cr
      -- 
    cr_641_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_641_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(41), ack => ptr_deref_125_load_0_req_1); -- 
    maxPool4_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 16) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_markings: IntegerArray(0 to 16)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_delays: IntegerArray(0 to 16) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 17); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(43) & maxPool4_CP_346_elements(118) & maxPool4_CP_346_elements(122) & maxPool4_CP_346_elements(126) & maxPool4_CP_346_elements(130) & maxPool4_CP_346_elements(134) & maxPool4_CP_346_elements(138) & maxPool4_CP_346_elements(142) & maxPool4_CP_346_elements(146) & maxPool4_CP_346_elements(150) & maxPool4_CP_346_elements(154) & maxPool4_CP_346_elements(158) & maxPool4_CP_346_elements(162) & maxPool4_CP_346_elements(166) & maxPool4_CP_346_elements(170) & maxPool4_CP_346_elements(174) & maxPool4_CP_346_elements(178);
      gj_maxPool4_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 17, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	40 
    -- CP-element group 42: successors 
    -- CP-element group 42: marked-successors 
    -- CP-element group 42: 	40 
    -- CP-element group 42: 	16 
    -- CP-element group 42:  members (5) 
      -- CP-element group 42: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_125_sample_completed_
      -- CP-element group 42: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_125_Sample/$exit
      -- CP-element group 42: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_125_Sample/word_access_start/$exit
      -- CP-element group 42: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_125_Sample/word_access_start/word_0/$exit
      -- CP-element group 42: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_125_Sample/word_access_start/word_0/ra
      -- 
    ra_631_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_125_load_0_ack_0, ack => maxPool4_CP_346_elements(42)); -- 
    -- CP-element group 43:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	41 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	116 
    -- CP-element group 43: 	120 
    -- CP-element group 43: 	124 
    -- CP-element group 43: 	128 
    -- CP-element group 43: 	132 
    -- CP-element group 43: 	136 
    -- CP-element group 43: 	140 
    -- CP-element group 43: 	144 
    -- CP-element group 43: 	148 
    -- CP-element group 43: 	152 
    -- CP-element group 43: 	156 
    -- CP-element group 43: 	160 
    -- CP-element group 43: 	164 
    -- CP-element group 43: 	168 
    -- CP-element group 43: 	172 
    -- CP-element group 43: 	176 
    -- CP-element group 43: marked-successors 
    -- CP-element group 43: 	41 
    -- CP-element group 43:  members (9) 
      -- CP-element group 43: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_125_update_completed_
      -- CP-element group 43: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_125_Update/$exit
      -- CP-element group 43: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_125_Update/word_access_complete/$exit
      -- CP-element group 43: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_125_Update/word_access_complete/word_0/$exit
      -- CP-element group 43: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_125_Update/word_access_complete/word_0/ca
      -- CP-element group 43: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_125_Update/ptr_deref_125_Merge/$entry
      -- CP-element group 43: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_125_Update/ptr_deref_125_Merge/$exit
      -- CP-element group 43: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_125_Update/ptr_deref_125_Merge/merge_req
      -- CP-element group 43: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_125_Update/ptr_deref_125_Merge/merge_ack
      -- 
    ca_642_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_125_load_0_ack_1, ack => maxPool4_CP_346_elements(43)); -- 
    -- CP-element group 44:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	28 
    -- CP-element group 44: marked-predecessors 
    -- CP-element group 44: 	46 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	46 
    -- CP-element group 44:  members (5) 
      -- CP-element group 44: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_129_sample_start_
      -- CP-element group 44: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_129_Sample/$entry
      -- CP-element group 44: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_129_Sample/word_access_start/$entry
      -- CP-element group 44: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_129_Sample/word_access_start/word_0/$entry
      -- CP-element group 44: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_129_Sample/word_access_start/word_0/rr
      -- 
    rr_680_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_680_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(44), ack => ptr_deref_129_load_0_req_0); -- 
    maxPool4_cp_element_group_44: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_44"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(28) & maxPool4_CP_346_elements(46);
      gj_maxPool4_cp_element_group_44 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(44), clk => clk, reset => reset); --
    end block;
    -- CP-element group 45:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: marked-predecessors 
    -- CP-element group 45: 	47 
    -- CP-element group 45: 	182 
    -- CP-element group 45: 	186 
    -- CP-element group 45: 	190 
    -- CP-element group 45: 	194 
    -- CP-element group 45: 	198 
    -- CP-element group 45: 	202 
    -- CP-element group 45: 	206 
    -- CP-element group 45: 	210 
    -- CP-element group 45: 	214 
    -- CP-element group 45: 	218 
    -- CP-element group 45: 	222 
    -- CP-element group 45: 	226 
    -- CP-element group 45: 	230 
    -- CP-element group 45: 	234 
    -- CP-element group 45: 	238 
    -- CP-element group 45: 	242 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	47 
    -- CP-element group 45:  members (5) 
      -- CP-element group 45: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_129_update_start_
      -- CP-element group 45: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_129_Update/$entry
      -- CP-element group 45: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_129_Update/word_access_complete/$entry
      -- CP-element group 45: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_129_Update/word_access_complete/word_0/$entry
      -- CP-element group 45: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_129_Update/word_access_complete/word_0/cr
      -- 
    cr_691_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_691_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(45), ack => ptr_deref_129_load_0_req_1); -- 
    maxPool4_cp_element_group_45: block -- 
      constant place_capacities: IntegerArray(0 to 16) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_markings: IntegerArray(0 to 16)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_delays: IntegerArray(0 to 16) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_45"; 
      signal preds: BooleanArray(1 to 17); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(47) & maxPool4_CP_346_elements(182) & maxPool4_CP_346_elements(186) & maxPool4_CP_346_elements(190) & maxPool4_CP_346_elements(194) & maxPool4_CP_346_elements(198) & maxPool4_CP_346_elements(202) & maxPool4_CP_346_elements(206) & maxPool4_CP_346_elements(210) & maxPool4_CP_346_elements(214) & maxPool4_CP_346_elements(218) & maxPool4_CP_346_elements(222) & maxPool4_CP_346_elements(226) & maxPool4_CP_346_elements(230) & maxPool4_CP_346_elements(234) & maxPool4_CP_346_elements(238) & maxPool4_CP_346_elements(242);
      gj_maxPool4_cp_element_group_45 : generic_join generic map(name => joinName, number_of_predecessors => 17, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(45), clk => clk, reset => reset); --
    end block;
    -- CP-element group 46:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	44 
    -- CP-element group 46: successors 
    -- CP-element group 46: marked-successors 
    -- CP-element group 46: 	44 
    -- CP-element group 46: 	23 
    -- CP-element group 46:  members (5) 
      -- CP-element group 46: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_129_sample_completed_
      -- CP-element group 46: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_129_Sample/$exit
      -- CP-element group 46: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_129_Sample/word_access_start/$exit
      -- CP-element group 46: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_129_Sample/word_access_start/word_0/$exit
      -- CP-element group 46: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_129_Sample/word_access_start/word_0/ra
      -- 
    ra_681_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_129_load_0_ack_0, ack => maxPool4_CP_346_elements(46)); -- 
    -- CP-element group 47:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	45 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	180 
    -- CP-element group 47: 	184 
    -- CP-element group 47: 	188 
    -- CP-element group 47: 	192 
    -- CP-element group 47: 	196 
    -- CP-element group 47: 	200 
    -- CP-element group 47: 	204 
    -- CP-element group 47: 	208 
    -- CP-element group 47: 	212 
    -- CP-element group 47: 	216 
    -- CP-element group 47: 	220 
    -- CP-element group 47: 	224 
    -- CP-element group 47: 	228 
    -- CP-element group 47: 	232 
    -- CP-element group 47: 	236 
    -- CP-element group 47: 	240 
    -- CP-element group 47: marked-successors 
    -- CP-element group 47: 	45 
    -- CP-element group 47:  members (9) 
      -- CP-element group 47: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_129_update_completed_
      -- CP-element group 47: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_129_Update/$exit
      -- CP-element group 47: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_129_Update/word_access_complete/$exit
      -- CP-element group 47: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_129_Update/word_access_complete/word_0/$exit
      -- CP-element group 47: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_129_Update/word_access_complete/word_0/ca
      -- CP-element group 47: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_129_Update/ptr_deref_129_Merge/$entry
      -- CP-element group 47: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_129_Update/ptr_deref_129_Merge/$exit
      -- CP-element group 47: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_129_Update/ptr_deref_129_Merge/merge_req
      -- CP-element group 47: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_129_Update/ptr_deref_129_Merge/merge_ack
      -- 
    ca_692_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_129_load_0_ack_1, ack => maxPool4_CP_346_elements(47)); -- 
    -- CP-element group 48:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	35 
    -- CP-element group 48: marked-predecessors 
    -- CP-element group 48: 	50 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	50 
    -- CP-element group 48:  members (5) 
      -- CP-element group 48: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_133_sample_start_
      -- CP-element group 48: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_133_Sample/$entry
      -- CP-element group 48: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_133_Sample/word_access_start/$entry
      -- CP-element group 48: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_133_Sample/word_access_start/word_0/$entry
      -- CP-element group 48: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_133_Sample/word_access_start/word_0/rr
      -- 
    rr_730_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_730_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(48), ack => ptr_deref_133_load_0_req_0); -- 
    maxPool4_cp_element_group_48: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_48"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(35) & maxPool4_CP_346_elements(50);
      gj_maxPool4_cp_element_group_48 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(48), clk => clk, reset => reset); --
    end block;
    -- CP-element group 49:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: marked-predecessors 
    -- CP-element group 49: 	51 
    -- CP-element group 49: 	246 
    -- CP-element group 49: 	250 
    -- CP-element group 49: 	254 
    -- CP-element group 49: 	258 
    -- CP-element group 49: 	262 
    -- CP-element group 49: 	266 
    -- CP-element group 49: 	270 
    -- CP-element group 49: 	274 
    -- CP-element group 49: 	278 
    -- CP-element group 49: 	282 
    -- CP-element group 49: 	286 
    -- CP-element group 49: 	290 
    -- CP-element group 49: 	294 
    -- CP-element group 49: 	298 
    -- CP-element group 49: 	302 
    -- CP-element group 49: 	306 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (5) 
      -- CP-element group 49: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_133_update_start_
      -- CP-element group 49: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_133_Update/$entry
      -- CP-element group 49: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_133_Update/word_access_complete/$entry
      -- CP-element group 49: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_133_Update/word_access_complete/word_0/$entry
      -- CP-element group 49: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_133_Update/word_access_complete/word_0/cr
      -- 
    cr_741_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_741_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(49), ack => ptr_deref_133_load_0_req_1); -- 
    maxPool4_cp_element_group_49: block -- 
      constant place_capacities: IntegerArray(0 to 16) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_markings: IntegerArray(0 to 16)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_delays: IntegerArray(0 to 16) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_49"; 
      signal preds: BooleanArray(1 to 17); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(51) & maxPool4_CP_346_elements(246) & maxPool4_CP_346_elements(250) & maxPool4_CP_346_elements(254) & maxPool4_CP_346_elements(258) & maxPool4_CP_346_elements(262) & maxPool4_CP_346_elements(266) & maxPool4_CP_346_elements(270) & maxPool4_CP_346_elements(274) & maxPool4_CP_346_elements(278) & maxPool4_CP_346_elements(282) & maxPool4_CP_346_elements(286) & maxPool4_CP_346_elements(290) & maxPool4_CP_346_elements(294) & maxPool4_CP_346_elements(298) & maxPool4_CP_346_elements(302) & maxPool4_CP_346_elements(306);
      gj_maxPool4_cp_element_group_49 : generic_join generic map(name => joinName, number_of_predecessors => 17, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(49), clk => clk, reset => reset); --
    end block;
    -- CP-element group 50:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	48 
    -- CP-element group 50: successors 
    -- CP-element group 50: marked-successors 
    -- CP-element group 50: 	48 
    -- CP-element group 50: 	30 
    -- CP-element group 50:  members (5) 
      -- CP-element group 50: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_133_sample_completed_
      -- CP-element group 50: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_133_Sample/$exit
      -- CP-element group 50: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_133_Sample/word_access_start/$exit
      -- CP-element group 50: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_133_Sample/word_access_start/word_0/$exit
      -- CP-element group 50: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_133_Sample/word_access_start/word_0/ra
      -- 
    ra_731_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_133_load_0_ack_0, ack => maxPool4_CP_346_elements(50)); -- 
    -- CP-element group 51:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	244 
    -- CP-element group 51: 	248 
    -- CP-element group 51: 	252 
    -- CP-element group 51: 	256 
    -- CP-element group 51: 	260 
    -- CP-element group 51: 	264 
    -- CP-element group 51: 	268 
    -- CP-element group 51: 	272 
    -- CP-element group 51: 	276 
    -- CP-element group 51: 	280 
    -- CP-element group 51: 	284 
    -- CP-element group 51: 	288 
    -- CP-element group 51: 	292 
    -- CP-element group 51: 	296 
    -- CP-element group 51: 	300 
    -- CP-element group 51: 	304 
    -- CP-element group 51: marked-successors 
    -- CP-element group 51: 	49 
    -- CP-element group 51:  members (9) 
      -- CP-element group 51: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_133_update_completed_
      -- CP-element group 51: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_133_Update/$exit
      -- CP-element group 51: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_133_Update/word_access_complete/$exit
      -- CP-element group 51: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_133_Update/word_access_complete/word_0/$exit
      -- CP-element group 51: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_133_Update/word_access_complete/word_0/ca
      -- CP-element group 51: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_133_Update/ptr_deref_133_Merge/$entry
      -- CP-element group 51: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_133_Update/ptr_deref_133_Merge/$exit
      -- CP-element group 51: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_133_Update/ptr_deref_133_Merge/merge_req
      -- CP-element group 51: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_133_Update/ptr_deref_133_Merge/merge_ack
      -- 
    ca_742_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_133_load_0_ack_1, ack => maxPool4_CP_346_elements(51)); -- 
    -- CP-element group 52:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	39 
    -- CP-element group 52: marked-predecessors 
    -- CP-element group 52: 	54 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 assign_stmt_97_to_assign_stmt_1138/slice_138_sample_start_
      -- CP-element group 52: 	 assign_stmt_97_to_assign_stmt_1138/slice_138_Sample/$entry
      -- CP-element group 52: 	 assign_stmt_97_to_assign_stmt_1138/slice_138_Sample/rr
      -- 
    rr_755_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_755_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(52), ack => slice_138_inst_req_0); -- 
    maxPool4_cp_element_group_52: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_52"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(39) & maxPool4_CP_346_elements(54);
      gj_maxPool4_cp_element_group_52 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(52), clk => clk, reset => reset); --
    end block;
    -- CP-element group 53:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: marked-predecessors 
    -- CP-element group 53: 	55 
    -- CP-element group 53: 	321 
    -- CP-element group 53: 	386 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 assign_stmt_97_to_assign_stmt_1138/slice_138_update_start_
      -- CP-element group 53: 	 assign_stmt_97_to_assign_stmt_1138/slice_138_Update/$entry
      -- CP-element group 53: 	 assign_stmt_97_to_assign_stmt_1138/slice_138_Update/cr
      -- 
    cr_760_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_760_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(53), ack => slice_138_inst_req_1); -- 
    maxPool4_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(55) & maxPool4_CP_346_elements(321) & maxPool4_CP_346_elements(386);
      gj_maxPool4_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54: marked-successors 
    -- CP-element group 54: 	37 
    -- CP-element group 54: 	52 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 assign_stmt_97_to_assign_stmt_1138/slice_138_sample_completed_
      -- CP-element group 54: 	 assign_stmt_97_to_assign_stmt_1138/slice_138_Sample/$exit
      -- CP-element group 54: 	 assign_stmt_97_to_assign_stmt_1138/slice_138_Sample/ra
      -- 
    ra_756_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_138_inst_ack_0, ack => maxPool4_CP_346_elements(54)); -- 
    -- CP-element group 55:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	319 
    -- CP-element group 55: 	384 
    -- CP-element group 55: marked-successors 
    -- CP-element group 55: 	53 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 assign_stmt_97_to_assign_stmt_1138/slice_138_update_completed_
      -- CP-element group 55: 	 assign_stmt_97_to_assign_stmt_1138/slice_138_Update/$exit
      -- CP-element group 55: 	 assign_stmt_97_to_assign_stmt_1138/slice_138_Update/ca
      -- 
    ca_761_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_138_inst_ack_1, ack => maxPool4_CP_346_elements(55)); -- 
    -- CP-element group 56:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	39 
    -- CP-element group 56: marked-predecessors 
    -- CP-element group 56: 	58 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	58 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 assign_stmt_97_to_assign_stmt_1138/slice_142_sample_start_
      -- CP-element group 56: 	 assign_stmt_97_to_assign_stmt_1138/slice_142_Sample/$entry
      -- CP-element group 56: 	 assign_stmt_97_to_assign_stmt_1138/slice_142_Sample/rr
      -- 
    rr_769_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_769_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(56), ack => slice_142_inst_req_0); -- 
    maxPool4_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(39) & maxPool4_CP_346_elements(58);
      gj_maxPool4_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: marked-predecessors 
    -- CP-element group 57: 	59 
    -- CP-element group 57: 	321 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	59 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 assign_stmt_97_to_assign_stmt_1138/slice_142_update_start_
      -- CP-element group 57: 	 assign_stmt_97_to_assign_stmt_1138/slice_142_Update/$entry
      -- CP-element group 57: 	 assign_stmt_97_to_assign_stmt_1138/slice_142_Update/cr
      -- 
    cr_774_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_774_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(57), ack => slice_142_inst_req_1); -- 
    maxPool4_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(59) & maxPool4_CP_346_elements(321);
      gj_maxPool4_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	56 
    -- CP-element group 58: successors 
    -- CP-element group 58: marked-successors 
    -- CP-element group 58: 	37 
    -- CP-element group 58: 	56 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 assign_stmt_97_to_assign_stmt_1138/slice_142_sample_completed_
      -- CP-element group 58: 	 assign_stmt_97_to_assign_stmt_1138/slice_142_Sample/$exit
      -- CP-element group 58: 	 assign_stmt_97_to_assign_stmt_1138/slice_142_Sample/ra
      -- 
    ra_770_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_142_inst_ack_0, ack => maxPool4_CP_346_elements(58)); -- 
    -- CP-element group 59:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	57 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	319 
    -- CP-element group 59: marked-successors 
    -- CP-element group 59: 	57 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 assign_stmt_97_to_assign_stmt_1138/slice_142_update_completed_
      -- CP-element group 59: 	 assign_stmt_97_to_assign_stmt_1138/slice_142_Update/$exit
      -- CP-element group 59: 	 assign_stmt_97_to_assign_stmt_1138/slice_142_Update/ca
      -- 
    ca_775_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_142_inst_ack_1, ack => maxPool4_CP_346_elements(59)); -- 
    -- CP-element group 60:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	39 
    -- CP-element group 60: marked-predecessors 
    -- CP-element group 60: 	62 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	62 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 assign_stmt_97_to_assign_stmt_1138/slice_146_sample_start_
      -- CP-element group 60: 	 assign_stmt_97_to_assign_stmt_1138/slice_146_Sample/$entry
      -- CP-element group 60: 	 assign_stmt_97_to_assign_stmt_1138/slice_146_Sample/rr
      -- 
    rr_783_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_783_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(60), ack => slice_146_inst_req_0); -- 
    maxPool4_cp_element_group_60: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_60"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(39) & maxPool4_CP_346_elements(62);
      gj_maxPool4_cp_element_group_60 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(60), clk => clk, reset => reset); --
    end block;
    -- CP-element group 61:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: marked-predecessors 
    -- CP-element group 61: 	63 
    -- CP-element group 61: 	321 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	63 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 assign_stmt_97_to_assign_stmt_1138/slice_146_update_start_
      -- CP-element group 61: 	 assign_stmt_97_to_assign_stmt_1138/slice_146_Update/$entry
      -- CP-element group 61: 	 assign_stmt_97_to_assign_stmt_1138/slice_146_Update/cr
      -- 
    cr_788_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_788_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(61), ack => slice_146_inst_req_1); -- 
    maxPool4_cp_element_group_61: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_61"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(63) & maxPool4_CP_346_elements(321);
      gj_maxPool4_cp_element_group_61 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(61), clk => clk, reset => reset); --
    end block;
    -- CP-element group 62:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	60 
    -- CP-element group 62: successors 
    -- CP-element group 62: marked-successors 
    -- CP-element group 62: 	37 
    -- CP-element group 62: 	60 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 assign_stmt_97_to_assign_stmt_1138/slice_146_sample_completed_
      -- CP-element group 62: 	 assign_stmt_97_to_assign_stmt_1138/slice_146_Sample/$exit
      -- CP-element group 62: 	 assign_stmt_97_to_assign_stmt_1138/slice_146_Sample/ra
      -- 
    ra_784_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_146_inst_ack_0, ack => maxPool4_CP_346_elements(62)); -- 
    -- CP-element group 63:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	61 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	319 
    -- CP-element group 63: marked-successors 
    -- CP-element group 63: 	61 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 assign_stmt_97_to_assign_stmt_1138/slice_146_update_completed_
      -- CP-element group 63: 	 assign_stmt_97_to_assign_stmt_1138/slice_146_Update/$exit
      -- CP-element group 63: 	 assign_stmt_97_to_assign_stmt_1138/slice_146_Update/ca
      -- 
    ca_789_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_146_inst_ack_1, ack => maxPool4_CP_346_elements(63)); -- 
    -- CP-element group 64:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	39 
    -- CP-element group 64: marked-predecessors 
    -- CP-element group 64: 	66 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	66 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 assign_stmt_97_to_assign_stmt_1138/slice_150_sample_start_
      -- CP-element group 64: 	 assign_stmt_97_to_assign_stmt_1138/slice_150_Sample/$entry
      -- CP-element group 64: 	 assign_stmt_97_to_assign_stmt_1138/slice_150_Sample/rr
      -- 
    rr_797_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_797_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(64), ack => slice_150_inst_req_0); -- 
    maxPool4_cp_element_group_64: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_64"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(39) & maxPool4_CP_346_elements(66);
      gj_maxPool4_cp_element_group_64 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(64), clk => clk, reset => reset); --
    end block;
    -- CP-element group 65:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: marked-predecessors 
    -- CP-element group 65: 	67 
    -- CP-element group 65: 	321 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	67 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 assign_stmt_97_to_assign_stmt_1138/slice_150_update_start_
      -- CP-element group 65: 	 assign_stmt_97_to_assign_stmt_1138/slice_150_Update/$entry
      -- CP-element group 65: 	 assign_stmt_97_to_assign_stmt_1138/slice_150_Update/cr
      -- 
    cr_802_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_802_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(65), ack => slice_150_inst_req_1); -- 
    maxPool4_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(67) & maxPool4_CP_346_elements(321);
      gj_maxPool4_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	64 
    -- CP-element group 66: successors 
    -- CP-element group 66: marked-successors 
    -- CP-element group 66: 	37 
    -- CP-element group 66: 	64 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 assign_stmt_97_to_assign_stmt_1138/slice_150_sample_completed_
      -- CP-element group 66: 	 assign_stmt_97_to_assign_stmt_1138/slice_150_Sample/$exit
      -- CP-element group 66: 	 assign_stmt_97_to_assign_stmt_1138/slice_150_Sample/ra
      -- 
    ra_798_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_150_inst_ack_0, ack => maxPool4_CP_346_elements(66)); -- 
    -- CP-element group 67:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	65 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	319 
    -- CP-element group 67: marked-successors 
    -- CP-element group 67: 	65 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 assign_stmt_97_to_assign_stmt_1138/slice_150_update_completed_
      -- CP-element group 67: 	 assign_stmt_97_to_assign_stmt_1138/slice_150_Update/$exit
      -- CP-element group 67: 	 assign_stmt_97_to_assign_stmt_1138/slice_150_Update/ca
      -- 
    ca_803_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_150_inst_ack_1, ack => maxPool4_CP_346_elements(67)); -- 
    -- CP-element group 68:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	39 
    -- CP-element group 68: marked-predecessors 
    -- CP-element group 68: 	70 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 assign_stmt_97_to_assign_stmt_1138/slice_154_sample_start_
      -- CP-element group 68: 	 assign_stmt_97_to_assign_stmt_1138/slice_154_Sample/$entry
      -- CP-element group 68: 	 assign_stmt_97_to_assign_stmt_1138/slice_154_Sample/rr
      -- 
    rr_811_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_811_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(68), ack => slice_154_inst_req_0); -- 
    maxPool4_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(39) & maxPool4_CP_346_elements(70);
      gj_maxPool4_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: marked-predecessors 
    -- CP-element group 69: 	71 
    -- CP-element group 69: 	340 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	71 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 assign_stmt_97_to_assign_stmt_1138/slice_154_update_start_
      -- CP-element group 69: 	 assign_stmt_97_to_assign_stmt_1138/slice_154_Update/$entry
      -- CP-element group 69: 	 assign_stmt_97_to_assign_stmt_1138/slice_154_Update/cr
      -- 
    cr_816_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_816_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(69), ack => slice_154_inst_req_1); -- 
    maxPool4_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(71) & maxPool4_CP_346_elements(340);
      gj_maxPool4_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: marked-successors 
    -- CP-element group 70: 	37 
    -- CP-element group 70: 	68 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 assign_stmt_97_to_assign_stmt_1138/slice_154_sample_completed_
      -- CP-element group 70: 	 assign_stmt_97_to_assign_stmt_1138/slice_154_Sample/$exit
      -- CP-element group 70: 	 assign_stmt_97_to_assign_stmt_1138/slice_154_Sample/ra
      -- 
    ra_812_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_154_inst_ack_0, ack => maxPool4_CP_346_elements(70)); -- 
    -- CP-element group 71:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	69 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	338 
    -- CP-element group 71: marked-successors 
    -- CP-element group 71: 	69 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 assign_stmt_97_to_assign_stmt_1138/slice_154_update_completed_
      -- CP-element group 71: 	 assign_stmt_97_to_assign_stmt_1138/slice_154_Update/$exit
      -- CP-element group 71: 	 assign_stmt_97_to_assign_stmt_1138/slice_154_Update/ca
      -- 
    ca_817_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_154_inst_ack_1, ack => maxPool4_CP_346_elements(71)); -- 
    -- CP-element group 72:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	39 
    -- CP-element group 72: marked-predecessors 
    -- CP-element group 72: 	74 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	74 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 assign_stmt_97_to_assign_stmt_1138/slice_158_sample_start_
      -- CP-element group 72: 	 assign_stmt_97_to_assign_stmt_1138/slice_158_Sample/$entry
      -- CP-element group 72: 	 assign_stmt_97_to_assign_stmt_1138/slice_158_Sample/rr
      -- 
    rr_825_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_825_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(72), ack => slice_158_inst_req_0); -- 
    maxPool4_cp_element_group_72: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_72"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(39) & maxPool4_CP_346_elements(74);
      gj_maxPool4_cp_element_group_72 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(72), clk => clk, reset => reset); --
    end block;
    -- CP-element group 73:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: marked-predecessors 
    -- CP-element group 73: 	75 
    -- CP-element group 73: 	340 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	75 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 assign_stmt_97_to_assign_stmt_1138/slice_158_update_start_
      -- CP-element group 73: 	 assign_stmt_97_to_assign_stmt_1138/slice_158_Update/$entry
      -- CP-element group 73: 	 assign_stmt_97_to_assign_stmt_1138/slice_158_Update/cr
      -- 
    cr_830_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_830_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(73), ack => slice_158_inst_req_1); -- 
    maxPool4_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(75) & maxPool4_CP_346_elements(340);
      gj_maxPool4_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	72 
    -- CP-element group 74: successors 
    -- CP-element group 74: marked-successors 
    -- CP-element group 74: 	37 
    -- CP-element group 74: 	72 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 assign_stmt_97_to_assign_stmt_1138/slice_158_sample_completed_
      -- CP-element group 74: 	 assign_stmt_97_to_assign_stmt_1138/slice_158_Sample/$exit
      -- CP-element group 74: 	 assign_stmt_97_to_assign_stmt_1138/slice_158_Sample/ra
      -- 
    ra_826_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_158_inst_ack_0, ack => maxPool4_CP_346_elements(74)); -- 
    -- CP-element group 75:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	73 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	338 
    -- CP-element group 75: marked-successors 
    -- CP-element group 75: 	73 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 assign_stmt_97_to_assign_stmt_1138/slice_158_update_completed_
      -- CP-element group 75: 	 assign_stmt_97_to_assign_stmt_1138/slice_158_Update/$exit
      -- CP-element group 75: 	 assign_stmt_97_to_assign_stmt_1138/slice_158_Update/ca
      -- 
    ca_831_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_158_inst_ack_1, ack => maxPool4_CP_346_elements(75)); -- 
    -- CP-element group 76:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	39 
    -- CP-element group 76: marked-predecessors 
    -- CP-element group 76: 	78 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	78 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 assign_stmt_97_to_assign_stmt_1138/slice_162_sample_start_
      -- CP-element group 76: 	 assign_stmt_97_to_assign_stmt_1138/slice_162_Sample/$entry
      -- CP-element group 76: 	 assign_stmt_97_to_assign_stmt_1138/slice_162_Sample/rr
      -- 
    rr_839_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_839_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(76), ack => slice_162_inst_req_0); -- 
    maxPool4_cp_element_group_76: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_76"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(39) & maxPool4_CP_346_elements(78);
      gj_maxPool4_cp_element_group_76 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(76), clk => clk, reset => reset); --
    end block;
    -- CP-element group 77:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: marked-predecessors 
    -- CP-element group 77: 	79 
    -- CP-element group 77: 	340 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	79 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 assign_stmt_97_to_assign_stmt_1138/slice_162_update_start_
      -- CP-element group 77: 	 assign_stmt_97_to_assign_stmt_1138/slice_162_Update/$entry
      -- CP-element group 77: 	 assign_stmt_97_to_assign_stmt_1138/slice_162_Update/cr
      -- 
    cr_844_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_844_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(77), ack => slice_162_inst_req_1); -- 
    maxPool4_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(79) & maxPool4_CP_346_elements(340);
      gj_maxPool4_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	76 
    -- CP-element group 78: successors 
    -- CP-element group 78: marked-successors 
    -- CP-element group 78: 	37 
    -- CP-element group 78: 	76 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 assign_stmt_97_to_assign_stmt_1138/slice_162_sample_completed_
      -- CP-element group 78: 	 assign_stmt_97_to_assign_stmt_1138/slice_162_Sample/$exit
      -- CP-element group 78: 	 assign_stmt_97_to_assign_stmt_1138/slice_162_Sample/ra
      -- 
    ra_840_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_162_inst_ack_0, ack => maxPool4_CP_346_elements(78)); -- 
    -- CP-element group 79:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	77 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	338 
    -- CP-element group 79: marked-successors 
    -- CP-element group 79: 	77 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 assign_stmt_97_to_assign_stmt_1138/slice_162_update_completed_
      -- CP-element group 79: 	 assign_stmt_97_to_assign_stmt_1138/slice_162_Update/$exit
      -- CP-element group 79: 	 assign_stmt_97_to_assign_stmt_1138/slice_162_Update/ca
      -- 
    ca_845_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_162_inst_ack_1, ack => maxPool4_CP_346_elements(79)); -- 
    -- CP-element group 80:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	39 
    -- CP-element group 80: marked-predecessors 
    -- CP-element group 80: 	82 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	82 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 assign_stmt_97_to_assign_stmt_1138/slice_166_sample_start_
      -- CP-element group 80: 	 assign_stmt_97_to_assign_stmt_1138/slice_166_Sample/$entry
      -- CP-element group 80: 	 assign_stmt_97_to_assign_stmt_1138/slice_166_Sample/rr
      -- 
    rr_853_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_853_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(80), ack => slice_166_inst_req_0); -- 
    maxPool4_cp_element_group_80: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_80"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(39) & maxPool4_CP_346_elements(82);
      gj_maxPool4_cp_element_group_80 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(80), clk => clk, reset => reset); --
    end block;
    -- CP-element group 81:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: marked-predecessors 
    -- CP-element group 81: 	83 
    -- CP-element group 81: 	340 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	83 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 assign_stmt_97_to_assign_stmt_1138/slice_166_update_start_
      -- CP-element group 81: 	 assign_stmt_97_to_assign_stmt_1138/slice_166_Update/$entry
      -- CP-element group 81: 	 assign_stmt_97_to_assign_stmt_1138/slice_166_Update/cr
      -- 
    cr_858_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_858_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(81), ack => slice_166_inst_req_1); -- 
    maxPool4_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(83) & maxPool4_CP_346_elements(340);
      gj_maxPool4_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	80 
    -- CP-element group 82: successors 
    -- CP-element group 82: marked-successors 
    -- CP-element group 82: 	37 
    -- CP-element group 82: 	80 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 assign_stmt_97_to_assign_stmt_1138/slice_166_sample_completed_
      -- CP-element group 82: 	 assign_stmt_97_to_assign_stmt_1138/slice_166_Sample/$exit
      -- CP-element group 82: 	 assign_stmt_97_to_assign_stmt_1138/slice_166_Sample/ra
      -- 
    ra_854_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_166_inst_ack_0, ack => maxPool4_CP_346_elements(82)); -- 
    -- CP-element group 83:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	81 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	338 
    -- CP-element group 83: marked-successors 
    -- CP-element group 83: 	81 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 assign_stmt_97_to_assign_stmt_1138/slice_166_update_completed_
      -- CP-element group 83: 	 assign_stmt_97_to_assign_stmt_1138/slice_166_Update/$exit
      -- CP-element group 83: 	 assign_stmt_97_to_assign_stmt_1138/slice_166_Update/ca
      -- 
    ca_859_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_166_inst_ack_1, ack => maxPool4_CP_346_elements(83)); -- 
    -- CP-element group 84:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	39 
    -- CP-element group 84: marked-predecessors 
    -- CP-element group 84: 	86 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 assign_stmt_97_to_assign_stmt_1138/slice_170_sample_start_
      -- CP-element group 84: 	 assign_stmt_97_to_assign_stmt_1138/slice_170_Sample/$entry
      -- CP-element group 84: 	 assign_stmt_97_to_assign_stmt_1138/slice_170_Sample/rr
      -- 
    rr_867_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_867_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(84), ack => slice_170_inst_req_0); -- 
    maxPool4_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(39) & maxPool4_CP_346_elements(86);
      gj_maxPool4_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: marked-predecessors 
    -- CP-element group 85: 	87 
    -- CP-element group 85: 	359 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 assign_stmt_97_to_assign_stmt_1138/slice_170_update_start_
      -- CP-element group 85: 	 assign_stmt_97_to_assign_stmt_1138/slice_170_Update/$entry
      -- CP-element group 85: 	 assign_stmt_97_to_assign_stmt_1138/slice_170_Update/cr
      -- 
    cr_872_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_872_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(85), ack => slice_170_inst_req_1); -- 
    maxPool4_cp_element_group_85: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_85"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(87) & maxPool4_CP_346_elements(359);
      gj_maxPool4_cp_element_group_85 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(85), clk => clk, reset => reset); --
    end block;
    -- CP-element group 86:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: successors 
    -- CP-element group 86: marked-successors 
    -- CP-element group 86: 	37 
    -- CP-element group 86: 	84 
    -- CP-element group 86:  members (3) 
      -- CP-element group 86: 	 assign_stmt_97_to_assign_stmt_1138/slice_170_sample_completed_
      -- CP-element group 86: 	 assign_stmt_97_to_assign_stmt_1138/slice_170_Sample/$exit
      -- CP-element group 86: 	 assign_stmt_97_to_assign_stmt_1138/slice_170_Sample/ra
      -- 
    ra_868_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_170_inst_ack_0, ack => maxPool4_CP_346_elements(86)); -- 
    -- CP-element group 87:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	357 
    -- CP-element group 87: marked-successors 
    -- CP-element group 87: 	85 
    -- CP-element group 87:  members (3) 
      -- CP-element group 87: 	 assign_stmt_97_to_assign_stmt_1138/slice_170_update_completed_
      -- CP-element group 87: 	 assign_stmt_97_to_assign_stmt_1138/slice_170_Update/$exit
      -- CP-element group 87: 	 assign_stmt_97_to_assign_stmt_1138/slice_170_Update/ca
      -- 
    ca_873_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_170_inst_ack_1, ack => maxPool4_CP_346_elements(87)); -- 
    -- CP-element group 88:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	39 
    -- CP-element group 88: marked-predecessors 
    -- CP-element group 88: 	90 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	90 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 assign_stmt_97_to_assign_stmt_1138/slice_174_sample_start_
      -- CP-element group 88: 	 assign_stmt_97_to_assign_stmt_1138/slice_174_Sample/$entry
      -- CP-element group 88: 	 assign_stmt_97_to_assign_stmt_1138/slice_174_Sample/rr
      -- 
    rr_881_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_881_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(88), ack => slice_174_inst_req_0); -- 
    maxPool4_cp_element_group_88: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_88"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(39) & maxPool4_CP_346_elements(90);
      gj_maxPool4_cp_element_group_88 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(88), clk => clk, reset => reset); --
    end block;
    -- CP-element group 89:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: marked-predecessors 
    -- CP-element group 89: 	91 
    -- CP-element group 89: 	359 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 assign_stmt_97_to_assign_stmt_1138/slice_174_update_start_
      -- CP-element group 89: 	 assign_stmt_97_to_assign_stmt_1138/slice_174_Update/$entry
      -- CP-element group 89: 	 assign_stmt_97_to_assign_stmt_1138/slice_174_Update/cr
      -- 
    cr_886_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_886_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(89), ack => slice_174_inst_req_1); -- 
    maxPool4_cp_element_group_89: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_89"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(91) & maxPool4_CP_346_elements(359);
      gj_maxPool4_cp_element_group_89 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(89), clk => clk, reset => reset); --
    end block;
    -- CP-element group 90:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	88 
    -- CP-element group 90: successors 
    -- CP-element group 90: marked-successors 
    -- CP-element group 90: 	37 
    -- CP-element group 90: 	88 
    -- CP-element group 90:  members (3) 
      -- CP-element group 90: 	 assign_stmt_97_to_assign_stmt_1138/slice_174_sample_completed_
      -- CP-element group 90: 	 assign_stmt_97_to_assign_stmt_1138/slice_174_Sample/$exit
      -- CP-element group 90: 	 assign_stmt_97_to_assign_stmt_1138/slice_174_Sample/ra
      -- 
    ra_882_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_174_inst_ack_0, ack => maxPool4_CP_346_elements(90)); -- 
    -- CP-element group 91:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	357 
    -- CP-element group 91: marked-successors 
    -- CP-element group 91: 	89 
    -- CP-element group 91:  members (3) 
      -- CP-element group 91: 	 assign_stmt_97_to_assign_stmt_1138/slice_174_update_completed_
      -- CP-element group 91: 	 assign_stmt_97_to_assign_stmt_1138/slice_174_Update/$exit
      -- CP-element group 91: 	 assign_stmt_97_to_assign_stmt_1138/slice_174_Update/ca
      -- 
    ca_887_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_174_inst_ack_1, ack => maxPool4_CP_346_elements(91)); -- 
    -- CP-element group 92:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	39 
    -- CP-element group 92: marked-predecessors 
    -- CP-element group 92: 	94 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	94 
    -- CP-element group 92:  members (3) 
      -- CP-element group 92: 	 assign_stmt_97_to_assign_stmt_1138/slice_178_sample_start_
      -- CP-element group 92: 	 assign_stmt_97_to_assign_stmt_1138/slice_178_Sample/$entry
      -- CP-element group 92: 	 assign_stmt_97_to_assign_stmt_1138/slice_178_Sample/rr
      -- 
    rr_895_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_895_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(92), ack => slice_178_inst_req_0); -- 
    maxPool4_cp_element_group_92: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_92"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(39) & maxPool4_CP_346_elements(94);
      gj_maxPool4_cp_element_group_92 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(92), clk => clk, reset => reset); --
    end block;
    -- CP-element group 93:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: marked-predecessors 
    -- CP-element group 93: 	95 
    -- CP-element group 93: 	359 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 assign_stmt_97_to_assign_stmt_1138/slice_178_update_start_
      -- CP-element group 93: 	 assign_stmt_97_to_assign_stmt_1138/slice_178_Update/$entry
      -- CP-element group 93: 	 assign_stmt_97_to_assign_stmt_1138/slice_178_Update/cr
      -- 
    cr_900_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_900_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(93), ack => slice_178_inst_req_1); -- 
    maxPool4_cp_element_group_93: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_93"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(95) & maxPool4_CP_346_elements(359);
      gj_maxPool4_cp_element_group_93 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(93), clk => clk, reset => reset); --
    end block;
    -- CP-element group 94:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	92 
    -- CP-element group 94: successors 
    -- CP-element group 94: marked-successors 
    -- CP-element group 94: 	37 
    -- CP-element group 94: 	92 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 assign_stmt_97_to_assign_stmt_1138/slice_178_sample_completed_
      -- CP-element group 94: 	 assign_stmt_97_to_assign_stmt_1138/slice_178_Sample/$exit
      -- CP-element group 94: 	 assign_stmt_97_to_assign_stmt_1138/slice_178_Sample/ra
      -- 
    ra_896_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_178_inst_ack_0, ack => maxPool4_CP_346_elements(94)); -- 
    -- CP-element group 95:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	357 
    -- CP-element group 95: marked-successors 
    -- CP-element group 95: 	93 
    -- CP-element group 95:  members (3) 
      -- CP-element group 95: 	 assign_stmt_97_to_assign_stmt_1138/slice_178_update_completed_
      -- CP-element group 95: 	 assign_stmt_97_to_assign_stmt_1138/slice_178_Update/$exit
      -- CP-element group 95: 	 assign_stmt_97_to_assign_stmt_1138/slice_178_Update/ca
      -- 
    ca_901_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_178_inst_ack_1, ack => maxPool4_CP_346_elements(95)); -- 
    -- CP-element group 96:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	39 
    -- CP-element group 96: marked-predecessors 
    -- CP-element group 96: 	98 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	98 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 assign_stmt_97_to_assign_stmt_1138/slice_182_sample_start_
      -- CP-element group 96: 	 assign_stmt_97_to_assign_stmt_1138/slice_182_Sample/$entry
      -- CP-element group 96: 	 assign_stmt_97_to_assign_stmt_1138/slice_182_Sample/rr
      -- 
    rr_909_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_909_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(96), ack => slice_182_inst_req_0); -- 
    maxPool4_cp_element_group_96: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_96"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(39) & maxPool4_CP_346_elements(98);
      gj_maxPool4_cp_element_group_96 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(96), clk => clk, reset => reset); --
    end block;
    -- CP-element group 97:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: marked-predecessors 
    -- CP-element group 97: 	99 
    -- CP-element group 97: 	359 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	99 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 assign_stmt_97_to_assign_stmt_1138/slice_182_update_start_
      -- CP-element group 97: 	 assign_stmt_97_to_assign_stmt_1138/slice_182_Update/$entry
      -- CP-element group 97: 	 assign_stmt_97_to_assign_stmt_1138/slice_182_Update/cr
      -- 
    cr_914_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_914_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(97), ack => slice_182_inst_req_1); -- 
    maxPool4_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "maxPool4_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(99) & maxPool4_CP_346_elements(359);
      gj_maxPool4_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	96 
    -- CP-element group 98: successors 
    -- CP-element group 98: marked-successors 
    -- CP-element group 98: 	37 
    -- CP-element group 98: 	96 
    -- CP-element group 98:  members (3) 
      -- CP-element group 98: 	 assign_stmt_97_to_assign_stmt_1138/slice_182_sample_completed_
      -- CP-element group 98: 	 assign_stmt_97_to_assign_stmt_1138/slice_182_Sample/$exit
      -- CP-element group 98: 	 assign_stmt_97_to_assign_stmt_1138/slice_182_Sample/ra
      -- 
    ra_910_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_182_inst_ack_0, ack => maxPool4_CP_346_elements(98)); -- 
    -- CP-element group 99:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	97 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	357 
    -- CP-element group 99: marked-successors 
    -- CP-element group 99: 	97 
    -- CP-element group 99:  members (3) 
      -- CP-element group 99: 	 assign_stmt_97_to_assign_stmt_1138/slice_182_update_completed_
      -- CP-element group 99: 	 assign_stmt_97_to_assign_stmt_1138/slice_182_Update/$exit
      -- CP-element group 99: 	 assign_stmt_97_to_assign_stmt_1138/slice_182_Update/ca
      -- 
    ca_915_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_182_inst_ack_1, ack => maxPool4_CP_346_elements(99)); -- 
    -- CP-element group 100:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	39 
    -- CP-element group 100: marked-predecessors 
    -- CP-element group 100: 	102 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	102 
    -- CP-element group 100:  members (3) 
      -- CP-element group 100: 	 assign_stmt_97_to_assign_stmt_1138/slice_186_sample_start_
      -- CP-element group 100: 	 assign_stmt_97_to_assign_stmt_1138/slice_186_Sample/$entry
      -- CP-element group 100: 	 assign_stmt_97_to_assign_stmt_1138/slice_186_Sample/rr
      -- 
    rr_923_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_923_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(100), ack => slice_186_inst_req_0); -- 
    maxPool4_cp_element_group_100: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_100"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(39) & maxPool4_CP_346_elements(102);
      gj_maxPool4_cp_element_group_100 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(100), clk => clk, reset => reset); --
    end block;
    -- CP-element group 101:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: marked-predecessors 
    -- CP-element group 101: 	103 
    -- CP-element group 101: 	378 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	103 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 assign_stmt_97_to_assign_stmt_1138/slice_186_update_start_
      -- CP-element group 101: 	 assign_stmt_97_to_assign_stmt_1138/slice_186_Update/$entry
      -- CP-element group 101: 	 assign_stmt_97_to_assign_stmt_1138/slice_186_Update/cr
      -- 
    cr_928_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_928_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(101), ack => slice_186_inst_req_1); -- 
    maxPool4_cp_element_group_101: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_101"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(103) & maxPool4_CP_346_elements(378);
      gj_maxPool4_cp_element_group_101 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(101), clk => clk, reset => reset); --
    end block;
    -- CP-element group 102:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	100 
    -- CP-element group 102: successors 
    -- CP-element group 102: marked-successors 
    -- CP-element group 102: 	37 
    -- CP-element group 102: 	100 
    -- CP-element group 102:  members (3) 
      -- CP-element group 102: 	 assign_stmt_97_to_assign_stmt_1138/slice_186_sample_completed_
      -- CP-element group 102: 	 assign_stmt_97_to_assign_stmt_1138/slice_186_Sample/$exit
      -- CP-element group 102: 	 assign_stmt_97_to_assign_stmt_1138/slice_186_Sample/ra
      -- 
    ra_924_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_186_inst_ack_0, ack => maxPool4_CP_346_elements(102)); -- 
    -- CP-element group 103:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	101 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	376 
    -- CP-element group 103: marked-successors 
    -- CP-element group 103: 	101 
    -- CP-element group 103:  members (3) 
      -- CP-element group 103: 	 assign_stmt_97_to_assign_stmt_1138/slice_186_update_completed_
      -- CP-element group 103: 	 assign_stmt_97_to_assign_stmt_1138/slice_186_Update/$exit
      -- CP-element group 103: 	 assign_stmt_97_to_assign_stmt_1138/slice_186_Update/ca
      -- 
    ca_929_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_186_inst_ack_1, ack => maxPool4_CP_346_elements(103)); -- 
    -- CP-element group 104:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	39 
    -- CP-element group 104: marked-predecessors 
    -- CP-element group 104: 	106 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	106 
    -- CP-element group 104:  members (3) 
      -- CP-element group 104: 	 assign_stmt_97_to_assign_stmt_1138/slice_190_sample_start_
      -- CP-element group 104: 	 assign_stmt_97_to_assign_stmt_1138/slice_190_Sample/$entry
      -- CP-element group 104: 	 assign_stmt_97_to_assign_stmt_1138/slice_190_Sample/rr
      -- 
    rr_937_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_937_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(104), ack => slice_190_inst_req_0); -- 
    maxPool4_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(39) & maxPool4_CP_346_elements(106);
      gj_maxPool4_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: marked-predecessors 
    -- CP-element group 105: 	107 
    -- CP-element group 105: 	378 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	107 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 assign_stmt_97_to_assign_stmt_1138/slice_190_update_start_
      -- CP-element group 105: 	 assign_stmt_97_to_assign_stmt_1138/slice_190_Update/$entry
      -- CP-element group 105: 	 assign_stmt_97_to_assign_stmt_1138/slice_190_Update/cr
      -- 
    cr_942_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_942_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(105), ack => slice_190_inst_req_1); -- 
    maxPool4_cp_element_group_105: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_105"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(107) & maxPool4_CP_346_elements(378);
      gj_maxPool4_cp_element_group_105 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(105), clk => clk, reset => reset); --
    end block;
    -- CP-element group 106:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	104 
    -- CP-element group 106: successors 
    -- CP-element group 106: marked-successors 
    -- CP-element group 106: 	37 
    -- CP-element group 106: 	104 
    -- CP-element group 106:  members (3) 
      -- CP-element group 106: 	 assign_stmt_97_to_assign_stmt_1138/slice_190_sample_completed_
      -- CP-element group 106: 	 assign_stmt_97_to_assign_stmt_1138/slice_190_Sample/$exit
      -- CP-element group 106: 	 assign_stmt_97_to_assign_stmt_1138/slice_190_Sample/ra
      -- 
    ra_938_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_190_inst_ack_0, ack => maxPool4_CP_346_elements(106)); -- 
    -- CP-element group 107:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	105 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	376 
    -- CP-element group 107: marked-successors 
    -- CP-element group 107: 	105 
    -- CP-element group 107:  members (3) 
      -- CP-element group 107: 	 assign_stmt_97_to_assign_stmt_1138/slice_190_update_completed_
      -- CP-element group 107: 	 assign_stmt_97_to_assign_stmt_1138/slice_190_Update/$exit
      -- CP-element group 107: 	 assign_stmt_97_to_assign_stmt_1138/slice_190_Update/ca
      -- 
    ca_943_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_190_inst_ack_1, ack => maxPool4_CP_346_elements(107)); -- 
    -- CP-element group 108:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	39 
    -- CP-element group 108: marked-predecessors 
    -- CP-element group 108: 	110 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	110 
    -- CP-element group 108:  members (3) 
      -- CP-element group 108: 	 assign_stmt_97_to_assign_stmt_1138/slice_194_sample_start_
      -- CP-element group 108: 	 assign_stmt_97_to_assign_stmt_1138/slice_194_Sample/$entry
      -- CP-element group 108: 	 assign_stmt_97_to_assign_stmt_1138/slice_194_Sample/rr
      -- 
    rr_951_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_951_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(108), ack => slice_194_inst_req_0); -- 
    maxPool4_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(39) & maxPool4_CP_346_elements(110);
      gj_maxPool4_cp_element_group_108 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: marked-predecessors 
    -- CP-element group 109: 	111 
    -- CP-element group 109: 	378 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 assign_stmt_97_to_assign_stmt_1138/slice_194_update_start_
      -- CP-element group 109: 	 assign_stmt_97_to_assign_stmt_1138/slice_194_Update/$entry
      -- CP-element group 109: 	 assign_stmt_97_to_assign_stmt_1138/slice_194_Update/cr
      -- 
    cr_956_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_956_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(109), ack => slice_194_inst_req_1); -- 
    maxPool4_cp_element_group_109: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_109"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(111) & maxPool4_CP_346_elements(378);
      gj_maxPool4_cp_element_group_109 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(109), clk => clk, reset => reset); --
    end block;
    -- CP-element group 110:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	108 
    -- CP-element group 110: successors 
    -- CP-element group 110: marked-successors 
    -- CP-element group 110: 	37 
    -- CP-element group 110: 	108 
    -- CP-element group 110:  members (3) 
      -- CP-element group 110: 	 assign_stmt_97_to_assign_stmt_1138/slice_194_sample_completed_
      -- CP-element group 110: 	 assign_stmt_97_to_assign_stmt_1138/slice_194_Sample/$exit
      -- CP-element group 110: 	 assign_stmt_97_to_assign_stmt_1138/slice_194_Sample/ra
      -- 
    ra_952_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_194_inst_ack_0, ack => maxPool4_CP_346_elements(110)); -- 
    -- CP-element group 111:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	376 
    -- CP-element group 111: marked-successors 
    -- CP-element group 111: 	109 
    -- CP-element group 111:  members (3) 
      -- CP-element group 111: 	 assign_stmt_97_to_assign_stmt_1138/slice_194_update_completed_
      -- CP-element group 111: 	 assign_stmt_97_to_assign_stmt_1138/slice_194_Update/$exit
      -- CP-element group 111: 	 assign_stmt_97_to_assign_stmt_1138/slice_194_Update/ca
      -- 
    ca_957_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_194_inst_ack_1, ack => maxPool4_CP_346_elements(111)); -- 
    -- CP-element group 112:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	39 
    -- CP-element group 112: marked-predecessors 
    -- CP-element group 112: 	114 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	114 
    -- CP-element group 112:  members (3) 
      -- CP-element group 112: 	 assign_stmt_97_to_assign_stmt_1138/slice_198_sample_start_
      -- CP-element group 112: 	 assign_stmt_97_to_assign_stmt_1138/slice_198_Sample/$entry
      -- CP-element group 112: 	 assign_stmt_97_to_assign_stmt_1138/slice_198_Sample/rr
      -- 
    rr_965_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_965_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(112), ack => slice_198_inst_req_0); -- 
    maxPool4_cp_element_group_112: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_112"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(39) & maxPool4_CP_346_elements(114);
      gj_maxPool4_cp_element_group_112 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(112), clk => clk, reset => reset); --
    end block;
    -- CP-element group 113:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: marked-predecessors 
    -- CP-element group 113: 	115 
    -- CP-element group 113: 	378 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 assign_stmt_97_to_assign_stmt_1138/slice_198_update_start_
      -- CP-element group 113: 	 assign_stmt_97_to_assign_stmt_1138/slice_198_Update/$entry
      -- CP-element group 113: 	 assign_stmt_97_to_assign_stmt_1138/slice_198_Update/cr
      -- 
    cr_970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(113), ack => slice_198_inst_req_1); -- 
    maxPool4_cp_element_group_113: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_113"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(115) & maxPool4_CP_346_elements(378);
      gj_maxPool4_cp_element_group_113 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(113), clk => clk, reset => reset); --
    end block;
    -- CP-element group 114:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	112 
    -- CP-element group 114: successors 
    -- CP-element group 114: marked-successors 
    -- CP-element group 114: 	37 
    -- CP-element group 114: 	112 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 assign_stmt_97_to_assign_stmt_1138/slice_198_sample_completed_
      -- CP-element group 114: 	 assign_stmt_97_to_assign_stmt_1138/slice_198_Sample/$exit
      -- CP-element group 114: 	 assign_stmt_97_to_assign_stmt_1138/slice_198_Sample/ra
      -- 
    ra_966_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_198_inst_ack_0, ack => maxPool4_CP_346_elements(114)); -- 
    -- CP-element group 115:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	376 
    -- CP-element group 115: marked-successors 
    -- CP-element group 115: 	113 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 assign_stmt_97_to_assign_stmt_1138/slice_198_update_completed_
      -- CP-element group 115: 	 assign_stmt_97_to_assign_stmt_1138/slice_198_Update/$exit
      -- CP-element group 115: 	 assign_stmt_97_to_assign_stmt_1138/slice_198_Update/ca
      -- 
    ca_971_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_198_inst_ack_1, ack => maxPool4_CP_346_elements(115)); -- 
    -- CP-element group 116:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	43 
    -- CP-element group 116: marked-predecessors 
    -- CP-element group 116: 	118 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	118 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 assign_stmt_97_to_assign_stmt_1138/slice_202_sample_start_
      -- CP-element group 116: 	 assign_stmt_97_to_assign_stmt_1138/slice_202_Sample/$entry
      -- CP-element group 116: 	 assign_stmt_97_to_assign_stmt_1138/slice_202_Sample/rr
      -- 
    rr_979_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_979_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(116), ack => slice_202_inst_req_0); -- 
    maxPool4_cp_element_group_116: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_116"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(43) & maxPool4_CP_346_elements(118);
      gj_maxPool4_cp_element_group_116 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(116), clk => clk, reset => reset); --
    end block;
    -- CP-element group 117:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: marked-predecessors 
    -- CP-element group 117: 	119 
    -- CP-element group 117: 	321 
    -- CP-element group 117: 	386 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	119 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 assign_stmt_97_to_assign_stmt_1138/slice_202_update_start_
      -- CP-element group 117: 	 assign_stmt_97_to_assign_stmt_1138/slice_202_Update/$entry
      -- CP-element group 117: 	 assign_stmt_97_to_assign_stmt_1138/slice_202_Update/cr
      -- 
    cr_984_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_984_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(117), ack => slice_202_inst_req_1); -- 
    maxPool4_cp_element_group_117: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_117"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(119) & maxPool4_CP_346_elements(321) & maxPool4_CP_346_elements(386);
      gj_maxPool4_cp_element_group_117 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(117), clk => clk, reset => reset); --
    end block;
    -- CP-element group 118:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	116 
    -- CP-element group 118: successors 
    -- CP-element group 118: marked-successors 
    -- CP-element group 118: 	41 
    -- CP-element group 118: 	116 
    -- CP-element group 118:  members (3) 
      -- CP-element group 118: 	 assign_stmt_97_to_assign_stmt_1138/slice_202_sample_completed_
      -- CP-element group 118: 	 assign_stmt_97_to_assign_stmt_1138/slice_202_Sample/$exit
      -- CP-element group 118: 	 assign_stmt_97_to_assign_stmt_1138/slice_202_Sample/ra
      -- 
    ra_980_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_202_inst_ack_0, ack => maxPool4_CP_346_elements(118)); -- 
    -- CP-element group 119:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	117 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	319 
    -- CP-element group 119: 	384 
    -- CP-element group 119: marked-successors 
    -- CP-element group 119: 	117 
    -- CP-element group 119:  members (3) 
      -- CP-element group 119: 	 assign_stmt_97_to_assign_stmt_1138/slice_202_update_completed_
      -- CP-element group 119: 	 assign_stmt_97_to_assign_stmt_1138/slice_202_Update/$exit
      -- CP-element group 119: 	 assign_stmt_97_to_assign_stmt_1138/slice_202_Update/ca
      -- 
    ca_985_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_202_inst_ack_1, ack => maxPool4_CP_346_elements(119)); -- 
    -- CP-element group 120:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	43 
    -- CP-element group 120: marked-predecessors 
    -- CP-element group 120: 	122 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	122 
    -- CP-element group 120:  members (3) 
      -- CP-element group 120: 	 assign_stmt_97_to_assign_stmt_1138/slice_206_sample_start_
      -- CP-element group 120: 	 assign_stmt_97_to_assign_stmt_1138/slice_206_Sample/$entry
      -- CP-element group 120: 	 assign_stmt_97_to_assign_stmt_1138/slice_206_Sample/rr
      -- 
    rr_993_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_993_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(120), ack => slice_206_inst_req_0); -- 
    maxPool4_cp_element_group_120: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_120"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(43) & maxPool4_CP_346_elements(122);
      gj_maxPool4_cp_element_group_120 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(120), clk => clk, reset => reset); --
    end block;
    -- CP-element group 121:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: marked-predecessors 
    -- CP-element group 121: 	123 
    -- CP-element group 121: 	321 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	123 
    -- CP-element group 121:  members (3) 
      -- CP-element group 121: 	 assign_stmt_97_to_assign_stmt_1138/slice_206_Update/cr
      -- CP-element group 121: 	 assign_stmt_97_to_assign_stmt_1138/slice_206_update_start_
      -- CP-element group 121: 	 assign_stmt_97_to_assign_stmt_1138/slice_206_Update/$entry
      -- 
    cr_998_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_998_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(121), ack => slice_206_inst_req_1); -- 
    maxPool4_cp_element_group_121: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_121"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(123) & maxPool4_CP_346_elements(321);
      gj_maxPool4_cp_element_group_121 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(121), clk => clk, reset => reset); --
    end block;
    -- CP-element group 122:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	120 
    -- CP-element group 122: successors 
    -- CP-element group 122: marked-successors 
    -- CP-element group 122: 	41 
    -- CP-element group 122: 	120 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 assign_stmt_97_to_assign_stmt_1138/slice_206_sample_completed_
      -- CP-element group 122: 	 assign_stmt_97_to_assign_stmt_1138/slice_206_Sample/$exit
      -- CP-element group 122: 	 assign_stmt_97_to_assign_stmt_1138/slice_206_Sample/ra
      -- 
    ra_994_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_206_inst_ack_0, ack => maxPool4_CP_346_elements(122)); -- 
    -- CP-element group 123:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	121 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	319 
    -- CP-element group 123: marked-successors 
    -- CP-element group 123: 	121 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 assign_stmt_97_to_assign_stmt_1138/slice_206_Update/ca
      -- CP-element group 123: 	 assign_stmt_97_to_assign_stmt_1138/slice_206_update_completed_
      -- CP-element group 123: 	 assign_stmt_97_to_assign_stmt_1138/slice_206_Update/$exit
      -- 
    ca_999_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_206_inst_ack_1, ack => maxPool4_CP_346_elements(123)); -- 
    -- CP-element group 124:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	43 
    -- CP-element group 124: marked-predecessors 
    -- CP-element group 124: 	126 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	126 
    -- CP-element group 124:  members (3) 
      -- CP-element group 124: 	 assign_stmt_97_to_assign_stmt_1138/slice_210_Sample/$entry
      -- CP-element group 124: 	 assign_stmt_97_to_assign_stmt_1138/slice_210_Sample/rr
      -- CP-element group 124: 	 assign_stmt_97_to_assign_stmt_1138/slice_210_sample_start_
      -- 
    rr_1007_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1007_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(124), ack => slice_210_inst_req_0); -- 
    maxPool4_cp_element_group_124: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_124"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(43) & maxPool4_CP_346_elements(126);
      gj_maxPool4_cp_element_group_124 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(124), clk => clk, reset => reset); --
    end block;
    -- CP-element group 125:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: marked-predecessors 
    -- CP-element group 125: 	127 
    -- CP-element group 125: 	321 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	127 
    -- CP-element group 125:  members (3) 
      -- CP-element group 125: 	 assign_stmt_97_to_assign_stmt_1138/slice_210_Update/$entry
      -- CP-element group 125: 	 assign_stmt_97_to_assign_stmt_1138/slice_210_Update/cr
      -- CP-element group 125: 	 assign_stmt_97_to_assign_stmt_1138/slice_210_update_start_
      -- 
    cr_1012_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1012_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(125), ack => slice_210_inst_req_1); -- 
    maxPool4_cp_element_group_125: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_125"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(127) & maxPool4_CP_346_elements(321);
      gj_maxPool4_cp_element_group_125 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(125), clk => clk, reset => reset); --
    end block;
    -- CP-element group 126:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	124 
    -- CP-element group 126: successors 
    -- CP-element group 126: marked-successors 
    -- CP-element group 126: 	41 
    -- CP-element group 126: 	124 
    -- CP-element group 126:  members (3) 
      -- CP-element group 126: 	 assign_stmt_97_to_assign_stmt_1138/slice_210_Sample/ra
      -- CP-element group 126: 	 assign_stmt_97_to_assign_stmt_1138/slice_210_Sample/$exit
      -- CP-element group 126: 	 assign_stmt_97_to_assign_stmt_1138/slice_210_sample_completed_
      -- 
    ra_1008_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_210_inst_ack_0, ack => maxPool4_CP_346_elements(126)); -- 
    -- CP-element group 127:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	125 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	319 
    -- CP-element group 127: marked-successors 
    -- CP-element group 127: 	125 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 assign_stmt_97_to_assign_stmt_1138/slice_210_update_completed_
      -- CP-element group 127: 	 assign_stmt_97_to_assign_stmt_1138/slice_210_Update/ca
      -- CP-element group 127: 	 assign_stmt_97_to_assign_stmt_1138/slice_210_Update/$exit
      -- 
    ca_1013_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_210_inst_ack_1, ack => maxPool4_CP_346_elements(127)); -- 
    -- CP-element group 128:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	43 
    -- CP-element group 128: marked-predecessors 
    -- CP-element group 128: 	130 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	130 
    -- CP-element group 128:  members (3) 
      -- CP-element group 128: 	 assign_stmt_97_to_assign_stmt_1138/slice_214_Sample/rr
      -- CP-element group 128: 	 assign_stmt_97_to_assign_stmt_1138/slice_214_Sample/$entry
      -- CP-element group 128: 	 assign_stmt_97_to_assign_stmt_1138/slice_214_sample_start_
      -- 
    rr_1021_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1021_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(128), ack => slice_214_inst_req_0); -- 
    maxPool4_cp_element_group_128: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_128"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(43) & maxPool4_CP_346_elements(130);
      gj_maxPool4_cp_element_group_128 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(128), clk => clk, reset => reset); --
    end block;
    -- CP-element group 129:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: marked-predecessors 
    -- CP-element group 129: 	131 
    -- CP-element group 129: 	321 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	131 
    -- CP-element group 129:  members (3) 
      -- CP-element group 129: 	 assign_stmt_97_to_assign_stmt_1138/slice_214_Update/$entry
      -- CP-element group 129: 	 assign_stmt_97_to_assign_stmt_1138/slice_214_update_start_
      -- CP-element group 129: 	 assign_stmt_97_to_assign_stmt_1138/slice_214_Update/cr
      -- 
    cr_1026_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1026_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(129), ack => slice_214_inst_req_1); -- 
    maxPool4_cp_element_group_129: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_129"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(131) & maxPool4_CP_346_elements(321);
      gj_maxPool4_cp_element_group_129 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(129), clk => clk, reset => reset); --
    end block;
    -- CP-element group 130:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	128 
    -- CP-element group 130: successors 
    -- CP-element group 130: marked-successors 
    -- CP-element group 130: 	41 
    -- CP-element group 130: 	128 
    -- CP-element group 130:  members (3) 
      -- CP-element group 130: 	 assign_stmt_97_to_assign_stmt_1138/slice_214_Sample/ra
      -- CP-element group 130: 	 assign_stmt_97_to_assign_stmt_1138/slice_214_Sample/$exit
      -- CP-element group 130: 	 assign_stmt_97_to_assign_stmt_1138/slice_214_sample_completed_
      -- 
    ra_1022_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_214_inst_ack_0, ack => maxPool4_CP_346_elements(130)); -- 
    -- CP-element group 131:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	129 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	319 
    -- CP-element group 131: marked-successors 
    -- CP-element group 131: 	129 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 assign_stmt_97_to_assign_stmt_1138/slice_214_update_completed_
      -- CP-element group 131: 	 assign_stmt_97_to_assign_stmt_1138/slice_214_Update/ca
      -- CP-element group 131: 	 assign_stmt_97_to_assign_stmt_1138/slice_214_Update/$exit
      -- 
    ca_1027_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_214_inst_ack_1, ack => maxPool4_CP_346_elements(131)); -- 
    -- CP-element group 132:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	43 
    -- CP-element group 132: marked-predecessors 
    -- CP-element group 132: 	134 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	134 
    -- CP-element group 132:  members (3) 
      -- CP-element group 132: 	 assign_stmt_97_to_assign_stmt_1138/slice_218_Sample/rr
      -- CP-element group 132: 	 assign_stmt_97_to_assign_stmt_1138/slice_218_Sample/$entry
      -- CP-element group 132: 	 assign_stmt_97_to_assign_stmt_1138/slice_218_sample_start_
      -- 
    rr_1035_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1035_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(132), ack => slice_218_inst_req_0); -- 
    maxPool4_cp_element_group_132: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_132"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(43) & maxPool4_CP_346_elements(134);
      gj_maxPool4_cp_element_group_132 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(132), clk => clk, reset => reset); --
    end block;
    -- CP-element group 133:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: marked-predecessors 
    -- CP-element group 133: 	135 
    -- CP-element group 133: 	340 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	135 
    -- CP-element group 133:  members (3) 
      -- CP-element group 133: 	 assign_stmt_97_to_assign_stmt_1138/slice_218_Update/cr
      -- CP-element group 133: 	 assign_stmt_97_to_assign_stmt_1138/slice_218_Update/$entry
      -- CP-element group 133: 	 assign_stmt_97_to_assign_stmt_1138/slice_218_update_start_
      -- 
    cr_1040_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1040_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(133), ack => slice_218_inst_req_1); -- 
    maxPool4_cp_element_group_133: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_133"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(135) & maxPool4_CP_346_elements(340);
      gj_maxPool4_cp_element_group_133 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(133), clk => clk, reset => reset); --
    end block;
    -- CP-element group 134:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	132 
    -- CP-element group 134: successors 
    -- CP-element group 134: marked-successors 
    -- CP-element group 134: 	41 
    -- CP-element group 134: 	132 
    -- CP-element group 134:  members (3) 
      -- CP-element group 134: 	 assign_stmt_97_to_assign_stmt_1138/slice_218_Sample/$exit
      -- CP-element group 134: 	 assign_stmt_97_to_assign_stmt_1138/slice_218_Sample/ra
      -- CP-element group 134: 	 assign_stmt_97_to_assign_stmt_1138/slice_218_sample_completed_
      -- 
    ra_1036_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_218_inst_ack_0, ack => maxPool4_CP_346_elements(134)); -- 
    -- CP-element group 135:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	133 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	338 
    -- CP-element group 135: marked-successors 
    -- CP-element group 135: 	133 
    -- CP-element group 135:  members (3) 
      -- CP-element group 135: 	 assign_stmt_97_to_assign_stmt_1138/slice_218_Update/ca
      -- CP-element group 135: 	 assign_stmt_97_to_assign_stmt_1138/slice_218_Update/$exit
      -- CP-element group 135: 	 assign_stmt_97_to_assign_stmt_1138/slice_218_update_completed_
      -- 
    ca_1041_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_218_inst_ack_1, ack => maxPool4_CP_346_elements(135)); -- 
    -- CP-element group 136:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	43 
    -- CP-element group 136: marked-predecessors 
    -- CP-element group 136: 	138 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	138 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 assign_stmt_97_to_assign_stmt_1138/slice_222_Sample/rr
      -- CP-element group 136: 	 assign_stmt_97_to_assign_stmt_1138/slice_222_Sample/$entry
      -- CP-element group 136: 	 assign_stmt_97_to_assign_stmt_1138/slice_222_sample_start_
      -- 
    rr_1049_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1049_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(136), ack => slice_222_inst_req_0); -- 
    maxPool4_cp_element_group_136: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_136"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(43) & maxPool4_CP_346_elements(138);
      gj_maxPool4_cp_element_group_136 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(136), clk => clk, reset => reset); --
    end block;
    -- CP-element group 137:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: marked-predecessors 
    -- CP-element group 137: 	139 
    -- CP-element group 137: 	340 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	139 
    -- CP-element group 137:  members (3) 
      -- CP-element group 137: 	 assign_stmt_97_to_assign_stmt_1138/slice_222_Update/$entry
      -- CP-element group 137: 	 assign_stmt_97_to_assign_stmt_1138/slice_222_update_start_
      -- CP-element group 137: 	 assign_stmt_97_to_assign_stmt_1138/slice_222_Update/cr
      -- 
    cr_1054_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1054_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(137), ack => slice_222_inst_req_1); -- 
    maxPool4_cp_element_group_137: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_137"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(139) & maxPool4_CP_346_elements(340);
      gj_maxPool4_cp_element_group_137 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(137), clk => clk, reset => reset); --
    end block;
    -- CP-element group 138:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	136 
    -- CP-element group 138: successors 
    -- CP-element group 138: marked-successors 
    -- CP-element group 138: 	41 
    -- CP-element group 138: 	136 
    -- CP-element group 138:  members (3) 
      -- CP-element group 138: 	 assign_stmt_97_to_assign_stmt_1138/slice_222_Sample/ra
      -- CP-element group 138: 	 assign_stmt_97_to_assign_stmt_1138/slice_222_Sample/$exit
      -- CP-element group 138: 	 assign_stmt_97_to_assign_stmt_1138/slice_222_sample_completed_
      -- 
    ra_1050_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_222_inst_ack_0, ack => maxPool4_CP_346_elements(138)); -- 
    -- CP-element group 139:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	137 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	338 
    -- CP-element group 139: marked-successors 
    -- CP-element group 139: 	137 
    -- CP-element group 139:  members (3) 
      -- CP-element group 139: 	 assign_stmt_97_to_assign_stmt_1138/slice_222_Update/$exit
      -- CP-element group 139: 	 assign_stmt_97_to_assign_stmt_1138/slice_222_update_completed_
      -- CP-element group 139: 	 assign_stmt_97_to_assign_stmt_1138/slice_222_Update/ca
      -- 
    ca_1055_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_222_inst_ack_1, ack => maxPool4_CP_346_elements(139)); -- 
    -- CP-element group 140:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	43 
    -- CP-element group 140: marked-predecessors 
    -- CP-element group 140: 	142 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	142 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 assign_stmt_97_to_assign_stmt_1138/slice_226_Sample/rr
      -- CP-element group 140: 	 assign_stmt_97_to_assign_stmt_1138/slice_226_Sample/$entry
      -- CP-element group 140: 	 assign_stmt_97_to_assign_stmt_1138/slice_226_sample_start_
      -- 
    rr_1063_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1063_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(140), ack => slice_226_inst_req_0); -- 
    maxPool4_cp_element_group_140: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_140"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(43) & maxPool4_CP_346_elements(142);
      gj_maxPool4_cp_element_group_140 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(140), clk => clk, reset => reset); --
    end block;
    -- CP-element group 141:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: marked-predecessors 
    -- CP-element group 141: 	143 
    -- CP-element group 141: 	340 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	143 
    -- CP-element group 141:  members (3) 
      -- CP-element group 141: 	 assign_stmt_97_to_assign_stmt_1138/slice_226_Update/cr
      -- CP-element group 141: 	 assign_stmt_97_to_assign_stmt_1138/slice_226_Update/$entry
      -- CP-element group 141: 	 assign_stmt_97_to_assign_stmt_1138/slice_226_update_start_
      -- 
    cr_1068_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1068_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(141), ack => slice_226_inst_req_1); -- 
    maxPool4_cp_element_group_141: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_141"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(143) & maxPool4_CP_346_elements(340);
      gj_maxPool4_cp_element_group_141 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(141), clk => clk, reset => reset); --
    end block;
    -- CP-element group 142:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	140 
    -- CP-element group 142: successors 
    -- CP-element group 142: marked-successors 
    -- CP-element group 142: 	41 
    -- CP-element group 142: 	140 
    -- CP-element group 142:  members (3) 
      -- CP-element group 142: 	 assign_stmt_97_to_assign_stmt_1138/slice_226_Sample/ra
      -- CP-element group 142: 	 assign_stmt_97_to_assign_stmt_1138/slice_226_Sample/$exit
      -- CP-element group 142: 	 assign_stmt_97_to_assign_stmt_1138/slice_226_sample_completed_
      -- 
    ra_1064_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_226_inst_ack_0, ack => maxPool4_CP_346_elements(142)); -- 
    -- CP-element group 143:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	141 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	338 
    -- CP-element group 143: marked-successors 
    -- CP-element group 143: 	141 
    -- CP-element group 143:  members (3) 
      -- CP-element group 143: 	 assign_stmt_97_to_assign_stmt_1138/slice_226_Update/$exit
      -- CP-element group 143: 	 assign_stmt_97_to_assign_stmt_1138/slice_226_update_completed_
      -- CP-element group 143: 	 assign_stmt_97_to_assign_stmt_1138/slice_226_Update/ca
      -- 
    ca_1069_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_226_inst_ack_1, ack => maxPool4_CP_346_elements(143)); -- 
    -- CP-element group 144:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	43 
    -- CP-element group 144: marked-predecessors 
    -- CP-element group 144: 	146 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	146 
    -- CP-element group 144:  members (3) 
      -- CP-element group 144: 	 assign_stmt_97_to_assign_stmt_1138/slice_230_Sample/rr
      -- CP-element group 144: 	 assign_stmt_97_to_assign_stmt_1138/slice_230_Sample/$entry
      -- CP-element group 144: 	 assign_stmt_97_to_assign_stmt_1138/slice_230_sample_start_
      -- 
    rr_1077_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1077_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(144), ack => slice_230_inst_req_0); -- 
    maxPool4_cp_element_group_144: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_144"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(43) & maxPool4_CP_346_elements(146);
      gj_maxPool4_cp_element_group_144 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(144), clk => clk, reset => reset); --
    end block;
    -- CP-element group 145:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: marked-predecessors 
    -- CP-element group 145: 	147 
    -- CP-element group 145: 	340 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	147 
    -- CP-element group 145:  members (3) 
      -- CP-element group 145: 	 assign_stmt_97_to_assign_stmt_1138/slice_230_Update/cr
      -- CP-element group 145: 	 assign_stmt_97_to_assign_stmt_1138/slice_230_Update/$entry
      -- CP-element group 145: 	 assign_stmt_97_to_assign_stmt_1138/slice_230_update_start_
      -- 
    cr_1082_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1082_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(145), ack => slice_230_inst_req_1); -- 
    maxPool4_cp_element_group_145: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_145"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(147) & maxPool4_CP_346_elements(340);
      gj_maxPool4_cp_element_group_145 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(145), clk => clk, reset => reset); --
    end block;
    -- CP-element group 146:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	144 
    -- CP-element group 146: successors 
    -- CP-element group 146: marked-successors 
    -- CP-element group 146: 	41 
    -- CP-element group 146: 	144 
    -- CP-element group 146:  members (3) 
      -- CP-element group 146: 	 assign_stmt_97_to_assign_stmt_1138/slice_230_Sample/ra
      -- CP-element group 146: 	 assign_stmt_97_to_assign_stmt_1138/slice_230_Sample/$exit
      -- CP-element group 146: 	 assign_stmt_97_to_assign_stmt_1138/slice_230_sample_completed_
      -- 
    ra_1078_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_230_inst_ack_0, ack => maxPool4_CP_346_elements(146)); -- 
    -- CP-element group 147:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	145 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	338 
    -- CP-element group 147: marked-successors 
    -- CP-element group 147: 	145 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 assign_stmt_97_to_assign_stmt_1138/slice_230_Update/ca
      -- CP-element group 147: 	 assign_stmt_97_to_assign_stmt_1138/slice_230_Update/$exit
      -- CP-element group 147: 	 assign_stmt_97_to_assign_stmt_1138/slice_230_update_completed_
      -- 
    ca_1083_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_230_inst_ack_1, ack => maxPool4_CP_346_elements(147)); -- 
    -- CP-element group 148:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	43 
    -- CP-element group 148: marked-predecessors 
    -- CP-element group 148: 	150 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	150 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 assign_stmt_97_to_assign_stmt_1138/slice_234_Sample/rr
      -- CP-element group 148: 	 assign_stmt_97_to_assign_stmt_1138/slice_234_Sample/$entry
      -- CP-element group 148: 	 assign_stmt_97_to_assign_stmt_1138/slice_234_sample_start_
      -- 
    rr_1091_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1091_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(148), ack => slice_234_inst_req_0); -- 
    maxPool4_cp_element_group_148: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_148"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(43) & maxPool4_CP_346_elements(150);
      gj_maxPool4_cp_element_group_148 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(148), clk => clk, reset => reset); --
    end block;
    -- CP-element group 149:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: marked-predecessors 
    -- CP-element group 149: 	151 
    -- CP-element group 149: 	359 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	151 
    -- CP-element group 149:  members (3) 
      -- CP-element group 149: 	 assign_stmt_97_to_assign_stmt_1138/slice_234_Update/cr
      -- CP-element group 149: 	 assign_stmt_97_to_assign_stmt_1138/slice_234_Update/$entry
      -- CP-element group 149: 	 assign_stmt_97_to_assign_stmt_1138/slice_234_update_start_
      -- 
    cr_1096_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1096_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(149), ack => slice_234_inst_req_1); -- 
    maxPool4_cp_element_group_149: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_149"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(151) & maxPool4_CP_346_elements(359);
      gj_maxPool4_cp_element_group_149 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(149), clk => clk, reset => reset); --
    end block;
    -- CP-element group 150:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	148 
    -- CP-element group 150: successors 
    -- CP-element group 150: marked-successors 
    -- CP-element group 150: 	41 
    -- CP-element group 150: 	148 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 assign_stmt_97_to_assign_stmt_1138/slice_234_Sample/ra
      -- CP-element group 150: 	 assign_stmt_97_to_assign_stmt_1138/slice_234_Sample/$exit
      -- CP-element group 150: 	 assign_stmt_97_to_assign_stmt_1138/slice_234_sample_completed_
      -- 
    ra_1092_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_234_inst_ack_0, ack => maxPool4_CP_346_elements(150)); -- 
    -- CP-element group 151:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	149 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	357 
    -- CP-element group 151: marked-successors 
    -- CP-element group 151: 	149 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 assign_stmt_97_to_assign_stmt_1138/slice_234_Update/ca
      -- CP-element group 151: 	 assign_stmt_97_to_assign_stmt_1138/slice_234_Update/$exit
      -- CP-element group 151: 	 assign_stmt_97_to_assign_stmt_1138/slice_234_update_completed_
      -- 
    ca_1097_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_234_inst_ack_1, ack => maxPool4_CP_346_elements(151)); -- 
    -- CP-element group 152:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	43 
    -- CP-element group 152: marked-predecessors 
    -- CP-element group 152: 	154 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	154 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 assign_stmt_97_to_assign_stmt_1138/slice_238_Sample/rr
      -- CP-element group 152: 	 assign_stmt_97_to_assign_stmt_1138/slice_238_Sample/$entry
      -- CP-element group 152: 	 assign_stmt_97_to_assign_stmt_1138/slice_238_sample_start_
      -- 
    rr_1105_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1105_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(152), ack => slice_238_inst_req_0); -- 
    maxPool4_cp_element_group_152: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_152"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(43) & maxPool4_CP_346_elements(154);
      gj_maxPool4_cp_element_group_152 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(152), clk => clk, reset => reset); --
    end block;
    -- CP-element group 153:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: marked-predecessors 
    -- CP-element group 153: 	155 
    -- CP-element group 153: 	359 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	155 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 assign_stmt_97_to_assign_stmt_1138/slice_238_Update/cr
      -- CP-element group 153: 	 assign_stmt_97_to_assign_stmt_1138/slice_238_Update/$entry
      -- CP-element group 153: 	 assign_stmt_97_to_assign_stmt_1138/slice_238_update_start_
      -- 
    cr_1110_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1110_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(153), ack => slice_238_inst_req_1); -- 
    maxPool4_cp_element_group_153: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_153"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(155) & maxPool4_CP_346_elements(359);
      gj_maxPool4_cp_element_group_153 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(153), clk => clk, reset => reset); --
    end block;
    -- CP-element group 154:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	152 
    -- CP-element group 154: successors 
    -- CP-element group 154: marked-successors 
    -- CP-element group 154: 	41 
    -- CP-element group 154: 	152 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 assign_stmt_97_to_assign_stmt_1138/slice_238_Sample/ra
      -- CP-element group 154: 	 assign_stmt_97_to_assign_stmt_1138/slice_238_Sample/$exit
      -- CP-element group 154: 	 assign_stmt_97_to_assign_stmt_1138/slice_238_sample_completed_
      -- 
    ra_1106_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_238_inst_ack_0, ack => maxPool4_CP_346_elements(154)); -- 
    -- CP-element group 155:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	153 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	357 
    -- CP-element group 155: marked-successors 
    -- CP-element group 155: 	153 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 assign_stmt_97_to_assign_stmt_1138/slice_238_Update/$exit
      -- CP-element group 155: 	 assign_stmt_97_to_assign_stmt_1138/slice_238_update_completed_
      -- CP-element group 155: 	 assign_stmt_97_to_assign_stmt_1138/slice_238_Update/ca
      -- 
    ca_1111_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_238_inst_ack_1, ack => maxPool4_CP_346_elements(155)); -- 
    -- CP-element group 156:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	43 
    -- CP-element group 156: marked-predecessors 
    -- CP-element group 156: 	158 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	158 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 assign_stmt_97_to_assign_stmt_1138/slice_242_sample_start_
      -- CP-element group 156: 	 assign_stmt_97_to_assign_stmt_1138/slice_242_Sample/rr
      -- CP-element group 156: 	 assign_stmt_97_to_assign_stmt_1138/slice_242_Sample/$entry
      -- 
    rr_1119_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1119_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(156), ack => slice_242_inst_req_0); -- 
    maxPool4_cp_element_group_156: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_156"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(43) & maxPool4_CP_346_elements(158);
      gj_maxPool4_cp_element_group_156 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(156), clk => clk, reset => reset); --
    end block;
    -- CP-element group 157:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: marked-predecessors 
    -- CP-element group 157: 	159 
    -- CP-element group 157: 	359 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	159 
    -- CP-element group 157:  members (3) 
      -- CP-element group 157: 	 assign_stmt_97_to_assign_stmt_1138/slice_242_update_start_
      -- CP-element group 157: 	 assign_stmt_97_to_assign_stmt_1138/slice_242_Update/cr
      -- CP-element group 157: 	 assign_stmt_97_to_assign_stmt_1138/slice_242_Update/$entry
      -- 
    cr_1124_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1124_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(157), ack => slice_242_inst_req_1); -- 
    maxPool4_cp_element_group_157: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_157"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(159) & maxPool4_CP_346_elements(359);
      gj_maxPool4_cp_element_group_157 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(157), clk => clk, reset => reset); --
    end block;
    -- CP-element group 158:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	156 
    -- CP-element group 158: successors 
    -- CP-element group 158: marked-successors 
    -- CP-element group 158: 	41 
    -- CP-element group 158: 	156 
    -- CP-element group 158:  members (3) 
      -- CP-element group 158: 	 assign_stmt_97_to_assign_stmt_1138/slice_242_sample_completed_
      -- CP-element group 158: 	 assign_stmt_97_to_assign_stmt_1138/slice_242_Sample/ra
      -- CP-element group 158: 	 assign_stmt_97_to_assign_stmt_1138/slice_242_Sample/$exit
      -- 
    ra_1120_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_242_inst_ack_0, ack => maxPool4_CP_346_elements(158)); -- 
    -- CP-element group 159:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	157 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	357 
    -- CP-element group 159: marked-successors 
    -- CP-element group 159: 	157 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 assign_stmt_97_to_assign_stmt_1138/slice_242_Update/ca
      -- CP-element group 159: 	 assign_stmt_97_to_assign_stmt_1138/slice_242_Update/$exit
      -- CP-element group 159: 	 assign_stmt_97_to_assign_stmt_1138/slice_242_update_completed_
      -- 
    ca_1125_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_242_inst_ack_1, ack => maxPool4_CP_346_elements(159)); -- 
    -- CP-element group 160:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	43 
    -- CP-element group 160: marked-predecessors 
    -- CP-element group 160: 	162 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	162 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 assign_stmt_97_to_assign_stmt_1138/slice_246_Sample/rr
      -- CP-element group 160: 	 assign_stmt_97_to_assign_stmt_1138/slice_246_Sample/$entry
      -- CP-element group 160: 	 assign_stmt_97_to_assign_stmt_1138/slice_246_sample_start_
      -- 
    rr_1133_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1133_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(160), ack => slice_246_inst_req_0); -- 
    maxPool4_cp_element_group_160: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_160"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(43) & maxPool4_CP_346_elements(162);
      gj_maxPool4_cp_element_group_160 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(160), clk => clk, reset => reset); --
    end block;
    -- CP-element group 161:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: marked-predecessors 
    -- CP-element group 161: 	163 
    -- CP-element group 161: 	359 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	163 
    -- CP-element group 161:  members (3) 
      -- CP-element group 161: 	 assign_stmt_97_to_assign_stmt_1138/slice_246_update_start_
      -- CP-element group 161: 	 assign_stmt_97_to_assign_stmt_1138/slice_246_Update/cr
      -- CP-element group 161: 	 assign_stmt_97_to_assign_stmt_1138/slice_246_Update/$entry
      -- 
    cr_1138_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1138_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(161), ack => slice_246_inst_req_1); -- 
    maxPool4_cp_element_group_161: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_161"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(163) & maxPool4_CP_346_elements(359);
      gj_maxPool4_cp_element_group_161 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(161), clk => clk, reset => reset); --
    end block;
    -- CP-element group 162:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	160 
    -- CP-element group 162: successors 
    -- CP-element group 162: marked-successors 
    -- CP-element group 162: 	41 
    -- CP-element group 162: 	160 
    -- CP-element group 162:  members (3) 
      -- CP-element group 162: 	 assign_stmt_97_to_assign_stmt_1138/slice_246_Sample/ra
      -- CP-element group 162: 	 assign_stmt_97_to_assign_stmt_1138/slice_246_Sample/$exit
      -- CP-element group 162: 	 assign_stmt_97_to_assign_stmt_1138/slice_246_sample_completed_
      -- 
    ra_1134_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_246_inst_ack_0, ack => maxPool4_CP_346_elements(162)); -- 
    -- CP-element group 163:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	161 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	357 
    -- CP-element group 163: marked-successors 
    -- CP-element group 163: 	161 
    -- CP-element group 163:  members (3) 
      -- CP-element group 163: 	 assign_stmt_97_to_assign_stmt_1138/slice_246_Update/ca
      -- CP-element group 163: 	 assign_stmt_97_to_assign_stmt_1138/slice_246_update_completed_
      -- CP-element group 163: 	 assign_stmt_97_to_assign_stmt_1138/slice_246_Update/$exit
      -- 
    ca_1139_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_246_inst_ack_1, ack => maxPool4_CP_346_elements(163)); -- 
    -- CP-element group 164:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	43 
    -- CP-element group 164: marked-predecessors 
    -- CP-element group 164: 	166 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	166 
    -- CP-element group 164:  members (3) 
      -- CP-element group 164: 	 assign_stmt_97_to_assign_stmt_1138/slice_250_sample_start_
      -- CP-element group 164: 	 assign_stmt_97_to_assign_stmt_1138/slice_250_Sample/rr
      -- CP-element group 164: 	 assign_stmt_97_to_assign_stmt_1138/slice_250_Sample/$entry
      -- 
    rr_1147_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1147_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(164), ack => slice_250_inst_req_0); -- 
    maxPool4_cp_element_group_164: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_164"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(43) & maxPool4_CP_346_elements(166);
      gj_maxPool4_cp_element_group_164 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(164), clk => clk, reset => reset); --
    end block;
    -- CP-element group 165:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: marked-predecessors 
    -- CP-element group 165: 	167 
    -- CP-element group 165: 	378 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	167 
    -- CP-element group 165:  members (3) 
      -- CP-element group 165: 	 assign_stmt_97_to_assign_stmt_1138/slice_250_update_start_
      -- CP-element group 165: 	 assign_stmt_97_to_assign_stmt_1138/slice_250_Update/cr
      -- CP-element group 165: 	 assign_stmt_97_to_assign_stmt_1138/slice_250_Update/$entry
      -- 
    cr_1152_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1152_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(165), ack => slice_250_inst_req_1); -- 
    maxPool4_cp_element_group_165: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_165"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(167) & maxPool4_CP_346_elements(378);
      gj_maxPool4_cp_element_group_165 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(165), clk => clk, reset => reset); --
    end block;
    -- CP-element group 166:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	164 
    -- CP-element group 166: successors 
    -- CP-element group 166: marked-successors 
    -- CP-element group 166: 	41 
    -- CP-element group 166: 	164 
    -- CP-element group 166:  members (3) 
      -- CP-element group 166: 	 assign_stmt_97_to_assign_stmt_1138/slice_250_Sample/ra
      -- CP-element group 166: 	 assign_stmt_97_to_assign_stmt_1138/slice_250_Sample/$exit
      -- CP-element group 166: 	 assign_stmt_97_to_assign_stmt_1138/slice_250_sample_completed_
      -- 
    ra_1148_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_250_inst_ack_0, ack => maxPool4_CP_346_elements(166)); -- 
    -- CP-element group 167:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	165 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	376 
    -- CP-element group 167: marked-successors 
    -- CP-element group 167: 	165 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 assign_stmt_97_to_assign_stmt_1138/slice_250_Update/ca
      -- CP-element group 167: 	 assign_stmt_97_to_assign_stmt_1138/slice_250_Update/$exit
      -- CP-element group 167: 	 assign_stmt_97_to_assign_stmt_1138/slice_250_update_completed_
      -- 
    ca_1153_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_250_inst_ack_1, ack => maxPool4_CP_346_elements(167)); -- 
    -- CP-element group 168:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	43 
    -- CP-element group 168: marked-predecessors 
    -- CP-element group 168: 	170 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	170 
    -- CP-element group 168:  members (3) 
      -- CP-element group 168: 	 assign_stmt_97_to_assign_stmt_1138/slice_254_sample_start_
      -- CP-element group 168: 	 assign_stmt_97_to_assign_stmt_1138/slice_254_Sample/$entry
      -- CP-element group 168: 	 assign_stmt_97_to_assign_stmt_1138/slice_254_Sample/rr
      -- 
    rr_1161_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1161_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(168), ack => slice_254_inst_req_0); -- 
    maxPool4_cp_element_group_168: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_168"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(43) & maxPool4_CP_346_elements(170);
      gj_maxPool4_cp_element_group_168 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(168), clk => clk, reset => reset); --
    end block;
    -- CP-element group 169:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: marked-predecessors 
    -- CP-element group 169: 	171 
    -- CP-element group 169: 	378 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	171 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 assign_stmt_97_to_assign_stmt_1138/slice_254_Update/$entry
      -- CP-element group 169: 	 assign_stmt_97_to_assign_stmt_1138/slice_254_update_start_
      -- CP-element group 169: 	 assign_stmt_97_to_assign_stmt_1138/slice_254_Update/cr
      -- 
    cr_1166_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1166_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(169), ack => slice_254_inst_req_1); -- 
    maxPool4_cp_element_group_169: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_169"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(171) & maxPool4_CP_346_elements(378);
      gj_maxPool4_cp_element_group_169 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(169), clk => clk, reset => reset); --
    end block;
    -- CP-element group 170:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	168 
    -- CP-element group 170: successors 
    -- CP-element group 170: marked-successors 
    -- CP-element group 170: 	41 
    -- CP-element group 170: 	168 
    -- CP-element group 170:  members (3) 
      -- CP-element group 170: 	 assign_stmt_97_to_assign_stmt_1138/slice_254_Sample/ra
      -- CP-element group 170: 	 assign_stmt_97_to_assign_stmt_1138/slice_254_sample_completed_
      -- CP-element group 170: 	 assign_stmt_97_to_assign_stmt_1138/slice_254_Sample/$exit
      -- 
    ra_1162_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_254_inst_ack_0, ack => maxPool4_CP_346_elements(170)); -- 
    -- CP-element group 171:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	169 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	376 
    -- CP-element group 171: marked-successors 
    -- CP-element group 171: 	169 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 assign_stmt_97_to_assign_stmt_1138/slice_254_Update/$exit
      -- CP-element group 171: 	 assign_stmt_97_to_assign_stmt_1138/slice_254_Update/ca
      -- CP-element group 171: 	 assign_stmt_97_to_assign_stmt_1138/slice_254_update_completed_
      -- 
    ca_1167_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_254_inst_ack_1, ack => maxPool4_CP_346_elements(171)); -- 
    -- CP-element group 172:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	43 
    -- CP-element group 172: marked-predecessors 
    -- CP-element group 172: 	174 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	174 
    -- CP-element group 172:  members (3) 
      -- CP-element group 172: 	 assign_stmt_97_to_assign_stmt_1138/slice_258_Sample/$entry
      -- CP-element group 172: 	 assign_stmt_97_to_assign_stmt_1138/slice_258_sample_start_
      -- CP-element group 172: 	 assign_stmt_97_to_assign_stmt_1138/slice_258_Sample/rr
      -- 
    rr_1175_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1175_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(172), ack => slice_258_inst_req_0); -- 
    maxPool4_cp_element_group_172: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_172"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(43) & maxPool4_CP_346_elements(174);
      gj_maxPool4_cp_element_group_172 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(172), clk => clk, reset => reset); --
    end block;
    -- CP-element group 173:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: marked-predecessors 
    -- CP-element group 173: 	175 
    -- CP-element group 173: 	378 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	175 
    -- CP-element group 173:  members (3) 
      -- CP-element group 173: 	 assign_stmt_97_to_assign_stmt_1138/slice_258_Update/$entry
      -- CP-element group 173: 	 assign_stmt_97_to_assign_stmt_1138/slice_258_Update/cr
      -- CP-element group 173: 	 assign_stmt_97_to_assign_stmt_1138/slice_258_update_start_
      -- 
    cr_1180_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1180_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(173), ack => slice_258_inst_req_1); -- 
    maxPool4_cp_element_group_173: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_173"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(175) & maxPool4_CP_346_elements(378);
      gj_maxPool4_cp_element_group_173 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(173), clk => clk, reset => reset); --
    end block;
    -- CP-element group 174:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	172 
    -- CP-element group 174: successors 
    -- CP-element group 174: marked-successors 
    -- CP-element group 174: 	41 
    -- CP-element group 174: 	172 
    -- CP-element group 174:  members (3) 
      -- CP-element group 174: 	 assign_stmt_97_to_assign_stmt_1138/slice_258_Sample/$exit
      -- CP-element group 174: 	 assign_stmt_97_to_assign_stmt_1138/slice_258_Sample/ra
      -- CP-element group 174: 	 assign_stmt_97_to_assign_stmt_1138/slice_258_sample_completed_
      -- 
    ra_1176_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_258_inst_ack_0, ack => maxPool4_CP_346_elements(174)); -- 
    -- CP-element group 175:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	173 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	376 
    -- CP-element group 175: marked-successors 
    -- CP-element group 175: 	173 
    -- CP-element group 175:  members (3) 
      -- CP-element group 175: 	 assign_stmt_97_to_assign_stmt_1138/slice_258_Update/$exit
      -- CP-element group 175: 	 assign_stmt_97_to_assign_stmt_1138/slice_258_Update/ca
      -- CP-element group 175: 	 assign_stmt_97_to_assign_stmt_1138/slice_258_update_completed_
      -- 
    ca_1181_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_258_inst_ack_1, ack => maxPool4_CP_346_elements(175)); -- 
    -- CP-element group 176:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	43 
    -- CP-element group 176: marked-predecessors 
    -- CP-element group 176: 	178 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	178 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 assign_stmt_97_to_assign_stmt_1138/slice_262_Sample/$entry
      -- CP-element group 176: 	 assign_stmt_97_to_assign_stmt_1138/slice_262_sample_start_
      -- CP-element group 176: 	 assign_stmt_97_to_assign_stmt_1138/slice_262_Sample/rr
      -- 
    rr_1189_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1189_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(176), ack => slice_262_inst_req_0); -- 
    maxPool4_cp_element_group_176: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_176"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(43) & maxPool4_CP_346_elements(178);
      gj_maxPool4_cp_element_group_176 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(176), clk => clk, reset => reset); --
    end block;
    -- CP-element group 177:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: marked-predecessors 
    -- CP-element group 177: 	179 
    -- CP-element group 177: 	378 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	179 
    -- CP-element group 177:  members (3) 
      -- CP-element group 177: 	 assign_stmt_97_to_assign_stmt_1138/slice_262_update_start_
      -- CP-element group 177: 	 assign_stmt_97_to_assign_stmt_1138/slice_262_Update/cr
      -- CP-element group 177: 	 assign_stmt_97_to_assign_stmt_1138/slice_262_Update/$entry
      -- 
    cr_1194_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1194_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(177), ack => slice_262_inst_req_1); -- 
    maxPool4_cp_element_group_177: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_177"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(179) & maxPool4_CP_346_elements(378);
      gj_maxPool4_cp_element_group_177 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(177), clk => clk, reset => reset); --
    end block;
    -- CP-element group 178:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	176 
    -- CP-element group 178: successors 
    -- CP-element group 178: marked-successors 
    -- CP-element group 178: 	41 
    -- CP-element group 178: 	176 
    -- CP-element group 178:  members (3) 
      -- CP-element group 178: 	 assign_stmt_97_to_assign_stmt_1138/slice_262_Sample/$exit
      -- CP-element group 178: 	 assign_stmt_97_to_assign_stmt_1138/slice_262_sample_completed_
      -- CP-element group 178: 	 assign_stmt_97_to_assign_stmt_1138/slice_262_Sample/ra
      -- 
    ra_1190_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_262_inst_ack_0, ack => maxPool4_CP_346_elements(178)); -- 
    -- CP-element group 179:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	177 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	376 
    -- CP-element group 179: marked-successors 
    -- CP-element group 179: 	177 
    -- CP-element group 179:  members (3) 
      -- CP-element group 179: 	 assign_stmt_97_to_assign_stmt_1138/slice_262_Update/ca
      -- CP-element group 179: 	 assign_stmt_97_to_assign_stmt_1138/slice_262_update_completed_
      -- CP-element group 179: 	 assign_stmt_97_to_assign_stmt_1138/slice_262_Update/$exit
      -- 
    ca_1195_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_262_inst_ack_1, ack => maxPool4_CP_346_elements(179)); -- 
    -- CP-element group 180:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	47 
    -- CP-element group 180: marked-predecessors 
    -- CP-element group 180: 	182 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	182 
    -- CP-element group 180:  members (3) 
      -- CP-element group 180: 	 assign_stmt_97_to_assign_stmt_1138/slice_266_Sample/$entry
      -- CP-element group 180: 	 assign_stmt_97_to_assign_stmt_1138/slice_266_Sample/rr
      -- CP-element group 180: 	 assign_stmt_97_to_assign_stmt_1138/slice_266_sample_start_
      -- 
    rr_1203_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1203_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(180), ack => slice_266_inst_req_0); -- 
    maxPool4_cp_element_group_180: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_180"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(47) & maxPool4_CP_346_elements(182);
      gj_maxPool4_cp_element_group_180 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(180), clk => clk, reset => reset); --
    end block;
    -- CP-element group 181:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: marked-predecessors 
    -- CP-element group 181: 	183 
    -- CP-element group 181: 	321 
    -- CP-element group 181: 	386 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	183 
    -- CP-element group 181:  members (3) 
      -- CP-element group 181: 	 assign_stmt_97_to_assign_stmt_1138/slice_266_Update/cr
      -- CP-element group 181: 	 assign_stmt_97_to_assign_stmt_1138/slice_266_update_start_
      -- CP-element group 181: 	 assign_stmt_97_to_assign_stmt_1138/slice_266_Update/$entry
      -- 
    cr_1208_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1208_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(181), ack => slice_266_inst_req_1); -- 
    maxPool4_cp_element_group_181: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_181"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(183) & maxPool4_CP_346_elements(321) & maxPool4_CP_346_elements(386);
      gj_maxPool4_cp_element_group_181 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(181), clk => clk, reset => reset); --
    end block;
    -- CP-element group 182:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	180 
    -- CP-element group 182: successors 
    -- CP-element group 182: marked-successors 
    -- CP-element group 182: 	45 
    -- CP-element group 182: 	180 
    -- CP-element group 182:  members (3) 
      -- CP-element group 182: 	 assign_stmt_97_to_assign_stmt_1138/slice_266_Sample/ra
      -- CP-element group 182: 	 assign_stmt_97_to_assign_stmt_1138/slice_266_sample_completed_
      -- CP-element group 182: 	 assign_stmt_97_to_assign_stmt_1138/slice_266_Sample/$exit
      -- 
    ra_1204_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_266_inst_ack_0, ack => maxPool4_CP_346_elements(182)); -- 
    -- CP-element group 183:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	181 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	319 
    -- CP-element group 183: 	384 
    -- CP-element group 183: marked-successors 
    -- CP-element group 183: 	181 
    -- CP-element group 183:  members (3) 
      -- CP-element group 183: 	 assign_stmt_97_to_assign_stmt_1138/slice_266_update_completed_
      -- CP-element group 183: 	 assign_stmt_97_to_assign_stmt_1138/slice_266_Update/ca
      -- CP-element group 183: 	 assign_stmt_97_to_assign_stmt_1138/slice_266_Update/$exit
      -- 
    ca_1209_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_266_inst_ack_1, ack => maxPool4_CP_346_elements(183)); -- 
    -- CP-element group 184:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	47 
    -- CP-element group 184: marked-predecessors 
    -- CP-element group 184: 	186 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	186 
    -- CP-element group 184:  members (3) 
      -- CP-element group 184: 	 assign_stmt_97_to_assign_stmt_1138/slice_270_sample_start_
      -- CP-element group 184: 	 assign_stmt_97_to_assign_stmt_1138/slice_270_Sample/$entry
      -- CP-element group 184: 	 assign_stmt_97_to_assign_stmt_1138/slice_270_Sample/rr
      -- 
    rr_1217_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1217_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(184), ack => slice_270_inst_req_0); -- 
    maxPool4_cp_element_group_184: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_184"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(47) & maxPool4_CP_346_elements(186);
      gj_maxPool4_cp_element_group_184 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(184), clk => clk, reset => reset); --
    end block;
    -- CP-element group 185:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: marked-predecessors 
    -- CP-element group 185: 	187 
    -- CP-element group 185: 	321 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	187 
    -- CP-element group 185:  members (3) 
      -- CP-element group 185: 	 assign_stmt_97_to_assign_stmt_1138/slice_270_Update/$entry
      -- CP-element group 185: 	 assign_stmt_97_to_assign_stmt_1138/slice_270_Update/cr
      -- CP-element group 185: 	 assign_stmt_97_to_assign_stmt_1138/slice_270_update_start_
      -- 
    cr_1222_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1222_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(185), ack => slice_270_inst_req_1); -- 
    maxPool4_cp_element_group_185: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_185"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(187) & maxPool4_CP_346_elements(321);
      gj_maxPool4_cp_element_group_185 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(185), clk => clk, reset => reset); --
    end block;
    -- CP-element group 186:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	184 
    -- CP-element group 186: successors 
    -- CP-element group 186: marked-successors 
    -- CP-element group 186: 	45 
    -- CP-element group 186: 	184 
    -- CP-element group 186:  members (3) 
      -- CP-element group 186: 	 assign_stmt_97_to_assign_stmt_1138/slice_270_sample_completed_
      -- CP-element group 186: 	 assign_stmt_97_to_assign_stmt_1138/slice_270_Sample/$exit
      -- CP-element group 186: 	 assign_stmt_97_to_assign_stmt_1138/slice_270_Sample/ra
      -- 
    ra_1218_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_270_inst_ack_0, ack => maxPool4_CP_346_elements(186)); -- 
    -- CP-element group 187:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	185 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	319 
    -- CP-element group 187: marked-successors 
    -- CP-element group 187: 	185 
    -- CP-element group 187:  members (3) 
      -- CP-element group 187: 	 assign_stmt_97_to_assign_stmt_1138/slice_270_Update/ca
      -- CP-element group 187: 	 assign_stmt_97_to_assign_stmt_1138/slice_270_update_completed_
      -- CP-element group 187: 	 assign_stmt_97_to_assign_stmt_1138/slice_270_Update/$exit
      -- 
    ca_1223_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_270_inst_ack_1, ack => maxPool4_CP_346_elements(187)); -- 
    -- CP-element group 188:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	47 
    -- CP-element group 188: marked-predecessors 
    -- CP-element group 188: 	190 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	190 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 assign_stmt_97_to_assign_stmt_1138/slice_274_sample_start_
      -- CP-element group 188: 	 assign_stmt_97_to_assign_stmt_1138/slice_274_Sample/$entry
      -- CP-element group 188: 	 assign_stmt_97_to_assign_stmt_1138/slice_274_Sample/rr
      -- 
    rr_1231_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1231_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(188), ack => slice_274_inst_req_0); -- 
    maxPool4_cp_element_group_188: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_188"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(47) & maxPool4_CP_346_elements(190);
      gj_maxPool4_cp_element_group_188 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(188), clk => clk, reset => reset); --
    end block;
    -- CP-element group 189:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: marked-predecessors 
    -- CP-element group 189: 	191 
    -- CP-element group 189: 	321 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	191 
    -- CP-element group 189:  members (3) 
      -- CP-element group 189: 	 assign_stmt_97_to_assign_stmt_1138/slice_274_update_start_
      -- CP-element group 189: 	 assign_stmt_97_to_assign_stmt_1138/slice_274_Update/$entry
      -- CP-element group 189: 	 assign_stmt_97_to_assign_stmt_1138/slice_274_Update/cr
      -- 
    cr_1236_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1236_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(189), ack => slice_274_inst_req_1); -- 
    maxPool4_cp_element_group_189: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_189"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(191) & maxPool4_CP_346_elements(321);
      gj_maxPool4_cp_element_group_189 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(189), clk => clk, reset => reset); --
    end block;
    -- CP-element group 190:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	188 
    -- CP-element group 190: successors 
    -- CP-element group 190: marked-successors 
    -- CP-element group 190: 	45 
    -- CP-element group 190: 	188 
    -- CP-element group 190:  members (3) 
      -- CP-element group 190: 	 assign_stmt_97_to_assign_stmt_1138/slice_274_sample_completed_
      -- CP-element group 190: 	 assign_stmt_97_to_assign_stmt_1138/slice_274_Sample/$exit
      -- CP-element group 190: 	 assign_stmt_97_to_assign_stmt_1138/slice_274_Sample/ra
      -- 
    ra_1232_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_274_inst_ack_0, ack => maxPool4_CP_346_elements(190)); -- 
    -- CP-element group 191:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	189 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	319 
    -- CP-element group 191: marked-successors 
    -- CP-element group 191: 	189 
    -- CP-element group 191:  members (3) 
      -- CP-element group 191: 	 assign_stmt_97_to_assign_stmt_1138/slice_274_update_completed_
      -- CP-element group 191: 	 assign_stmt_97_to_assign_stmt_1138/slice_274_Update/$exit
      -- CP-element group 191: 	 assign_stmt_97_to_assign_stmt_1138/slice_274_Update/ca
      -- 
    ca_1237_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_274_inst_ack_1, ack => maxPool4_CP_346_elements(191)); -- 
    -- CP-element group 192:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	47 
    -- CP-element group 192: marked-predecessors 
    -- CP-element group 192: 	194 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	194 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 assign_stmt_97_to_assign_stmt_1138/slice_278_sample_start_
      -- CP-element group 192: 	 assign_stmt_97_to_assign_stmt_1138/slice_278_Sample/$entry
      -- CP-element group 192: 	 assign_stmt_97_to_assign_stmt_1138/slice_278_Sample/rr
      -- 
    rr_1245_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1245_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(192), ack => slice_278_inst_req_0); -- 
    maxPool4_cp_element_group_192: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_192"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(47) & maxPool4_CP_346_elements(194);
      gj_maxPool4_cp_element_group_192 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(192), clk => clk, reset => reset); --
    end block;
    -- CP-element group 193:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: marked-predecessors 
    -- CP-element group 193: 	195 
    -- CP-element group 193: 	321 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	195 
    -- CP-element group 193:  members (3) 
      -- CP-element group 193: 	 assign_stmt_97_to_assign_stmt_1138/slice_278_update_start_
      -- CP-element group 193: 	 assign_stmt_97_to_assign_stmt_1138/slice_278_Update/$entry
      -- CP-element group 193: 	 assign_stmt_97_to_assign_stmt_1138/slice_278_Update/cr
      -- 
    cr_1250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(193), ack => slice_278_inst_req_1); -- 
    maxPool4_cp_element_group_193: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_193"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(195) & maxPool4_CP_346_elements(321);
      gj_maxPool4_cp_element_group_193 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(193), clk => clk, reset => reset); --
    end block;
    -- CP-element group 194:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	192 
    -- CP-element group 194: successors 
    -- CP-element group 194: marked-successors 
    -- CP-element group 194: 	45 
    -- CP-element group 194: 	192 
    -- CP-element group 194:  members (3) 
      -- CP-element group 194: 	 assign_stmt_97_to_assign_stmt_1138/slice_278_sample_completed_
      -- CP-element group 194: 	 assign_stmt_97_to_assign_stmt_1138/slice_278_Sample/$exit
      -- CP-element group 194: 	 assign_stmt_97_to_assign_stmt_1138/slice_278_Sample/ra
      -- 
    ra_1246_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_278_inst_ack_0, ack => maxPool4_CP_346_elements(194)); -- 
    -- CP-element group 195:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	193 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	319 
    -- CP-element group 195: marked-successors 
    -- CP-element group 195: 	193 
    -- CP-element group 195:  members (3) 
      -- CP-element group 195: 	 assign_stmt_97_to_assign_stmt_1138/slice_278_update_completed_
      -- CP-element group 195: 	 assign_stmt_97_to_assign_stmt_1138/slice_278_Update/$exit
      -- CP-element group 195: 	 assign_stmt_97_to_assign_stmt_1138/slice_278_Update/ca
      -- 
    ca_1251_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_278_inst_ack_1, ack => maxPool4_CP_346_elements(195)); -- 
    -- CP-element group 196:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	47 
    -- CP-element group 196: marked-predecessors 
    -- CP-element group 196: 	198 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	198 
    -- CP-element group 196:  members (3) 
      -- CP-element group 196: 	 assign_stmt_97_to_assign_stmt_1138/slice_282_sample_start_
      -- CP-element group 196: 	 assign_stmt_97_to_assign_stmt_1138/slice_282_Sample/$entry
      -- CP-element group 196: 	 assign_stmt_97_to_assign_stmt_1138/slice_282_Sample/rr
      -- 
    rr_1259_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1259_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(196), ack => slice_282_inst_req_0); -- 
    maxPool4_cp_element_group_196: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_196"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(47) & maxPool4_CP_346_elements(198);
      gj_maxPool4_cp_element_group_196 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(196), clk => clk, reset => reset); --
    end block;
    -- CP-element group 197:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: marked-predecessors 
    -- CP-element group 197: 	199 
    -- CP-element group 197: 	340 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	199 
    -- CP-element group 197:  members (3) 
      -- CP-element group 197: 	 assign_stmt_97_to_assign_stmt_1138/slice_282_update_start_
      -- CP-element group 197: 	 assign_stmt_97_to_assign_stmt_1138/slice_282_Update/$entry
      -- CP-element group 197: 	 assign_stmt_97_to_assign_stmt_1138/slice_282_Update/cr
      -- 
    cr_1264_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1264_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(197), ack => slice_282_inst_req_1); -- 
    maxPool4_cp_element_group_197: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_197"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(199) & maxPool4_CP_346_elements(340);
      gj_maxPool4_cp_element_group_197 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(197), clk => clk, reset => reset); --
    end block;
    -- CP-element group 198:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	196 
    -- CP-element group 198: successors 
    -- CP-element group 198: marked-successors 
    -- CP-element group 198: 	45 
    -- CP-element group 198: 	196 
    -- CP-element group 198:  members (3) 
      -- CP-element group 198: 	 assign_stmt_97_to_assign_stmt_1138/slice_282_sample_completed_
      -- CP-element group 198: 	 assign_stmt_97_to_assign_stmt_1138/slice_282_Sample/$exit
      -- CP-element group 198: 	 assign_stmt_97_to_assign_stmt_1138/slice_282_Sample/ra
      -- 
    ra_1260_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_282_inst_ack_0, ack => maxPool4_CP_346_elements(198)); -- 
    -- CP-element group 199:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	197 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	338 
    -- CP-element group 199: marked-successors 
    -- CP-element group 199: 	197 
    -- CP-element group 199:  members (3) 
      -- CP-element group 199: 	 assign_stmt_97_to_assign_stmt_1138/slice_282_update_completed_
      -- CP-element group 199: 	 assign_stmt_97_to_assign_stmt_1138/slice_282_Update/$exit
      -- CP-element group 199: 	 assign_stmt_97_to_assign_stmt_1138/slice_282_Update/ca
      -- 
    ca_1265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_282_inst_ack_1, ack => maxPool4_CP_346_elements(199)); -- 
    -- CP-element group 200:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	47 
    -- CP-element group 200: marked-predecessors 
    -- CP-element group 200: 	202 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	202 
    -- CP-element group 200:  members (3) 
      -- CP-element group 200: 	 assign_stmt_97_to_assign_stmt_1138/slice_286_sample_start_
      -- CP-element group 200: 	 assign_stmt_97_to_assign_stmt_1138/slice_286_Sample/$entry
      -- CP-element group 200: 	 assign_stmt_97_to_assign_stmt_1138/slice_286_Sample/rr
      -- 
    rr_1273_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1273_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(200), ack => slice_286_inst_req_0); -- 
    maxPool4_cp_element_group_200: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_200"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(47) & maxPool4_CP_346_elements(202);
      gj_maxPool4_cp_element_group_200 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(200), clk => clk, reset => reset); --
    end block;
    -- CP-element group 201:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: marked-predecessors 
    -- CP-element group 201: 	203 
    -- CP-element group 201: 	340 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	203 
    -- CP-element group 201:  members (3) 
      -- CP-element group 201: 	 assign_stmt_97_to_assign_stmt_1138/slice_286_update_start_
      -- CP-element group 201: 	 assign_stmt_97_to_assign_stmt_1138/slice_286_Update/$entry
      -- CP-element group 201: 	 assign_stmt_97_to_assign_stmt_1138/slice_286_Update/cr
      -- 
    cr_1278_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1278_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(201), ack => slice_286_inst_req_1); -- 
    maxPool4_cp_element_group_201: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_201"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(203) & maxPool4_CP_346_elements(340);
      gj_maxPool4_cp_element_group_201 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(201), clk => clk, reset => reset); --
    end block;
    -- CP-element group 202:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	200 
    -- CP-element group 202: successors 
    -- CP-element group 202: marked-successors 
    -- CP-element group 202: 	45 
    -- CP-element group 202: 	200 
    -- CP-element group 202:  members (3) 
      -- CP-element group 202: 	 assign_stmt_97_to_assign_stmt_1138/slice_286_sample_completed_
      -- CP-element group 202: 	 assign_stmt_97_to_assign_stmt_1138/slice_286_Sample/$exit
      -- CP-element group 202: 	 assign_stmt_97_to_assign_stmt_1138/slice_286_Sample/ra
      -- 
    ra_1274_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_286_inst_ack_0, ack => maxPool4_CP_346_elements(202)); -- 
    -- CP-element group 203:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	201 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	338 
    -- CP-element group 203: marked-successors 
    -- CP-element group 203: 	201 
    -- CP-element group 203:  members (3) 
      -- CP-element group 203: 	 assign_stmt_97_to_assign_stmt_1138/slice_286_update_completed_
      -- CP-element group 203: 	 assign_stmt_97_to_assign_stmt_1138/slice_286_Update/$exit
      -- CP-element group 203: 	 assign_stmt_97_to_assign_stmt_1138/slice_286_Update/ca
      -- 
    ca_1279_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 203_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_286_inst_ack_1, ack => maxPool4_CP_346_elements(203)); -- 
    -- CP-element group 204:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	47 
    -- CP-element group 204: marked-predecessors 
    -- CP-element group 204: 	206 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	206 
    -- CP-element group 204:  members (3) 
      -- CP-element group 204: 	 assign_stmt_97_to_assign_stmt_1138/slice_290_sample_start_
      -- CP-element group 204: 	 assign_stmt_97_to_assign_stmt_1138/slice_290_Sample/$entry
      -- CP-element group 204: 	 assign_stmt_97_to_assign_stmt_1138/slice_290_Sample/rr
      -- 
    rr_1287_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1287_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(204), ack => slice_290_inst_req_0); -- 
    maxPool4_cp_element_group_204: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_204"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(47) & maxPool4_CP_346_elements(206);
      gj_maxPool4_cp_element_group_204 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(204), clk => clk, reset => reset); --
    end block;
    -- CP-element group 205:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: marked-predecessors 
    -- CP-element group 205: 	207 
    -- CP-element group 205: 	340 
    -- CP-element group 205: successors 
    -- CP-element group 205: 	207 
    -- CP-element group 205:  members (3) 
      -- CP-element group 205: 	 assign_stmt_97_to_assign_stmt_1138/slice_290_update_start_
      -- CP-element group 205: 	 assign_stmt_97_to_assign_stmt_1138/slice_290_Update/$entry
      -- CP-element group 205: 	 assign_stmt_97_to_assign_stmt_1138/slice_290_Update/cr
      -- 
    cr_1292_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1292_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(205), ack => slice_290_inst_req_1); -- 
    maxPool4_cp_element_group_205: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_205"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(207) & maxPool4_CP_346_elements(340);
      gj_maxPool4_cp_element_group_205 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(205), clk => clk, reset => reset); --
    end block;
    -- CP-element group 206:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	204 
    -- CP-element group 206: successors 
    -- CP-element group 206: marked-successors 
    -- CP-element group 206: 	45 
    -- CP-element group 206: 	204 
    -- CP-element group 206:  members (3) 
      -- CP-element group 206: 	 assign_stmt_97_to_assign_stmt_1138/slice_290_sample_completed_
      -- CP-element group 206: 	 assign_stmt_97_to_assign_stmt_1138/slice_290_Sample/$exit
      -- CP-element group 206: 	 assign_stmt_97_to_assign_stmt_1138/slice_290_Sample/ra
      -- 
    ra_1288_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 206_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_290_inst_ack_0, ack => maxPool4_CP_346_elements(206)); -- 
    -- CP-element group 207:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	205 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	338 
    -- CP-element group 207: marked-successors 
    -- CP-element group 207: 	205 
    -- CP-element group 207:  members (3) 
      -- CP-element group 207: 	 assign_stmt_97_to_assign_stmt_1138/slice_290_update_completed_
      -- CP-element group 207: 	 assign_stmt_97_to_assign_stmt_1138/slice_290_Update/$exit
      -- CP-element group 207: 	 assign_stmt_97_to_assign_stmt_1138/slice_290_Update/ca
      -- 
    ca_1293_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 207_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_290_inst_ack_1, ack => maxPool4_CP_346_elements(207)); -- 
    -- CP-element group 208:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	47 
    -- CP-element group 208: marked-predecessors 
    -- CP-element group 208: 	210 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	210 
    -- CP-element group 208:  members (3) 
      -- CP-element group 208: 	 assign_stmt_97_to_assign_stmt_1138/slice_294_sample_start_
      -- CP-element group 208: 	 assign_stmt_97_to_assign_stmt_1138/slice_294_Sample/$entry
      -- CP-element group 208: 	 assign_stmt_97_to_assign_stmt_1138/slice_294_Sample/rr
      -- 
    rr_1301_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1301_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(208), ack => slice_294_inst_req_0); -- 
    maxPool4_cp_element_group_208: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_208"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(47) & maxPool4_CP_346_elements(210);
      gj_maxPool4_cp_element_group_208 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(208), clk => clk, reset => reset); --
    end block;
    -- CP-element group 209:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: marked-predecessors 
    -- CP-element group 209: 	211 
    -- CP-element group 209: 	340 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	211 
    -- CP-element group 209:  members (3) 
      -- CP-element group 209: 	 assign_stmt_97_to_assign_stmt_1138/slice_294_update_start_
      -- CP-element group 209: 	 assign_stmt_97_to_assign_stmt_1138/slice_294_Update/$entry
      -- CP-element group 209: 	 assign_stmt_97_to_assign_stmt_1138/slice_294_Update/cr
      -- 
    cr_1306_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1306_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(209), ack => slice_294_inst_req_1); -- 
    maxPool4_cp_element_group_209: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_209"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(211) & maxPool4_CP_346_elements(340);
      gj_maxPool4_cp_element_group_209 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(209), clk => clk, reset => reset); --
    end block;
    -- CP-element group 210:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	208 
    -- CP-element group 210: successors 
    -- CP-element group 210: marked-successors 
    -- CP-element group 210: 	45 
    -- CP-element group 210: 	208 
    -- CP-element group 210:  members (3) 
      -- CP-element group 210: 	 assign_stmt_97_to_assign_stmt_1138/slice_294_sample_completed_
      -- CP-element group 210: 	 assign_stmt_97_to_assign_stmt_1138/slice_294_Sample/$exit
      -- CP-element group 210: 	 assign_stmt_97_to_assign_stmt_1138/slice_294_Sample/ra
      -- 
    ra_1302_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 210_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_294_inst_ack_0, ack => maxPool4_CP_346_elements(210)); -- 
    -- CP-element group 211:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	209 
    -- CP-element group 211: successors 
    -- CP-element group 211: 	338 
    -- CP-element group 211: marked-successors 
    -- CP-element group 211: 	209 
    -- CP-element group 211:  members (3) 
      -- CP-element group 211: 	 assign_stmt_97_to_assign_stmt_1138/slice_294_update_completed_
      -- CP-element group 211: 	 assign_stmt_97_to_assign_stmt_1138/slice_294_Update/$exit
      -- CP-element group 211: 	 assign_stmt_97_to_assign_stmt_1138/slice_294_Update/ca
      -- 
    ca_1307_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 211_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_294_inst_ack_1, ack => maxPool4_CP_346_elements(211)); -- 
    -- CP-element group 212:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	47 
    -- CP-element group 212: marked-predecessors 
    -- CP-element group 212: 	214 
    -- CP-element group 212: successors 
    -- CP-element group 212: 	214 
    -- CP-element group 212:  members (3) 
      -- CP-element group 212: 	 assign_stmt_97_to_assign_stmt_1138/slice_298_sample_start_
      -- CP-element group 212: 	 assign_stmt_97_to_assign_stmt_1138/slice_298_Sample/$entry
      -- CP-element group 212: 	 assign_stmt_97_to_assign_stmt_1138/slice_298_Sample/rr
      -- 
    rr_1315_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1315_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(212), ack => slice_298_inst_req_0); -- 
    maxPool4_cp_element_group_212: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_212"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(47) & maxPool4_CP_346_elements(214);
      gj_maxPool4_cp_element_group_212 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(212), clk => clk, reset => reset); --
    end block;
    -- CP-element group 213:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: marked-predecessors 
    -- CP-element group 213: 	215 
    -- CP-element group 213: 	359 
    -- CP-element group 213: successors 
    -- CP-element group 213: 	215 
    -- CP-element group 213:  members (3) 
      -- CP-element group 213: 	 assign_stmt_97_to_assign_stmt_1138/slice_298_update_start_
      -- CP-element group 213: 	 assign_stmt_97_to_assign_stmt_1138/slice_298_Update/$entry
      -- CP-element group 213: 	 assign_stmt_97_to_assign_stmt_1138/slice_298_Update/cr
      -- 
    cr_1320_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1320_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(213), ack => slice_298_inst_req_1); -- 
    maxPool4_cp_element_group_213: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_213"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(215) & maxPool4_CP_346_elements(359);
      gj_maxPool4_cp_element_group_213 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(213), clk => clk, reset => reset); --
    end block;
    -- CP-element group 214:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	212 
    -- CP-element group 214: successors 
    -- CP-element group 214: marked-successors 
    -- CP-element group 214: 	45 
    -- CP-element group 214: 	212 
    -- CP-element group 214:  members (3) 
      -- CP-element group 214: 	 assign_stmt_97_to_assign_stmt_1138/slice_298_sample_completed_
      -- CP-element group 214: 	 assign_stmt_97_to_assign_stmt_1138/slice_298_Sample/$exit
      -- CP-element group 214: 	 assign_stmt_97_to_assign_stmt_1138/slice_298_Sample/ra
      -- 
    ra_1316_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 214_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_298_inst_ack_0, ack => maxPool4_CP_346_elements(214)); -- 
    -- CP-element group 215:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	213 
    -- CP-element group 215: successors 
    -- CP-element group 215: 	357 
    -- CP-element group 215: marked-successors 
    -- CP-element group 215: 	213 
    -- CP-element group 215:  members (3) 
      -- CP-element group 215: 	 assign_stmt_97_to_assign_stmt_1138/slice_298_update_completed_
      -- CP-element group 215: 	 assign_stmt_97_to_assign_stmt_1138/slice_298_Update/$exit
      -- CP-element group 215: 	 assign_stmt_97_to_assign_stmt_1138/slice_298_Update/ca
      -- 
    ca_1321_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 215_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_298_inst_ack_1, ack => maxPool4_CP_346_elements(215)); -- 
    -- CP-element group 216:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	47 
    -- CP-element group 216: marked-predecessors 
    -- CP-element group 216: 	218 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	218 
    -- CP-element group 216:  members (3) 
      -- CP-element group 216: 	 assign_stmt_97_to_assign_stmt_1138/slice_302_sample_start_
      -- CP-element group 216: 	 assign_stmt_97_to_assign_stmt_1138/slice_302_Sample/$entry
      -- CP-element group 216: 	 assign_stmt_97_to_assign_stmt_1138/slice_302_Sample/rr
      -- 
    rr_1329_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1329_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(216), ack => slice_302_inst_req_0); -- 
    maxPool4_cp_element_group_216: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_216"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(47) & maxPool4_CP_346_elements(218);
      gj_maxPool4_cp_element_group_216 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(216), clk => clk, reset => reset); --
    end block;
    -- CP-element group 217:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: marked-predecessors 
    -- CP-element group 217: 	219 
    -- CP-element group 217: 	359 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	219 
    -- CP-element group 217:  members (3) 
      -- CP-element group 217: 	 assign_stmt_97_to_assign_stmt_1138/slice_302_update_start_
      -- CP-element group 217: 	 assign_stmt_97_to_assign_stmt_1138/slice_302_Update/$entry
      -- CP-element group 217: 	 assign_stmt_97_to_assign_stmt_1138/slice_302_Update/cr
      -- 
    cr_1334_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1334_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(217), ack => slice_302_inst_req_1); -- 
    maxPool4_cp_element_group_217: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_217"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(219) & maxPool4_CP_346_elements(359);
      gj_maxPool4_cp_element_group_217 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(217), clk => clk, reset => reset); --
    end block;
    -- CP-element group 218:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	216 
    -- CP-element group 218: successors 
    -- CP-element group 218: marked-successors 
    -- CP-element group 218: 	45 
    -- CP-element group 218: 	216 
    -- CP-element group 218:  members (3) 
      -- CP-element group 218: 	 assign_stmt_97_to_assign_stmt_1138/slice_302_sample_completed_
      -- CP-element group 218: 	 assign_stmt_97_to_assign_stmt_1138/slice_302_Sample/$exit
      -- CP-element group 218: 	 assign_stmt_97_to_assign_stmt_1138/slice_302_Sample/ra
      -- 
    ra_1330_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 218_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_302_inst_ack_0, ack => maxPool4_CP_346_elements(218)); -- 
    -- CP-element group 219:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	217 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	357 
    -- CP-element group 219: marked-successors 
    -- CP-element group 219: 	217 
    -- CP-element group 219:  members (3) 
      -- CP-element group 219: 	 assign_stmt_97_to_assign_stmt_1138/slice_302_update_completed_
      -- CP-element group 219: 	 assign_stmt_97_to_assign_stmt_1138/slice_302_Update/$exit
      -- CP-element group 219: 	 assign_stmt_97_to_assign_stmt_1138/slice_302_Update/ca
      -- 
    ca_1335_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 219_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_302_inst_ack_1, ack => maxPool4_CP_346_elements(219)); -- 
    -- CP-element group 220:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	47 
    -- CP-element group 220: marked-predecessors 
    -- CP-element group 220: 	222 
    -- CP-element group 220: successors 
    -- CP-element group 220: 	222 
    -- CP-element group 220:  members (3) 
      -- CP-element group 220: 	 assign_stmt_97_to_assign_stmt_1138/slice_306_sample_start_
      -- CP-element group 220: 	 assign_stmt_97_to_assign_stmt_1138/slice_306_Sample/$entry
      -- CP-element group 220: 	 assign_stmt_97_to_assign_stmt_1138/slice_306_Sample/rr
      -- 
    rr_1343_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1343_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(220), ack => slice_306_inst_req_0); -- 
    maxPool4_cp_element_group_220: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_220"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(47) & maxPool4_CP_346_elements(222);
      gj_maxPool4_cp_element_group_220 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(220), clk => clk, reset => reset); --
    end block;
    -- CP-element group 221:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: marked-predecessors 
    -- CP-element group 221: 	223 
    -- CP-element group 221: 	359 
    -- CP-element group 221: successors 
    -- CP-element group 221: 	223 
    -- CP-element group 221:  members (3) 
      -- CP-element group 221: 	 assign_stmt_97_to_assign_stmt_1138/slice_306_update_start_
      -- CP-element group 221: 	 assign_stmt_97_to_assign_stmt_1138/slice_306_Update/$entry
      -- CP-element group 221: 	 assign_stmt_97_to_assign_stmt_1138/slice_306_Update/cr
      -- 
    cr_1348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(221), ack => slice_306_inst_req_1); -- 
    maxPool4_cp_element_group_221: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_221"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(223) & maxPool4_CP_346_elements(359);
      gj_maxPool4_cp_element_group_221 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(221), clk => clk, reset => reset); --
    end block;
    -- CP-element group 222:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	220 
    -- CP-element group 222: successors 
    -- CP-element group 222: marked-successors 
    -- CP-element group 222: 	45 
    -- CP-element group 222: 	220 
    -- CP-element group 222:  members (3) 
      -- CP-element group 222: 	 assign_stmt_97_to_assign_stmt_1138/slice_306_sample_completed_
      -- CP-element group 222: 	 assign_stmt_97_to_assign_stmt_1138/slice_306_Sample/$exit
      -- CP-element group 222: 	 assign_stmt_97_to_assign_stmt_1138/slice_306_Sample/ra
      -- 
    ra_1344_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 222_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_306_inst_ack_0, ack => maxPool4_CP_346_elements(222)); -- 
    -- CP-element group 223:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	221 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	357 
    -- CP-element group 223: marked-successors 
    -- CP-element group 223: 	221 
    -- CP-element group 223:  members (3) 
      -- CP-element group 223: 	 assign_stmt_97_to_assign_stmt_1138/slice_306_update_completed_
      -- CP-element group 223: 	 assign_stmt_97_to_assign_stmt_1138/slice_306_Update/$exit
      -- CP-element group 223: 	 assign_stmt_97_to_assign_stmt_1138/slice_306_Update/ca
      -- 
    ca_1349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 223_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_306_inst_ack_1, ack => maxPool4_CP_346_elements(223)); -- 
    -- CP-element group 224:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	47 
    -- CP-element group 224: marked-predecessors 
    -- CP-element group 224: 	226 
    -- CP-element group 224: successors 
    -- CP-element group 224: 	226 
    -- CP-element group 224:  members (3) 
      -- CP-element group 224: 	 assign_stmt_97_to_assign_stmt_1138/slice_310_sample_start_
      -- CP-element group 224: 	 assign_stmt_97_to_assign_stmt_1138/slice_310_Sample/$entry
      -- CP-element group 224: 	 assign_stmt_97_to_assign_stmt_1138/slice_310_Sample/rr
      -- 
    rr_1357_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1357_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(224), ack => slice_310_inst_req_0); -- 
    maxPool4_cp_element_group_224: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_224"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(47) & maxPool4_CP_346_elements(226);
      gj_maxPool4_cp_element_group_224 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(224), clk => clk, reset => reset); --
    end block;
    -- CP-element group 225:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: marked-predecessors 
    -- CP-element group 225: 	227 
    -- CP-element group 225: 	359 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	227 
    -- CP-element group 225:  members (3) 
      -- CP-element group 225: 	 assign_stmt_97_to_assign_stmt_1138/slice_310_update_start_
      -- CP-element group 225: 	 assign_stmt_97_to_assign_stmt_1138/slice_310_Update/$entry
      -- CP-element group 225: 	 assign_stmt_97_to_assign_stmt_1138/slice_310_Update/cr
      -- 
    cr_1362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(225), ack => slice_310_inst_req_1); -- 
    maxPool4_cp_element_group_225: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_225"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(227) & maxPool4_CP_346_elements(359);
      gj_maxPool4_cp_element_group_225 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(225), clk => clk, reset => reset); --
    end block;
    -- CP-element group 226:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	224 
    -- CP-element group 226: successors 
    -- CP-element group 226: marked-successors 
    -- CP-element group 226: 	45 
    -- CP-element group 226: 	224 
    -- CP-element group 226:  members (3) 
      -- CP-element group 226: 	 assign_stmt_97_to_assign_stmt_1138/slice_310_sample_completed_
      -- CP-element group 226: 	 assign_stmt_97_to_assign_stmt_1138/slice_310_Sample/$exit
      -- CP-element group 226: 	 assign_stmt_97_to_assign_stmt_1138/slice_310_Sample/ra
      -- 
    ra_1358_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 226_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_310_inst_ack_0, ack => maxPool4_CP_346_elements(226)); -- 
    -- CP-element group 227:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	225 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	357 
    -- CP-element group 227: marked-successors 
    -- CP-element group 227: 	225 
    -- CP-element group 227:  members (3) 
      -- CP-element group 227: 	 assign_stmt_97_to_assign_stmt_1138/slice_310_update_completed_
      -- CP-element group 227: 	 assign_stmt_97_to_assign_stmt_1138/slice_310_Update/$exit
      -- CP-element group 227: 	 assign_stmt_97_to_assign_stmt_1138/slice_310_Update/ca
      -- 
    ca_1363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 227_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_310_inst_ack_1, ack => maxPool4_CP_346_elements(227)); -- 
    -- CP-element group 228:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	47 
    -- CP-element group 228: marked-predecessors 
    -- CP-element group 228: 	230 
    -- CP-element group 228: successors 
    -- CP-element group 228: 	230 
    -- CP-element group 228:  members (3) 
      -- CP-element group 228: 	 assign_stmt_97_to_assign_stmt_1138/slice_314_sample_start_
      -- CP-element group 228: 	 assign_stmt_97_to_assign_stmt_1138/slice_314_Sample/$entry
      -- CP-element group 228: 	 assign_stmt_97_to_assign_stmt_1138/slice_314_Sample/rr
      -- 
    rr_1371_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1371_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(228), ack => slice_314_inst_req_0); -- 
    maxPool4_cp_element_group_228: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_228"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(47) & maxPool4_CP_346_elements(230);
      gj_maxPool4_cp_element_group_228 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(228), clk => clk, reset => reset); --
    end block;
    -- CP-element group 229:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: marked-predecessors 
    -- CP-element group 229: 	231 
    -- CP-element group 229: 	378 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	231 
    -- CP-element group 229:  members (3) 
      -- CP-element group 229: 	 assign_stmt_97_to_assign_stmt_1138/slice_314_update_start_
      -- CP-element group 229: 	 assign_stmt_97_to_assign_stmt_1138/slice_314_Update/$entry
      -- CP-element group 229: 	 assign_stmt_97_to_assign_stmt_1138/slice_314_Update/cr
      -- 
    cr_1376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(229), ack => slice_314_inst_req_1); -- 
    maxPool4_cp_element_group_229: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_229"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(231) & maxPool4_CP_346_elements(378);
      gj_maxPool4_cp_element_group_229 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(229), clk => clk, reset => reset); --
    end block;
    -- CP-element group 230:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	228 
    -- CP-element group 230: successors 
    -- CP-element group 230: marked-successors 
    -- CP-element group 230: 	45 
    -- CP-element group 230: 	228 
    -- CP-element group 230:  members (3) 
      -- CP-element group 230: 	 assign_stmt_97_to_assign_stmt_1138/slice_314_sample_completed_
      -- CP-element group 230: 	 assign_stmt_97_to_assign_stmt_1138/slice_314_Sample/$exit
      -- CP-element group 230: 	 assign_stmt_97_to_assign_stmt_1138/slice_314_Sample/ra
      -- 
    ra_1372_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 230_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_314_inst_ack_0, ack => maxPool4_CP_346_elements(230)); -- 
    -- CP-element group 231:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	229 
    -- CP-element group 231: successors 
    -- CP-element group 231: 	376 
    -- CP-element group 231: marked-successors 
    -- CP-element group 231: 	229 
    -- CP-element group 231:  members (3) 
      -- CP-element group 231: 	 assign_stmt_97_to_assign_stmt_1138/slice_314_update_completed_
      -- CP-element group 231: 	 assign_stmt_97_to_assign_stmt_1138/slice_314_Update/$exit
      -- CP-element group 231: 	 assign_stmt_97_to_assign_stmt_1138/slice_314_Update/ca
      -- 
    ca_1377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 231_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_314_inst_ack_1, ack => maxPool4_CP_346_elements(231)); -- 
    -- CP-element group 232:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	47 
    -- CP-element group 232: marked-predecessors 
    -- CP-element group 232: 	234 
    -- CP-element group 232: successors 
    -- CP-element group 232: 	234 
    -- CP-element group 232:  members (3) 
      -- CP-element group 232: 	 assign_stmt_97_to_assign_stmt_1138/slice_318_sample_start_
      -- CP-element group 232: 	 assign_stmt_97_to_assign_stmt_1138/slice_318_Sample/$entry
      -- CP-element group 232: 	 assign_stmt_97_to_assign_stmt_1138/slice_318_Sample/rr
      -- 
    rr_1385_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1385_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(232), ack => slice_318_inst_req_0); -- 
    maxPool4_cp_element_group_232: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_232"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(47) & maxPool4_CP_346_elements(234);
      gj_maxPool4_cp_element_group_232 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(232), clk => clk, reset => reset); --
    end block;
    -- CP-element group 233:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: marked-predecessors 
    -- CP-element group 233: 	235 
    -- CP-element group 233: 	378 
    -- CP-element group 233: successors 
    -- CP-element group 233: 	235 
    -- CP-element group 233:  members (3) 
      -- CP-element group 233: 	 assign_stmt_97_to_assign_stmt_1138/slice_318_update_start_
      -- CP-element group 233: 	 assign_stmt_97_to_assign_stmt_1138/slice_318_Update/$entry
      -- CP-element group 233: 	 assign_stmt_97_to_assign_stmt_1138/slice_318_Update/cr
      -- 
    cr_1390_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1390_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(233), ack => slice_318_inst_req_1); -- 
    maxPool4_cp_element_group_233: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_233"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(235) & maxPool4_CP_346_elements(378);
      gj_maxPool4_cp_element_group_233 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(233), clk => clk, reset => reset); --
    end block;
    -- CP-element group 234:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	232 
    -- CP-element group 234: successors 
    -- CP-element group 234: marked-successors 
    -- CP-element group 234: 	45 
    -- CP-element group 234: 	232 
    -- CP-element group 234:  members (3) 
      -- CP-element group 234: 	 assign_stmt_97_to_assign_stmt_1138/slice_318_sample_completed_
      -- CP-element group 234: 	 assign_stmt_97_to_assign_stmt_1138/slice_318_Sample/$exit
      -- CP-element group 234: 	 assign_stmt_97_to_assign_stmt_1138/slice_318_Sample/ra
      -- 
    ra_1386_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 234_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_318_inst_ack_0, ack => maxPool4_CP_346_elements(234)); -- 
    -- CP-element group 235:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	233 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	376 
    -- CP-element group 235: marked-successors 
    -- CP-element group 235: 	233 
    -- CP-element group 235:  members (3) 
      -- CP-element group 235: 	 assign_stmt_97_to_assign_stmt_1138/slice_318_update_completed_
      -- CP-element group 235: 	 assign_stmt_97_to_assign_stmt_1138/slice_318_Update/$exit
      -- CP-element group 235: 	 assign_stmt_97_to_assign_stmt_1138/slice_318_Update/ca
      -- 
    ca_1391_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 235_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_318_inst_ack_1, ack => maxPool4_CP_346_elements(235)); -- 
    -- CP-element group 236:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	47 
    -- CP-element group 236: marked-predecessors 
    -- CP-element group 236: 	238 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	238 
    -- CP-element group 236:  members (3) 
      -- CP-element group 236: 	 assign_stmt_97_to_assign_stmt_1138/slice_322_sample_start_
      -- CP-element group 236: 	 assign_stmt_97_to_assign_stmt_1138/slice_322_Sample/$entry
      -- CP-element group 236: 	 assign_stmt_97_to_assign_stmt_1138/slice_322_Sample/rr
      -- 
    rr_1399_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1399_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(236), ack => slice_322_inst_req_0); -- 
    maxPool4_cp_element_group_236: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_236"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(47) & maxPool4_CP_346_elements(238);
      gj_maxPool4_cp_element_group_236 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(236), clk => clk, reset => reset); --
    end block;
    -- CP-element group 237:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: marked-predecessors 
    -- CP-element group 237: 	239 
    -- CP-element group 237: 	378 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	239 
    -- CP-element group 237:  members (3) 
      -- CP-element group 237: 	 assign_stmt_97_to_assign_stmt_1138/slice_322_update_start_
      -- CP-element group 237: 	 assign_stmt_97_to_assign_stmt_1138/slice_322_Update/$entry
      -- CP-element group 237: 	 assign_stmt_97_to_assign_stmt_1138/slice_322_Update/cr
      -- 
    cr_1404_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1404_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(237), ack => slice_322_inst_req_1); -- 
    maxPool4_cp_element_group_237: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_237"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(239) & maxPool4_CP_346_elements(378);
      gj_maxPool4_cp_element_group_237 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(237), clk => clk, reset => reset); --
    end block;
    -- CP-element group 238:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	236 
    -- CP-element group 238: successors 
    -- CP-element group 238: marked-successors 
    -- CP-element group 238: 	45 
    -- CP-element group 238: 	236 
    -- CP-element group 238:  members (3) 
      -- CP-element group 238: 	 assign_stmt_97_to_assign_stmt_1138/slice_322_sample_completed_
      -- CP-element group 238: 	 assign_stmt_97_to_assign_stmt_1138/slice_322_Sample/$exit
      -- CP-element group 238: 	 assign_stmt_97_to_assign_stmt_1138/slice_322_Sample/ra
      -- 
    ra_1400_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 238_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_322_inst_ack_0, ack => maxPool4_CP_346_elements(238)); -- 
    -- CP-element group 239:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	237 
    -- CP-element group 239: successors 
    -- CP-element group 239: 	376 
    -- CP-element group 239: marked-successors 
    -- CP-element group 239: 	237 
    -- CP-element group 239:  members (3) 
      -- CP-element group 239: 	 assign_stmt_97_to_assign_stmt_1138/slice_322_update_completed_
      -- CP-element group 239: 	 assign_stmt_97_to_assign_stmt_1138/slice_322_Update/$exit
      -- CP-element group 239: 	 assign_stmt_97_to_assign_stmt_1138/slice_322_Update/ca
      -- 
    ca_1405_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 239_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_322_inst_ack_1, ack => maxPool4_CP_346_elements(239)); -- 
    -- CP-element group 240:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	47 
    -- CP-element group 240: marked-predecessors 
    -- CP-element group 240: 	242 
    -- CP-element group 240: successors 
    -- CP-element group 240: 	242 
    -- CP-element group 240:  members (3) 
      -- CP-element group 240: 	 assign_stmt_97_to_assign_stmt_1138/slice_326_sample_start_
      -- CP-element group 240: 	 assign_stmt_97_to_assign_stmt_1138/slice_326_Sample/$entry
      -- CP-element group 240: 	 assign_stmt_97_to_assign_stmt_1138/slice_326_Sample/rr
      -- 
    rr_1413_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1413_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(240), ack => slice_326_inst_req_0); -- 
    maxPool4_cp_element_group_240: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_240"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(47) & maxPool4_CP_346_elements(242);
      gj_maxPool4_cp_element_group_240 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(240), clk => clk, reset => reset); --
    end block;
    -- CP-element group 241:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: marked-predecessors 
    -- CP-element group 241: 	243 
    -- CP-element group 241: 	378 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	243 
    -- CP-element group 241:  members (3) 
      -- CP-element group 241: 	 assign_stmt_97_to_assign_stmt_1138/slice_326_update_start_
      -- CP-element group 241: 	 assign_stmt_97_to_assign_stmt_1138/slice_326_Update/$entry
      -- CP-element group 241: 	 assign_stmt_97_to_assign_stmt_1138/slice_326_Update/cr
      -- 
    cr_1418_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1418_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(241), ack => slice_326_inst_req_1); -- 
    maxPool4_cp_element_group_241: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_241"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(243) & maxPool4_CP_346_elements(378);
      gj_maxPool4_cp_element_group_241 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(241), clk => clk, reset => reset); --
    end block;
    -- CP-element group 242:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	240 
    -- CP-element group 242: successors 
    -- CP-element group 242: marked-successors 
    -- CP-element group 242: 	45 
    -- CP-element group 242: 	240 
    -- CP-element group 242:  members (3) 
      -- CP-element group 242: 	 assign_stmt_97_to_assign_stmt_1138/slice_326_sample_completed_
      -- CP-element group 242: 	 assign_stmt_97_to_assign_stmt_1138/slice_326_Sample/$exit
      -- CP-element group 242: 	 assign_stmt_97_to_assign_stmt_1138/slice_326_Sample/ra
      -- 
    ra_1414_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 242_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_326_inst_ack_0, ack => maxPool4_CP_346_elements(242)); -- 
    -- CP-element group 243:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	241 
    -- CP-element group 243: successors 
    -- CP-element group 243: 	376 
    -- CP-element group 243: marked-successors 
    -- CP-element group 243: 	241 
    -- CP-element group 243:  members (3) 
      -- CP-element group 243: 	 assign_stmt_97_to_assign_stmt_1138/slice_326_update_completed_
      -- CP-element group 243: 	 assign_stmt_97_to_assign_stmt_1138/slice_326_Update/$exit
      -- CP-element group 243: 	 assign_stmt_97_to_assign_stmt_1138/slice_326_Update/ca
      -- 
    ca_1419_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 243_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_326_inst_ack_1, ack => maxPool4_CP_346_elements(243)); -- 
    -- CP-element group 244:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	51 
    -- CP-element group 244: marked-predecessors 
    -- CP-element group 244: 	246 
    -- CP-element group 244: successors 
    -- CP-element group 244: 	246 
    -- CP-element group 244:  members (3) 
      -- CP-element group 244: 	 assign_stmt_97_to_assign_stmt_1138/slice_330_sample_start_
      -- CP-element group 244: 	 assign_stmt_97_to_assign_stmt_1138/slice_330_Sample/$entry
      -- CP-element group 244: 	 assign_stmt_97_to_assign_stmt_1138/slice_330_Sample/rr
      -- 
    rr_1427_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1427_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(244), ack => slice_330_inst_req_0); -- 
    maxPool4_cp_element_group_244: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_244"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(51) & maxPool4_CP_346_elements(246);
      gj_maxPool4_cp_element_group_244 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(244), clk => clk, reset => reset); --
    end block;
    -- CP-element group 245:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: marked-predecessors 
    -- CP-element group 245: 	247 
    -- CP-element group 245: 	321 
    -- CP-element group 245: 	386 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	247 
    -- CP-element group 245:  members (3) 
      -- CP-element group 245: 	 assign_stmt_97_to_assign_stmt_1138/slice_330_update_start_
      -- CP-element group 245: 	 assign_stmt_97_to_assign_stmt_1138/slice_330_Update/$entry
      -- CP-element group 245: 	 assign_stmt_97_to_assign_stmt_1138/slice_330_Update/cr
      -- 
    cr_1432_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1432_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(245), ack => slice_330_inst_req_1); -- 
    maxPool4_cp_element_group_245: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_245"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(247) & maxPool4_CP_346_elements(321) & maxPool4_CP_346_elements(386);
      gj_maxPool4_cp_element_group_245 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(245), clk => clk, reset => reset); --
    end block;
    -- CP-element group 246:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	244 
    -- CP-element group 246: successors 
    -- CP-element group 246: marked-successors 
    -- CP-element group 246: 	49 
    -- CP-element group 246: 	244 
    -- CP-element group 246:  members (3) 
      -- CP-element group 246: 	 assign_stmt_97_to_assign_stmt_1138/slice_330_sample_completed_
      -- CP-element group 246: 	 assign_stmt_97_to_assign_stmt_1138/slice_330_Sample/$exit
      -- CP-element group 246: 	 assign_stmt_97_to_assign_stmt_1138/slice_330_Sample/ra
      -- 
    ra_1428_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 246_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_330_inst_ack_0, ack => maxPool4_CP_346_elements(246)); -- 
    -- CP-element group 247:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	245 
    -- CP-element group 247: successors 
    -- CP-element group 247: 	319 
    -- CP-element group 247: 	384 
    -- CP-element group 247: marked-successors 
    -- CP-element group 247: 	245 
    -- CP-element group 247:  members (3) 
      -- CP-element group 247: 	 assign_stmt_97_to_assign_stmt_1138/slice_330_update_completed_
      -- CP-element group 247: 	 assign_stmt_97_to_assign_stmt_1138/slice_330_Update/$exit
      -- CP-element group 247: 	 assign_stmt_97_to_assign_stmt_1138/slice_330_Update/ca
      -- 
    ca_1433_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 247_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_330_inst_ack_1, ack => maxPool4_CP_346_elements(247)); -- 
    -- CP-element group 248:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	51 
    -- CP-element group 248: marked-predecessors 
    -- CP-element group 248: 	250 
    -- CP-element group 248: successors 
    -- CP-element group 248: 	250 
    -- CP-element group 248:  members (3) 
      -- CP-element group 248: 	 assign_stmt_97_to_assign_stmt_1138/slice_334_sample_start_
      -- CP-element group 248: 	 assign_stmt_97_to_assign_stmt_1138/slice_334_Sample/$entry
      -- CP-element group 248: 	 assign_stmt_97_to_assign_stmt_1138/slice_334_Sample/rr
      -- 
    rr_1441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(248), ack => slice_334_inst_req_0); -- 
    maxPool4_cp_element_group_248: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_248"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(51) & maxPool4_CP_346_elements(250);
      gj_maxPool4_cp_element_group_248 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(248), clk => clk, reset => reset); --
    end block;
    -- CP-element group 249:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: marked-predecessors 
    -- CP-element group 249: 	251 
    -- CP-element group 249: 	321 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	251 
    -- CP-element group 249:  members (3) 
      -- CP-element group 249: 	 assign_stmt_97_to_assign_stmt_1138/slice_334_update_start_
      -- CP-element group 249: 	 assign_stmt_97_to_assign_stmt_1138/slice_334_Update/$entry
      -- CP-element group 249: 	 assign_stmt_97_to_assign_stmt_1138/slice_334_Update/cr
      -- 
    cr_1446_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1446_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(249), ack => slice_334_inst_req_1); -- 
    maxPool4_cp_element_group_249: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_249"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(251) & maxPool4_CP_346_elements(321);
      gj_maxPool4_cp_element_group_249 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(249), clk => clk, reset => reset); --
    end block;
    -- CP-element group 250:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	248 
    -- CP-element group 250: successors 
    -- CP-element group 250: marked-successors 
    -- CP-element group 250: 	49 
    -- CP-element group 250: 	248 
    -- CP-element group 250:  members (3) 
      -- CP-element group 250: 	 assign_stmt_97_to_assign_stmt_1138/slice_334_sample_completed_
      -- CP-element group 250: 	 assign_stmt_97_to_assign_stmt_1138/slice_334_Sample/$exit
      -- CP-element group 250: 	 assign_stmt_97_to_assign_stmt_1138/slice_334_Sample/ra
      -- 
    ra_1442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 250_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_334_inst_ack_0, ack => maxPool4_CP_346_elements(250)); -- 
    -- CP-element group 251:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	249 
    -- CP-element group 251: successors 
    -- CP-element group 251: 	319 
    -- CP-element group 251: marked-successors 
    -- CP-element group 251: 	249 
    -- CP-element group 251:  members (3) 
      -- CP-element group 251: 	 assign_stmt_97_to_assign_stmt_1138/slice_334_update_completed_
      -- CP-element group 251: 	 assign_stmt_97_to_assign_stmt_1138/slice_334_Update/$exit
      -- CP-element group 251: 	 assign_stmt_97_to_assign_stmt_1138/slice_334_Update/ca
      -- 
    ca_1447_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 251_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_334_inst_ack_1, ack => maxPool4_CP_346_elements(251)); -- 
    -- CP-element group 252:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	51 
    -- CP-element group 252: marked-predecessors 
    -- CP-element group 252: 	254 
    -- CP-element group 252: successors 
    -- CP-element group 252: 	254 
    -- CP-element group 252:  members (3) 
      -- CP-element group 252: 	 assign_stmt_97_to_assign_stmt_1138/slice_338_sample_start_
      -- CP-element group 252: 	 assign_stmt_97_to_assign_stmt_1138/slice_338_Sample/$entry
      -- CP-element group 252: 	 assign_stmt_97_to_assign_stmt_1138/slice_338_Sample/rr
      -- 
    rr_1455_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1455_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(252), ack => slice_338_inst_req_0); -- 
    maxPool4_cp_element_group_252: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_252"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(51) & maxPool4_CP_346_elements(254);
      gj_maxPool4_cp_element_group_252 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(252), clk => clk, reset => reset); --
    end block;
    -- CP-element group 253:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: marked-predecessors 
    -- CP-element group 253: 	255 
    -- CP-element group 253: 	321 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	255 
    -- CP-element group 253:  members (3) 
      -- CP-element group 253: 	 assign_stmt_97_to_assign_stmt_1138/slice_338_update_start_
      -- CP-element group 253: 	 assign_stmt_97_to_assign_stmt_1138/slice_338_Update/$entry
      -- CP-element group 253: 	 assign_stmt_97_to_assign_stmt_1138/slice_338_Update/cr
      -- 
    cr_1460_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1460_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(253), ack => slice_338_inst_req_1); -- 
    maxPool4_cp_element_group_253: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_253"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(255) & maxPool4_CP_346_elements(321);
      gj_maxPool4_cp_element_group_253 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(253), clk => clk, reset => reset); --
    end block;
    -- CP-element group 254:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	252 
    -- CP-element group 254: successors 
    -- CP-element group 254: marked-successors 
    -- CP-element group 254: 	49 
    -- CP-element group 254: 	252 
    -- CP-element group 254:  members (3) 
      -- CP-element group 254: 	 assign_stmt_97_to_assign_stmt_1138/slice_338_sample_completed_
      -- CP-element group 254: 	 assign_stmt_97_to_assign_stmt_1138/slice_338_Sample/$exit
      -- CP-element group 254: 	 assign_stmt_97_to_assign_stmt_1138/slice_338_Sample/ra
      -- 
    ra_1456_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 254_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_338_inst_ack_0, ack => maxPool4_CP_346_elements(254)); -- 
    -- CP-element group 255:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	253 
    -- CP-element group 255: successors 
    -- CP-element group 255: 	319 
    -- CP-element group 255: marked-successors 
    -- CP-element group 255: 	253 
    -- CP-element group 255:  members (3) 
      -- CP-element group 255: 	 assign_stmt_97_to_assign_stmt_1138/slice_338_update_completed_
      -- CP-element group 255: 	 assign_stmt_97_to_assign_stmt_1138/slice_338_Update/$exit
      -- CP-element group 255: 	 assign_stmt_97_to_assign_stmt_1138/slice_338_Update/ca
      -- 
    ca_1461_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 255_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_338_inst_ack_1, ack => maxPool4_CP_346_elements(255)); -- 
    -- CP-element group 256:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	51 
    -- CP-element group 256: marked-predecessors 
    -- CP-element group 256: 	258 
    -- CP-element group 256: successors 
    -- CP-element group 256: 	258 
    -- CP-element group 256:  members (3) 
      -- CP-element group 256: 	 assign_stmt_97_to_assign_stmt_1138/slice_342_sample_start_
      -- CP-element group 256: 	 assign_stmt_97_to_assign_stmt_1138/slice_342_Sample/$entry
      -- CP-element group 256: 	 assign_stmt_97_to_assign_stmt_1138/slice_342_Sample/rr
      -- 
    rr_1469_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1469_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(256), ack => slice_342_inst_req_0); -- 
    maxPool4_cp_element_group_256: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_256"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(51) & maxPool4_CP_346_elements(258);
      gj_maxPool4_cp_element_group_256 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(256), clk => clk, reset => reset); --
    end block;
    -- CP-element group 257:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: marked-predecessors 
    -- CP-element group 257: 	259 
    -- CP-element group 257: 	321 
    -- CP-element group 257: successors 
    -- CP-element group 257: 	259 
    -- CP-element group 257:  members (3) 
      -- CP-element group 257: 	 assign_stmt_97_to_assign_stmt_1138/slice_342_update_start_
      -- CP-element group 257: 	 assign_stmt_97_to_assign_stmt_1138/slice_342_Update/$entry
      -- CP-element group 257: 	 assign_stmt_97_to_assign_stmt_1138/slice_342_Update/cr
      -- 
    cr_1474_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1474_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(257), ack => slice_342_inst_req_1); -- 
    maxPool4_cp_element_group_257: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_257"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(259) & maxPool4_CP_346_elements(321);
      gj_maxPool4_cp_element_group_257 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(257), clk => clk, reset => reset); --
    end block;
    -- CP-element group 258:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	256 
    -- CP-element group 258: successors 
    -- CP-element group 258: marked-successors 
    -- CP-element group 258: 	49 
    -- CP-element group 258: 	256 
    -- CP-element group 258:  members (3) 
      -- CP-element group 258: 	 assign_stmt_97_to_assign_stmt_1138/slice_342_sample_completed_
      -- CP-element group 258: 	 assign_stmt_97_to_assign_stmt_1138/slice_342_Sample/$exit
      -- CP-element group 258: 	 assign_stmt_97_to_assign_stmt_1138/slice_342_Sample/ra
      -- 
    ra_1470_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 258_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_342_inst_ack_0, ack => maxPool4_CP_346_elements(258)); -- 
    -- CP-element group 259:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	257 
    -- CP-element group 259: successors 
    -- CP-element group 259: 	319 
    -- CP-element group 259: marked-successors 
    -- CP-element group 259: 	257 
    -- CP-element group 259:  members (3) 
      -- CP-element group 259: 	 assign_stmt_97_to_assign_stmt_1138/slice_342_update_completed_
      -- CP-element group 259: 	 assign_stmt_97_to_assign_stmt_1138/slice_342_Update/$exit
      -- CP-element group 259: 	 assign_stmt_97_to_assign_stmt_1138/slice_342_Update/ca
      -- 
    ca_1475_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 259_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_342_inst_ack_1, ack => maxPool4_CP_346_elements(259)); -- 
    -- CP-element group 260:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	51 
    -- CP-element group 260: marked-predecessors 
    -- CP-element group 260: 	262 
    -- CP-element group 260: successors 
    -- CP-element group 260: 	262 
    -- CP-element group 260:  members (3) 
      -- CP-element group 260: 	 assign_stmt_97_to_assign_stmt_1138/slice_346_sample_start_
      -- CP-element group 260: 	 assign_stmt_97_to_assign_stmt_1138/slice_346_Sample/$entry
      -- CP-element group 260: 	 assign_stmt_97_to_assign_stmt_1138/slice_346_Sample/rr
      -- 
    rr_1483_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1483_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(260), ack => slice_346_inst_req_0); -- 
    maxPool4_cp_element_group_260: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_260"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(51) & maxPool4_CP_346_elements(262);
      gj_maxPool4_cp_element_group_260 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(260), clk => clk, reset => reset); --
    end block;
    -- CP-element group 261:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: marked-predecessors 
    -- CP-element group 261: 	263 
    -- CP-element group 261: 	340 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	263 
    -- CP-element group 261:  members (3) 
      -- CP-element group 261: 	 assign_stmt_97_to_assign_stmt_1138/slice_346_update_start_
      -- CP-element group 261: 	 assign_stmt_97_to_assign_stmt_1138/slice_346_Update/$entry
      -- CP-element group 261: 	 assign_stmt_97_to_assign_stmt_1138/slice_346_Update/cr
      -- 
    cr_1488_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1488_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(261), ack => slice_346_inst_req_1); -- 
    maxPool4_cp_element_group_261: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_261"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(263) & maxPool4_CP_346_elements(340);
      gj_maxPool4_cp_element_group_261 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(261), clk => clk, reset => reset); --
    end block;
    -- CP-element group 262:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	260 
    -- CP-element group 262: successors 
    -- CP-element group 262: marked-successors 
    -- CP-element group 262: 	49 
    -- CP-element group 262: 	260 
    -- CP-element group 262:  members (3) 
      -- CP-element group 262: 	 assign_stmt_97_to_assign_stmt_1138/slice_346_sample_completed_
      -- CP-element group 262: 	 assign_stmt_97_to_assign_stmt_1138/slice_346_Sample/$exit
      -- CP-element group 262: 	 assign_stmt_97_to_assign_stmt_1138/slice_346_Sample/ra
      -- 
    ra_1484_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 262_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_346_inst_ack_0, ack => maxPool4_CP_346_elements(262)); -- 
    -- CP-element group 263:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	261 
    -- CP-element group 263: successors 
    -- CP-element group 263: 	338 
    -- CP-element group 263: marked-successors 
    -- CP-element group 263: 	261 
    -- CP-element group 263:  members (3) 
      -- CP-element group 263: 	 assign_stmt_97_to_assign_stmt_1138/slice_346_update_completed_
      -- CP-element group 263: 	 assign_stmt_97_to_assign_stmt_1138/slice_346_Update/$exit
      -- CP-element group 263: 	 assign_stmt_97_to_assign_stmt_1138/slice_346_Update/ca
      -- 
    ca_1489_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 263_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_346_inst_ack_1, ack => maxPool4_CP_346_elements(263)); -- 
    -- CP-element group 264:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	51 
    -- CP-element group 264: marked-predecessors 
    -- CP-element group 264: 	266 
    -- CP-element group 264: successors 
    -- CP-element group 264: 	266 
    -- CP-element group 264:  members (3) 
      -- CP-element group 264: 	 assign_stmt_97_to_assign_stmt_1138/slice_350_sample_start_
      -- CP-element group 264: 	 assign_stmt_97_to_assign_stmt_1138/slice_350_Sample/$entry
      -- CP-element group 264: 	 assign_stmt_97_to_assign_stmt_1138/slice_350_Sample/rr
      -- 
    rr_1497_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1497_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(264), ack => slice_350_inst_req_0); -- 
    maxPool4_cp_element_group_264: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_264"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(51) & maxPool4_CP_346_elements(266);
      gj_maxPool4_cp_element_group_264 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(264), clk => clk, reset => reset); --
    end block;
    -- CP-element group 265:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: marked-predecessors 
    -- CP-element group 265: 	267 
    -- CP-element group 265: 	340 
    -- CP-element group 265: successors 
    -- CP-element group 265: 	267 
    -- CP-element group 265:  members (3) 
      -- CP-element group 265: 	 assign_stmt_97_to_assign_stmt_1138/slice_350_update_start_
      -- CP-element group 265: 	 assign_stmt_97_to_assign_stmt_1138/slice_350_Update/$entry
      -- CP-element group 265: 	 assign_stmt_97_to_assign_stmt_1138/slice_350_Update/cr
      -- 
    cr_1502_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1502_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(265), ack => slice_350_inst_req_1); -- 
    maxPool4_cp_element_group_265: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_265"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(267) & maxPool4_CP_346_elements(340);
      gj_maxPool4_cp_element_group_265 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(265), clk => clk, reset => reset); --
    end block;
    -- CP-element group 266:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	264 
    -- CP-element group 266: successors 
    -- CP-element group 266: marked-successors 
    -- CP-element group 266: 	49 
    -- CP-element group 266: 	264 
    -- CP-element group 266:  members (3) 
      -- CP-element group 266: 	 assign_stmt_97_to_assign_stmt_1138/slice_350_sample_completed_
      -- CP-element group 266: 	 assign_stmt_97_to_assign_stmt_1138/slice_350_Sample/$exit
      -- CP-element group 266: 	 assign_stmt_97_to_assign_stmt_1138/slice_350_Sample/ra
      -- 
    ra_1498_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 266_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_350_inst_ack_0, ack => maxPool4_CP_346_elements(266)); -- 
    -- CP-element group 267:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	265 
    -- CP-element group 267: successors 
    -- CP-element group 267: 	338 
    -- CP-element group 267: marked-successors 
    -- CP-element group 267: 	265 
    -- CP-element group 267:  members (3) 
      -- CP-element group 267: 	 assign_stmt_97_to_assign_stmt_1138/slice_350_update_completed_
      -- CP-element group 267: 	 assign_stmt_97_to_assign_stmt_1138/slice_350_Update/$exit
      -- CP-element group 267: 	 assign_stmt_97_to_assign_stmt_1138/slice_350_Update/ca
      -- 
    ca_1503_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 267_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_350_inst_ack_1, ack => maxPool4_CP_346_elements(267)); -- 
    -- CP-element group 268:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	51 
    -- CP-element group 268: marked-predecessors 
    -- CP-element group 268: 	270 
    -- CP-element group 268: successors 
    -- CP-element group 268: 	270 
    -- CP-element group 268:  members (3) 
      -- CP-element group 268: 	 assign_stmt_97_to_assign_stmt_1138/slice_354_sample_start_
      -- CP-element group 268: 	 assign_stmt_97_to_assign_stmt_1138/slice_354_Sample/$entry
      -- CP-element group 268: 	 assign_stmt_97_to_assign_stmt_1138/slice_354_Sample/rr
      -- 
    rr_1511_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1511_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(268), ack => slice_354_inst_req_0); -- 
    maxPool4_cp_element_group_268: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_268"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(51) & maxPool4_CP_346_elements(270);
      gj_maxPool4_cp_element_group_268 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(268), clk => clk, reset => reset); --
    end block;
    -- CP-element group 269:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: marked-predecessors 
    -- CP-element group 269: 	271 
    -- CP-element group 269: 	340 
    -- CP-element group 269: successors 
    -- CP-element group 269: 	271 
    -- CP-element group 269:  members (3) 
      -- CP-element group 269: 	 assign_stmt_97_to_assign_stmt_1138/slice_354_update_start_
      -- CP-element group 269: 	 assign_stmt_97_to_assign_stmt_1138/slice_354_Update/$entry
      -- CP-element group 269: 	 assign_stmt_97_to_assign_stmt_1138/slice_354_Update/cr
      -- 
    cr_1516_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1516_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(269), ack => slice_354_inst_req_1); -- 
    maxPool4_cp_element_group_269: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_269"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(271) & maxPool4_CP_346_elements(340);
      gj_maxPool4_cp_element_group_269 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(269), clk => clk, reset => reset); --
    end block;
    -- CP-element group 270:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	268 
    -- CP-element group 270: successors 
    -- CP-element group 270: marked-successors 
    -- CP-element group 270: 	49 
    -- CP-element group 270: 	268 
    -- CP-element group 270:  members (3) 
      -- CP-element group 270: 	 assign_stmt_97_to_assign_stmt_1138/slice_354_sample_completed_
      -- CP-element group 270: 	 assign_stmt_97_to_assign_stmt_1138/slice_354_Sample/$exit
      -- CP-element group 270: 	 assign_stmt_97_to_assign_stmt_1138/slice_354_Sample/ra
      -- 
    ra_1512_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 270_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_354_inst_ack_0, ack => maxPool4_CP_346_elements(270)); -- 
    -- CP-element group 271:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	269 
    -- CP-element group 271: successors 
    -- CP-element group 271: 	338 
    -- CP-element group 271: marked-successors 
    -- CP-element group 271: 	269 
    -- CP-element group 271:  members (3) 
      -- CP-element group 271: 	 assign_stmt_97_to_assign_stmt_1138/slice_354_update_completed_
      -- CP-element group 271: 	 assign_stmt_97_to_assign_stmt_1138/slice_354_Update/$exit
      -- CP-element group 271: 	 assign_stmt_97_to_assign_stmt_1138/slice_354_Update/ca
      -- 
    ca_1517_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 271_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_354_inst_ack_1, ack => maxPool4_CP_346_elements(271)); -- 
    -- CP-element group 272:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	51 
    -- CP-element group 272: marked-predecessors 
    -- CP-element group 272: 	274 
    -- CP-element group 272: successors 
    -- CP-element group 272: 	274 
    -- CP-element group 272:  members (3) 
      -- CP-element group 272: 	 assign_stmt_97_to_assign_stmt_1138/slice_358_sample_start_
      -- CP-element group 272: 	 assign_stmt_97_to_assign_stmt_1138/slice_358_Sample/$entry
      -- CP-element group 272: 	 assign_stmt_97_to_assign_stmt_1138/slice_358_Sample/rr
      -- 
    rr_1525_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1525_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(272), ack => slice_358_inst_req_0); -- 
    maxPool4_cp_element_group_272: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_272"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(51) & maxPool4_CP_346_elements(274);
      gj_maxPool4_cp_element_group_272 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(272), clk => clk, reset => reset); --
    end block;
    -- CP-element group 273:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: marked-predecessors 
    -- CP-element group 273: 	275 
    -- CP-element group 273: 	340 
    -- CP-element group 273: successors 
    -- CP-element group 273: 	275 
    -- CP-element group 273:  members (3) 
      -- CP-element group 273: 	 assign_stmt_97_to_assign_stmt_1138/slice_358_update_start_
      -- CP-element group 273: 	 assign_stmt_97_to_assign_stmt_1138/slice_358_Update/$entry
      -- CP-element group 273: 	 assign_stmt_97_to_assign_stmt_1138/slice_358_Update/cr
      -- 
    cr_1530_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1530_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(273), ack => slice_358_inst_req_1); -- 
    maxPool4_cp_element_group_273: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_273"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(275) & maxPool4_CP_346_elements(340);
      gj_maxPool4_cp_element_group_273 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(273), clk => clk, reset => reset); --
    end block;
    -- CP-element group 274:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	272 
    -- CP-element group 274: successors 
    -- CP-element group 274: marked-successors 
    -- CP-element group 274: 	49 
    -- CP-element group 274: 	272 
    -- CP-element group 274:  members (3) 
      -- CP-element group 274: 	 assign_stmt_97_to_assign_stmt_1138/slice_358_sample_completed_
      -- CP-element group 274: 	 assign_stmt_97_to_assign_stmt_1138/slice_358_Sample/$exit
      -- CP-element group 274: 	 assign_stmt_97_to_assign_stmt_1138/slice_358_Sample/ra
      -- 
    ra_1526_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 274_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_358_inst_ack_0, ack => maxPool4_CP_346_elements(274)); -- 
    -- CP-element group 275:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	273 
    -- CP-element group 275: successors 
    -- CP-element group 275: 	338 
    -- CP-element group 275: marked-successors 
    -- CP-element group 275: 	273 
    -- CP-element group 275:  members (3) 
      -- CP-element group 275: 	 assign_stmt_97_to_assign_stmt_1138/slice_358_update_completed_
      -- CP-element group 275: 	 assign_stmt_97_to_assign_stmt_1138/slice_358_Update/$exit
      -- CP-element group 275: 	 assign_stmt_97_to_assign_stmt_1138/slice_358_Update/ca
      -- 
    ca_1531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 275_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_358_inst_ack_1, ack => maxPool4_CP_346_elements(275)); -- 
    -- CP-element group 276:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	51 
    -- CP-element group 276: marked-predecessors 
    -- CP-element group 276: 	278 
    -- CP-element group 276: successors 
    -- CP-element group 276: 	278 
    -- CP-element group 276:  members (3) 
      -- CP-element group 276: 	 assign_stmt_97_to_assign_stmt_1138/slice_362_Sample/rr
      -- CP-element group 276: 	 assign_stmt_97_to_assign_stmt_1138/slice_362_Sample/$entry
      -- CP-element group 276: 	 assign_stmt_97_to_assign_stmt_1138/slice_362_sample_start_
      -- 
    rr_1539_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1539_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(276), ack => slice_362_inst_req_0); -- 
    maxPool4_cp_element_group_276: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_276"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(51) & maxPool4_CP_346_elements(278);
      gj_maxPool4_cp_element_group_276 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(276), clk => clk, reset => reset); --
    end block;
    -- CP-element group 277:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: marked-predecessors 
    -- CP-element group 277: 	279 
    -- CP-element group 277: 	359 
    -- CP-element group 277: successors 
    -- CP-element group 277: 	279 
    -- CP-element group 277:  members (3) 
      -- CP-element group 277: 	 assign_stmt_97_to_assign_stmt_1138/slice_362_Update/cr
      -- CP-element group 277: 	 assign_stmt_97_to_assign_stmt_1138/slice_362_Update/$entry
      -- CP-element group 277: 	 assign_stmt_97_to_assign_stmt_1138/slice_362_update_start_
      -- 
    cr_1544_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1544_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(277), ack => slice_362_inst_req_1); -- 
    maxPool4_cp_element_group_277: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_277"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(279) & maxPool4_CP_346_elements(359);
      gj_maxPool4_cp_element_group_277 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(277), clk => clk, reset => reset); --
    end block;
    -- CP-element group 278:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	276 
    -- CP-element group 278: successors 
    -- CP-element group 278: marked-successors 
    -- CP-element group 278: 	49 
    -- CP-element group 278: 	276 
    -- CP-element group 278:  members (3) 
      -- CP-element group 278: 	 assign_stmt_97_to_assign_stmt_1138/slice_362_Sample/ra
      -- CP-element group 278: 	 assign_stmt_97_to_assign_stmt_1138/slice_362_Sample/$exit
      -- CP-element group 278: 	 assign_stmt_97_to_assign_stmt_1138/slice_362_sample_completed_
      -- 
    ra_1540_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 278_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_362_inst_ack_0, ack => maxPool4_CP_346_elements(278)); -- 
    -- CP-element group 279:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	277 
    -- CP-element group 279: successors 
    -- CP-element group 279: 	357 
    -- CP-element group 279: marked-successors 
    -- CP-element group 279: 	277 
    -- CP-element group 279:  members (3) 
      -- CP-element group 279: 	 assign_stmt_97_to_assign_stmt_1138/slice_362_Update/ca
      -- CP-element group 279: 	 assign_stmt_97_to_assign_stmt_1138/slice_362_Update/$exit
      -- CP-element group 279: 	 assign_stmt_97_to_assign_stmt_1138/slice_362_update_completed_
      -- 
    ca_1545_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 279_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_362_inst_ack_1, ack => maxPool4_CP_346_elements(279)); -- 
    -- CP-element group 280:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	51 
    -- CP-element group 280: marked-predecessors 
    -- CP-element group 280: 	282 
    -- CP-element group 280: successors 
    -- CP-element group 280: 	282 
    -- CP-element group 280:  members (3) 
      -- CP-element group 280: 	 assign_stmt_97_to_assign_stmt_1138/slice_366_Sample/rr
      -- CP-element group 280: 	 assign_stmt_97_to_assign_stmt_1138/slice_366_Sample/$entry
      -- CP-element group 280: 	 assign_stmt_97_to_assign_stmt_1138/slice_366_sample_start_
      -- 
    rr_1553_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1553_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(280), ack => slice_366_inst_req_0); -- 
    maxPool4_cp_element_group_280: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_280"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(51) & maxPool4_CP_346_elements(282);
      gj_maxPool4_cp_element_group_280 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(280), clk => clk, reset => reset); --
    end block;
    -- CP-element group 281:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: marked-predecessors 
    -- CP-element group 281: 	283 
    -- CP-element group 281: 	359 
    -- CP-element group 281: successors 
    -- CP-element group 281: 	283 
    -- CP-element group 281:  members (3) 
      -- CP-element group 281: 	 assign_stmt_97_to_assign_stmt_1138/slice_366_Update/cr
      -- CP-element group 281: 	 assign_stmt_97_to_assign_stmt_1138/slice_366_Update/$entry
      -- CP-element group 281: 	 assign_stmt_97_to_assign_stmt_1138/slice_366_update_start_
      -- 
    cr_1558_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1558_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(281), ack => slice_366_inst_req_1); -- 
    maxPool4_cp_element_group_281: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_281"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(283) & maxPool4_CP_346_elements(359);
      gj_maxPool4_cp_element_group_281 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(281), clk => clk, reset => reset); --
    end block;
    -- CP-element group 282:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	280 
    -- CP-element group 282: successors 
    -- CP-element group 282: marked-successors 
    -- CP-element group 282: 	49 
    -- CP-element group 282: 	280 
    -- CP-element group 282:  members (3) 
      -- CP-element group 282: 	 assign_stmt_97_to_assign_stmt_1138/slice_366_Sample/ra
      -- CP-element group 282: 	 assign_stmt_97_to_assign_stmt_1138/slice_366_Sample/$exit
      -- CP-element group 282: 	 assign_stmt_97_to_assign_stmt_1138/slice_366_sample_completed_
      -- 
    ra_1554_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 282_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_366_inst_ack_0, ack => maxPool4_CP_346_elements(282)); -- 
    -- CP-element group 283:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: 	281 
    -- CP-element group 283: successors 
    -- CP-element group 283: 	357 
    -- CP-element group 283: marked-successors 
    -- CP-element group 283: 	281 
    -- CP-element group 283:  members (3) 
      -- CP-element group 283: 	 assign_stmt_97_to_assign_stmt_1138/slice_366_Update/$exit
      -- CP-element group 283: 	 assign_stmt_97_to_assign_stmt_1138/slice_366_Update/ca
      -- CP-element group 283: 	 assign_stmt_97_to_assign_stmt_1138/slice_366_update_completed_
      -- 
    ca_1559_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 283_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_366_inst_ack_1, ack => maxPool4_CP_346_elements(283)); -- 
    -- CP-element group 284:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	51 
    -- CP-element group 284: marked-predecessors 
    -- CP-element group 284: 	286 
    -- CP-element group 284: successors 
    -- CP-element group 284: 	286 
    -- CP-element group 284:  members (3) 
      -- CP-element group 284: 	 assign_stmt_97_to_assign_stmt_1138/slice_370_Sample/$entry
      -- CP-element group 284: 	 assign_stmt_97_to_assign_stmt_1138/slice_370_Sample/rr
      -- CP-element group 284: 	 assign_stmt_97_to_assign_stmt_1138/slice_370_sample_start_
      -- 
    rr_1567_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1567_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(284), ack => slice_370_inst_req_0); -- 
    maxPool4_cp_element_group_284: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_284"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(51) & maxPool4_CP_346_elements(286);
      gj_maxPool4_cp_element_group_284 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(284), clk => clk, reset => reset); --
    end block;
    -- CP-element group 285:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: marked-predecessors 
    -- CP-element group 285: 	287 
    -- CP-element group 285: 	359 
    -- CP-element group 285: successors 
    -- CP-element group 285: 	287 
    -- CP-element group 285:  members (3) 
      -- CP-element group 285: 	 assign_stmt_97_to_assign_stmt_1138/slice_370_update_start_
      -- CP-element group 285: 	 assign_stmt_97_to_assign_stmt_1138/slice_370_Update/$entry
      -- CP-element group 285: 	 assign_stmt_97_to_assign_stmt_1138/slice_370_Update/cr
      -- 
    cr_1572_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1572_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(285), ack => slice_370_inst_req_1); -- 
    maxPool4_cp_element_group_285: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_285"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(287) & maxPool4_CP_346_elements(359);
      gj_maxPool4_cp_element_group_285 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(285), clk => clk, reset => reset); --
    end block;
    -- CP-element group 286:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	284 
    -- CP-element group 286: successors 
    -- CP-element group 286: marked-successors 
    -- CP-element group 286: 	49 
    -- CP-element group 286: 	284 
    -- CP-element group 286:  members (3) 
      -- CP-element group 286: 	 assign_stmt_97_to_assign_stmt_1138/slice_370_Sample/$exit
      -- CP-element group 286: 	 assign_stmt_97_to_assign_stmt_1138/slice_370_sample_completed_
      -- CP-element group 286: 	 assign_stmt_97_to_assign_stmt_1138/slice_370_Sample/ra
      -- 
    ra_1568_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 286_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_370_inst_ack_0, ack => maxPool4_CP_346_elements(286)); -- 
    -- CP-element group 287:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	285 
    -- CP-element group 287: successors 
    -- CP-element group 287: 	357 
    -- CP-element group 287: marked-successors 
    -- CP-element group 287: 	285 
    -- CP-element group 287:  members (3) 
      -- CP-element group 287: 	 assign_stmt_97_to_assign_stmt_1138/slice_370_update_completed_
      -- CP-element group 287: 	 assign_stmt_97_to_assign_stmt_1138/slice_370_Update/$exit
      -- CP-element group 287: 	 assign_stmt_97_to_assign_stmt_1138/slice_370_Update/ca
      -- 
    ca_1573_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 287_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_370_inst_ack_1, ack => maxPool4_CP_346_elements(287)); -- 
    -- CP-element group 288:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	51 
    -- CP-element group 288: marked-predecessors 
    -- CP-element group 288: 	290 
    -- CP-element group 288: successors 
    -- CP-element group 288: 	290 
    -- CP-element group 288:  members (3) 
      -- CP-element group 288: 	 assign_stmt_97_to_assign_stmt_1138/slice_374_sample_start_
      -- CP-element group 288: 	 assign_stmt_97_to_assign_stmt_1138/slice_374_Sample/$entry
      -- CP-element group 288: 	 assign_stmt_97_to_assign_stmt_1138/slice_374_Sample/rr
      -- 
    rr_1581_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1581_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(288), ack => slice_374_inst_req_0); -- 
    maxPool4_cp_element_group_288: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_288"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(51) & maxPool4_CP_346_elements(290);
      gj_maxPool4_cp_element_group_288 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(288), clk => clk, reset => reset); --
    end block;
    -- CP-element group 289:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: marked-predecessors 
    -- CP-element group 289: 	291 
    -- CP-element group 289: 	359 
    -- CP-element group 289: successors 
    -- CP-element group 289: 	291 
    -- CP-element group 289:  members (3) 
      -- CP-element group 289: 	 assign_stmt_97_to_assign_stmt_1138/slice_374_update_start_
      -- CP-element group 289: 	 assign_stmt_97_to_assign_stmt_1138/slice_374_Update/$entry
      -- CP-element group 289: 	 assign_stmt_97_to_assign_stmt_1138/slice_374_Update/cr
      -- 
    cr_1586_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1586_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(289), ack => slice_374_inst_req_1); -- 
    maxPool4_cp_element_group_289: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_289"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(291) & maxPool4_CP_346_elements(359);
      gj_maxPool4_cp_element_group_289 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(289), clk => clk, reset => reset); --
    end block;
    -- CP-element group 290:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: 	288 
    -- CP-element group 290: successors 
    -- CP-element group 290: marked-successors 
    -- CP-element group 290: 	49 
    -- CP-element group 290: 	288 
    -- CP-element group 290:  members (3) 
      -- CP-element group 290: 	 assign_stmt_97_to_assign_stmt_1138/slice_374_sample_completed_
      -- CP-element group 290: 	 assign_stmt_97_to_assign_stmt_1138/slice_374_Sample/$exit
      -- CP-element group 290: 	 assign_stmt_97_to_assign_stmt_1138/slice_374_Sample/ra
      -- 
    ra_1582_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 290_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_374_inst_ack_0, ack => maxPool4_CP_346_elements(290)); -- 
    -- CP-element group 291:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	289 
    -- CP-element group 291: successors 
    -- CP-element group 291: 	357 
    -- CP-element group 291: marked-successors 
    -- CP-element group 291: 	289 
    -- CP-element group 291:  members (3) 
      -- CP-element group 291: 	 assign_stmt_97_to_assign_stmt_1138/slice_374_update_completed_
      -- CP-element group 291: 	 assign_stmt_97_to_assign_stmt_1138/slice_374_Update/$exit
      -- CP-element group 291: 	 assign_stmt_97_to_assign_stmt_1138/slice_374_Update/ca
      -- 
    ca_1587_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 291_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_374_inst_ack_1, ack => maxPool4_CP_346_elements(291)); -- 
    -- CP-element group 292:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	51 
    -- CP-element group 292: marked-predecessors 
    -- CP-element group 292: 	294 
    -- CP-element group 292: successors 
    -- CP-element group 292: 	294 
    -- CP-element group 292:  members (3) 
      -- CP-element group 292: 	 assign_stmt_97_to_assign_stmt_1138/slice_378_sample_start_
      -- CP-element group 292: 	 assign_stmt_97_to_assign_stmt_1138/slice_378_Sample/$entry
      -- CP-element group 292: 	 assign_stmt_97_to_assign_stmt_1138/slice_378_Sample/rr
      -- 
    rr_1595_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1595_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(292), ack => slice_378_inst_req_0); -- 
    maxPool4_cp_element_group_292: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_292"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(51) & maxPool4_CP_346_elements(294);
      gj_maxPool4_cp_element_group_292 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(292), clk => clk, reset => reset); --
    end block;
    -- CP-element group 293:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: marked-predecessors 
    -- CP-element group 293: 	295 
    -- CP-element group 293: 	378 
    -- CP-element group 293: successors 
    -- CP-element group 293: 	295 
    -- CP-element group 293:  members (3) 
      -- CP-element group 293: 	 assign_stmt_97_to_assign_stmt_1138/slice_378_Update/$entry
      -- CP-element group 293: 	 assign_stmt_97_to_assign_stmt_1138/slice_378_Update/cr
      -- CP-element group 293: 	 assign_stmt_97_to_assign_stmt_1138/slice_378_update_start_
      -- 
    cr_1600_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1600_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(293), ack => slice_378_inst_req_1); -- 
    maxPool4_cp_element_group_293: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_293"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(295) & maxPool4_CP_346_elements(378);
      gj_maxPool4_cp_element_group_293 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(293), clk => clk, reset => reset); --
    end block;
    -- CP-element group 294:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: 	292 
    -- CP-element group 294: successors 
    -- CP-element group 294: marked-successors 
    -- CP-element group 294: 	49 
    -- CP-element group 294: 	292 
    -- CP-element group 294:  members (3) 
      -- CP-element group 294: 	 assign_stmt_97_to_assign_stmt_1138/slice_378_sample_completed_
      -- CP-element group 294: 	 assign_stmt_97_to_assign_stmt_1138/slice_378_Sample/$exit
      -- CP-element group 294: 	 assign_stmt_97_to_assign_stmt_1138/slice_378_Sample/ra
      -- 
    ra_1596_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 294_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_378_inst_ack_0, ack => maxPool4_CP_346_elements(294)); -- 
    -- CP-element group 295:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 295: predecessors 
    -- CP-element group 295: 	293 
    -- CP-element group 295: successors 
    -- CP-element group 295: 	376 
    -- CP-element group 295: marked-successors 
    -- CP-element group 295: 	293 
    -- CP-element group 295:  members (3) 
      -- CP-element group 295: 	 assign_stmt_97_to_assign_stmt_1138/slice_378_Update/$exit
      -- CP-element group 295: 	 assign_stmt_97_to_assign_stmt_1138/slice_378_Update/ca
      -- CP-element group 295: 	 assign_stmt_97_to_assign_stmt_1138/slice_378_update_completed_
      -- 
    ca_1601_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 295_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_378_inst_ack_1, ack => maxPool4_CP_346_elements(295)); -- 
    -- CP-element group 296:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 296: predecessors 
    -- CP-element group 296: 	51 
    -- CP-element group 296: marked-predecessors 
    -- CP-element group 296: 	298 
    -- CP-element group 296: successors 
    -- CP-element group 296: 	298 
    -- CP-element group 296:  members (3) 
      -- CP-element group 296: 	 assign_stmt_97_to_assign_stmt_1138/slice_382_sample_start_
      -- CP-element group 296: 	 assign_stmt_97_to_assign_stmt_1138/slice_382_Sample/rr
      -- CP-element group 296: 	 assign_stmt_97_to_assign_stmt_1138/slice_382_Sample/$entry
      -- 
    rr_1609_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1609_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(296), ack => slice_382_inst_req_0); -- 
    maxPool4_cp_element_group_296: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_296"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(51) & maxPool4_CP_346_elements(298);
      gj_maxPool4_cp_element_group_296 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(296), clk => clk, reset => reset); --
    end block;
    -- CP-element group 297:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 297: predecessors 
    -- CP-element group 297: marked-predecessors 
    -- CP-element group 297: 	299 
    -- CP-element group 297: 	378 
    -- CP-element group 297: successors 
    -- CP-element group 297: 	299 
    -- CP-element group 297:  members (3) 
      -- CP-element group 297: 	 assign_stmt_97_to_assign_stmt_1138/slice_382_update_start_
      -- CP-element group 297: 	 assign_stmt_97_to_assign_stmt_1138/slice_382_Update/cr
      -- CP-element group 297: 	 assign_stmt_97_to_assign_stmt_1138/slice_382_Update/$entry
      -- 
    cr_1614_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1614_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(297), ack => slice_382_inst_req_1); -- 
    maxPool4_cp_element_group_297: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_297"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(299) & maxPool4_CP_346_elements(378);
      gj_maxPool4_cp_element_group_297 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(297), clk => clk, reset => reset); --
    end block;
    -- CP-element group 298:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 298: predecessors 
    -- CP-element group 298: 	296 
    -- CP-element group 298: successors 
    -- CP-element group 298: marked-successors 
    -- CP-element group 298: 	49 
    -- CP-element group 298: 	296 
    -- CP-element group 298:  members (3) 
      -- CP-element group 298: 	 assign_stmt_97_to_assign_stmt_1138/slice_382_sample_completed_
      -- CP-element group 298: 	 assign_stmt_97_to_assign_stmt_1138/slice_382_Sample/$exit
      -- CP-element group 298: 	 assign_stmt_97_to_assign_stmt_1138/slice_382_Sample/ra
      -- 
    ra_1610_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 298_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_382_inst_ack_0, ack => maxPool4_CP_346_elements(298)); -- 
    -- CP-element group 299:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 299: predecessors 
    -- CP-element group 299: 	297 
    -- CP-element group 299: successors 
    -- CP-element group 299: 	376 
    -- CP-element group 299: marked-successors 
    -- CP-element group 299: 	297 
    -- CP-element group 299:  members (3) 
      -- CP-element group 299: 	 assign_stmt_97_to_assign_stmt_1138/slice_382_update_completed_
      -- CP-element group 299: 	 assign_stmt_97_to_assign_stmt_1138/slice_382_Update/ca
      -- CP-element group 299: 	 assign_stmt_97_to_assign_stmt_1138/slice_382_Update/$exit
      -- 
    ca_1615_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 299_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_382_inst_ack_1, ack => maxPool4_CP_346_elements(299)); -- 
    -- CP-element group 300:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 300: predecessors 
    -- CP-element group 300: 	51 
    -- CP-element group 300: marked-predecessors 
    -- CP-element group 300: 	302 
    -- CP-element group 300: successors 
    -- CP-element group 300: 	302 
    -- CP-element group 300:  members (3) 
      -- CP-element group 300: 	 assign_stmt_97_to_assign_stmt_1138/slice_386_Sample/rr
      -- CP-element group 300: 	 assign_stmt_97_to_assign_stmt_1138/slice_386_Sample/$entry
      -- CP-element group 300: 	 assign_stmt_97_to_assign_stmt_1138/slice_386_sample_start_
      -- 
    rr_1623_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1623_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(300), ack => slice_386_inst_req_0); -- 
    maxPool4_cp_element_group_300: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_300"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(51) & maxPool4_CP_346_elements(302);
      gj_maxPool4_cp_element_group_300 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(300), clk => clk, reset => reset); --
    end block;
    -- CP-element group 301:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 301: predecessors 
    -- CP-element group 301: marked-predecessors 
    -- CP-element group 301: 	303 
    -- CP-element group 301: 	378 
    -- CP-element group 301: successors 
    -- CP-element group 301: 	303 
    -- CP-element group 301:  members (3) 
      -- CP-element group 301: 	 assign_stmt_97_to_assign_stmt_1138/slice_386_Update/cr
      -- CP-element group 301: 	 assign_stmt_97_to_assign_stmt_1138/slice_386_Update/$entry
      -- CP-element group 301: 	 assign_stmt_97_to_assign_stmt_1138/slice_386_update_start_
      -- 
    cr_1628_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1628_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(301), ack => slice_386_inst_req_1); -- 
    maxPool4_cp_element_group_301: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_301"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(303) & maxPool4_CP_346_elements(378);
      gj_maxPool4_cp_element_group_301 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(301), clk => clk, reset => reset); --
    end block;
    -- CP-element group 302:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 302: predecessors 
    -- CP-element group 302: 	300 
    -- CP-element group 302: successors 
    -- CP-element group 302: marked-successors 
    -- CP-element group 302: 	49 
    -- CP-element group 302: 	300 
    -- CP-element group 302:  members (3) 
      -- CP-element group 302: 	 assign_stmt_97_to_assign_stmt_1138/slice_386_Sample/ra
      -- CP-element group 302: 	 assign_stmt_97_to_assign_stmt_1138/slice_386_Sample/$exit
      -- CP-element group 302: 	 assign_stmt_97_to_assign_stmt_1138/slice_386_sample_completed_
      -- 
    ra_1624_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 302_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_386_inst_ack_0, ack => maxPool4_CP_346_elements(302)); -- 
    -- CP-element group 303:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 303: predecessors 
    -- CP-element group 303: 	301 
    -- CP-element group 303: successors 
    -- CP-element group 303: 	376 
    -- CP-element group 303: marked-successors 
    -- CP-element group 303: 	301 
    -- CP-element group 303:  members (3) 
      -- CP-element group 303: 	 assign_stmt_97_to_assign_stmt_1138/slice_386_Update/ca
      -- CP-element group 303: 	 assign_stmt_97_to_assign_stmt_1138/slice_386_Update/$exit
      -- CP-element group 303: 	 assign_stmt_97_to_assign_stmt_1138/slice_386_update_completed_
      -- 
    ca_1629_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 303_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_386_inst_ack_1, ack => maxPool4_CP_346_elements(303)); -- 
    -- CP-element group 304:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 304: predecessors 
    -- CP-element group 304: 	51 
    -- CP-element group 304: marked-predecessors 
    -- CP-element group 304: 	306 
    -- CP-element group 304: successors 
    -- CP-element group 304: 	306 
    -- CP-element group 304:  members (3) 
      -- CP-element group 304: 	 assign_stmt_97_to_assign_stmt_1138/slice_390_Sample/rr
      -- CP-element group 304: 	 assign_stmt_97_to_assign_stmt_1138/slice_390_Sample/$entry
      -- CP-element group 304: 	 assign_stmt_97_to_assign_stmt_1138/slice_390_sample_start_
      -- 
    rr_1637_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1637_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(304), ack => slice_390_inst_req_0); -- 
    maxPool4_cp_element_group_304: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_304"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(51) & maxPool4_CP_346_elements(306);
      gj_maxPool4_cp_element_group_304 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(304), clk => clk, reset => reset); --
    end block;
    -- CP-element group 305:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 305: predecessors 
    -- CP-element group 305: marked-predecessors 
    -- CP-element group 305: 	307 
    -- CP-element group 305: 	378 
    -- CP-element group 305: successors 
    -- CP-element group 305: 	307 
    -- CP-element group 305:  members (3) 
      -- CP-element group 305: 	 assign_stmt_97_to_assign_stmt_1138/slice_390_Update/$entry
      -- CP-element group 305: 	 assign_stmt_97_to_assign_stmt_1138/slice_390_Update/cr
      -- CP-element group 305: 	 assign_stmt_97_to_assign_stmt_1138/slice_390_update_start_
      -- 
    cr_1642_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1642_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(305), ack => slice_390_inst_req_1); -- 
    maxPool4_cp_element_group_305: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_305"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(307) & maxPool4_CP_346_elements(378);
      gj_maxPool4_cp_element_group_305 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(305), clk => clk, reset => reset); --
    end block;
    -- CP-element group 306:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 306: predecessors 
    -- CP-element group 306: 	304 
    -- CP-element group 306: successors 
    -- CP-element group 306: marked-successors 
    -- CP-element group 306: 	49 
    -- CP-element group 306: 	304 
    -- CP-element group 306:  members (3) 
      -- CP-element group 306: 	 assign_stmt_97_to_assign_stmt_1138/slice_390_Sample/ra
      -- CP-element group 306: 	 assign_stmt_97_to_assign_stmt_1138/slice_390_Sample/$exit
      -- CP-element group 306: 	 assign_stmt_97_to_assign_stmt_1138/slice_390_sample_completed_
      -- 
    ra_1638_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 306_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_390_inst_ack_0, ack => maxPool4_CP_346_elements(306)); -- 
    -- CP-element group 307:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 307: predecessors 
    -- CP-element group 307: 	305 
    -- CP-element group 307: successors 
    -- CP-element group 307: 	376 
    -- CP-element group 307: marked-successors 
    -- CP-element group 307: 	305 
    -- CP-element group 307:  members (3) 
      -- CP-element group 307: 	 assign_stmt_97_to_assign_stmt_1138/slice_390_Update/$exit
      -- CP-element group 307: 	 assign_stmt_97_to_assign_stmt_1138/slice_390_Update/ca
      -- CP-element group 307: 	 assign_stmt_97_to_assign_stmt_1138/slice_390_update_completed_
      -- 
    ca_1643_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 307_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_390_inst_ack_1, ack => maxPool4_CP_346_elements(307)); -- 
    -- CP-element group 308:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 308: predecessors 
    -- CP-element group 308: 	312 
    -- CP-element group 308: marked-predecessors 
    -- CP-element group 308: 	313 
    -- CP-element group 308: successors 
    -- CP-element group 308: 	313 
    -- CP-element group 308:  members (3) 
      -- CP-element group 308: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_1038_sample_start_
      -- CP-element group 308: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_1038_request/$entry
      -- CP-element group 308: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_1038_request/req
      -- 
    req_1683_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1683_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(308), ack => addr_of_1038_final_reg_req_0); -- 
    maxPool4_cp_element_group_308: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_308"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(312) & maxPool4_CP_346_elements(313);
      gj_maxPool4_cp_element_group_308 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(308), clk => clk, reset => reset); --
    end block;
    -- CP-element group 309:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 309: predecessors 
    -- CP-element group 309: 	1 
    -- CP-element group 309: marked-predecessors 
    -- CP-element group 309: 	314 
    -- CP-element group 309: 	317 
    -- CP-element group 309: successors 
    -- CP-element group 309: 	314 
    -- CP-element group 309:  members (3) 
      -- CP-element group 309: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_1038_update_start_
      -- CP-element group 309: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_1038_complete/$entry
      -- CP-element group 309: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_1038_complete/req
      -- 
    req_1688_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1688_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(309), ack => addr_of_1038_final_reg_req_1); -- 
    maxPool4_cp_element_group_309: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_309"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(1) & maxPool4_CP_346_elements(314) & maxPool4_CP_346_elements(317);
      gj_maxPool4_cp_element_group_309 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(309), clk => clk, reset => reset); --
    end block;
    -- CP-element group 310:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 310: predecessors 
    -- CP-element group 310: 	1 
    -- CP-element group 310: marked-predecessors 
    -- CP-element group 310: 	312 
    -- CP-element group 310: 	313 
    -- CP-element group 310: successors 
    -- CP-element group 310: 	312 
    -- CP-element group 310:  members (3) 
      -- CP-element group 310: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1037_final_index_sum_regn_update_start
      -- CP-element group 310: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1037_final_index_sum_regn_Update/$entry
      -- CP-element group 310: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1037_final_index_sum_regn_Update/req
      -- 
    req_1673_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1673_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(310), ack => array_obj_ref_1037_index_offset_req_1); -- 
    maxPool4_cp_element_group_310: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_310"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(1) & maxPool4_CP_346_elements(312) & maxPool4_CP_346_elements(313);
      gj_maxPool4_cp_element_group_310 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(310), clk => clk, reset => reset); --
    end block;
    -- CP-element group 311:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 311: predecessors 
    -- CP-element group 311: 	1 
    -- CP-element group 311: successors 
    -- CP-element group 311: 	391 
    -- CP-element group 311: marked-successors 
    -- CP-element group 311: 	2 
    -- CP-element group 311:  members (3) 
      -- CP-element group 311: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1037_final_index_sum_regn_sample_complete
      -- CP-element group 311: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1037_final_index_sum_regn_Sample/$exit
      -- CP-element group 311: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1037_final_index_sum_regn_Sample/ack
      -- 
    ack_1669_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 311_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1037_index_offset_ack_0, ack => maxPool4_CP_346_elements(311)); -- 
    -- CP-element group 312:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 312: predecessors 
    -- CP-element group 312: 	310 
    -- CP-element group 312: successors 
    -- CP-element group 312: 	308 
    -- CP-element group 312: marked-successors 
    -- CP-element group 312: 	310 
    -- CP-element group 312:  members (8) 
      -- CP-element group 312: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1037_root_address_calculated
      -- CP-element group 312: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1037_offset_calculated
      -- CP-element group 312: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1037_base_plus_offset/sum_rename_req
      -- CP-element group 312: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1037_final_index_sum_regn_Update/$exit
      -- CP-element group 312: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1037_final_index_sum_regn_Update/ack
      -- CP-element group 312: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1037_base_plus_offset/$entry
      -- CP-element group 312: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1037_base_plus_offset/$exit
      -- CP-element group 312: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1037_base_plus_offset/sum_rename_ack
      -- 
    ack_1674_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 312_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1037_index_offset_ack_1, ack => maxPool4_CP_346_elements(312)); -- 
    -- CP-element group 313:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 313: predecessors 
    -- CP-element group 313: 	308 
    -- CP-element group 313: successors 
    -- CP-element group 313: marked-successors 
    -- CP-element group 313: 	308 
    -- CP-element group 313: 	310 
    -- CP-element group 313:  members (3) 
      -- CP-element group 313: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_1038_sample_completed_
      -- CP-element group 313: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_1038_request/$exit
      -- CP-element group 313: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_1038_request/ack
      -- 
    ack_1684_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 313_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1038_final_reg_ack_0, ack => maxPool4_CP_346_elements(313)); -- 
    -- CP-element group 314:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 314: predecessors 
    -- CP-element group 314: 	309 
    -- CP-element group 314: successors 
    -- CP-element group 314: 	315 
    -- CP-element group 314: marked-successors 
    -- CP-element group 314: 	309 
    -- CP-element group 314:  members (3) 
      -- CP-element group 314: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_1038_update_completed_
      -- CP-element group 314: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_1038_complete/$exit
      -- CP-element group 314: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_1038_complete/ack
      -- 
    ack_1689_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 314_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1038_final_reg_ack_1, ack => maxPool4_CP_346_elements(314)); -- 
    -- CP-element group 315:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 315: predecessors 
    -- CP-element group 315: 	314 
    -- CP-element group 315: marked-predecessors 
    -- CP-element group 315: 	317 
    -- CP-element group 315: successors 
    -- CP-element group 315: 	317 
    -- CP-element group 315:  members (3) 
      -- CP-element group 315: 	 assign_stmt_97_to_assign_stmt_1138/assign_stmt_1042_Sample/$entry
      -- CP-element group 315: 	 assign_stmt_97_to_assign_stmt_1138/assign_stmt_1042_Sample/req
      -- CP-element group 315: 	 assign_stmt_97_to_assign_stmt_1138/assign_stmt_1042_sample_start_
      -- 
    req_1697_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1697_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(315), ack => W_myptr5_1040_delayed_8_0_1040_inst_req_0); -- 
    maxPool4_cp_element_group_315: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_315"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(314) & maxPool4_CP_346_elements(317);
      gj_maxPool4_cp_element_group_315 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(315), clk => clk, reset => reset); --
    end block;
    -- CP-element group 316:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 316: predecessors 
    -- CP-element group 316: marked-predecessors 
    -- CP-element group 316: 	318 
    -- CP-element group 316: 	325 
    -- CP-element group 316: successors 
    -- CP-element group 316: 	318 
    -- CP-element group 316:  members (3) 
      -- CP-element group 316: 	 assign_stmt_97_to_assign_stmt_1138/assign_stmt_1042_Update/$entry
      -- CP-element group 316: 	 assign_stmt_97_to_assign_stmt_1138/assign_stmt_1042_update_start_
      -- CP-element group 316: 	 assign_stmt_97_to_assign_stmt_1138/assign_stmt_1042_Update/req
      -- 
    req_1702_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1702_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(316), ack => W_myptr5_1040_delayed_8_0_1040_inst_req_1); -- 
    maxPool4_cp_element_group_316: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_316"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(318) & maxPool4_CP_346_elements(325);
      gj_maxPool4_cp_element_group_316 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(316), clk => clk, reset => reset); --
    end block;
    -- CP-element group 317:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 317: predecessors 
    -- CP-element group 317: 	315 
    -- CP-element group 317: successors 
    -- CP-element group 317: marked-successors 
    -- CP-element group 317: 	309 
    -- CP-element group 317: 	315 
    -- CP-element group 317:  members (3) 
      -- CP-element group 317: 	 assign_stmt_97_to_assign_stmt_1138/assign_stmt_1042_Sample/ack
      -- CP-element group 317: 	 assign_stmt_97_to_assign_stmt_1138/assign_stmt_1042_Sample/$exit
      -- CP-element group 317: 	 assign_stmt_97_to_assign_stmt_1138/assign_stmt_1042_sample_completed_
      -- 
    ack_1698_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 317_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_myptr5_1040_delayed_8_0_1040_inst_ack_0, ack => maxPool4_CP_346_elements(317)); -- 
    -- CP-element group 318:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 318: predecessors 
    -- CP-element group 318: 	316 
    -- CP-element group 318: successors 
    -- CP-element group 318: 	323 
    -- CP-element group 318: marked-successors 
    -- CP-element group 318: 	316 
    -- CP-element group 318:  members (19) 
      -- CP-element group 318: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1044_base_addr_resize/base_resize_ack
      -- CP-element group 318: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1044_base_plus_offset/$entry
      -- CP-element group 318: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1044_base_addr_resize/base_resize_req
      -- CP-element group 318: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1044_base_plus_offset/$exit
      -- CP-element group 318: 	 assign_stmt_97_to_assign_stmt_1138/assign_stmt_1042_update_completed_
      -- CP-element group 318: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1044_base_addr_resize/$exit
      -- CP-element group 318: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1044_base_plus_offset/sum_rename_req
      -- CP-element group 318: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1044_base_address_calculated
      -- CP-element group 318: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1044_base_address_resized
      -- CP-element group 318: 	 assign_stmt_97_to_assign_stmt_1138/assign_stmt_1042_Update/$exit
      -- CP-element group 318: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1044_base_addr_resize/$entry
      -- CP-element group 318: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1044_base_plus_offset/sum_rename_ack
      -- CP-element group 318: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1044_root_address_calculated
      -- CP-element group 318: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1044_word_address_calculated
      -- CP-element group 318: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1044_word_addrgen/$entry
      -- CP-element group 318: 	 assign_stmt_97_to_assign_stmt_1138/assign_stmt_1042_Update/ack
      -- CP-element group 318: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1044_word_addrgen/$exit
      -- CP-element group 318: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1044_word_addrgen/root_register_req
      -- CP-element group 318: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1044_word_addrgen/root_register_ack
      -- 
    ack_1703_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 318_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_myptr5_1040_delayed_8_0_1040_inst_ack_1, ack => maxPool4_CP_346_elements(318)); -- 
    -- CP-element group 319:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 319: predecessors 
    -- CP-element group 319: 	55 
    -- CP-element group 319: 	59 
    -- CP-element group 319: 	63 
    -- CP-element group 319: 	67 
    -- CP-element group 319: 	119 
    -- CP-element group 319: 	123 
    -- CP-element group 319: 	127 
    -- CP-element group 319: 	131 
    -- CP-element group 319: 	183 
    -- CP-element group 319: 	187 
    -- CP-element group 319: 	191 
    -- CP-element group 319: 	195 
    -- CP-element group 319: 	247 
    -- CP-element group 319: 	251 
    -- CP-element group 319: 	255 
    -- CP-element group 319: 	259 
    -- CP-element group 319: marked-predecessors 
    -- CP-element group 319: 	321 
    -- CP-element group 319: successors 
    -- CP-element group 319: 	321 
    -- CP-element group 319:  members (3) 
      -- CP-element group 319: 	 assign_stmt_97_to_assign_stmt_1138/CONCAT_u32_u64_1055_sample_start_
      -- CP-element group 319: 	 assign_stmt_97_to_assign_stmt_1138/CONCAT_u32_u64_1055_Sample/$entry
      -- CP-element group 319: 	 assign_stmt_97_to_assign_stmt_1138/CONCAT_u32_u64_1055_Sample/rr
      -- 
    rr_1711_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1711_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(319), ack => CONCAT_u32_u64_1055_inst_req_0); -- 
    maxPool4_cp_element_group_319: block -- 
      constant place_capacities: IntegerArray(0 to 16) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_markings: IntegerArray(0 to 16)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 1);
      constant place_delays: IntegerArray(0 to 16) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_319"; 
      signal preds: BooleanArray(1 to 17); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(55) & maxPool4_CP_346_elements(59) & maxPool4_CP_346_elements(63) & maxPool4_CP_346_elements(67) & maxPool4_CP_346_elements(119) & maxPool4_CP_346_elements(123) & maxPool4_CP_346_elements(127) & maxPool4_CP_346_elements(131) & maxPool4_CP_346_elements(183) & maxPool4_CP_346_elements(187) & maxPool4_CP_346_elements(191) & maxPool4_CP_346_elements(195) & maxPool4_CP_346_elements(247) & maxPool4_CP_346_elements(251) & maxPool4_CP_346_elements(255) & maxPool4_CP_346_elements(259) & maxPool4_CP_346_elements(321);
      gj_maxPool4_cp_element_group_319 : generic_join generic map(name => joinName, number_of_predecessors => 17, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(319), clk => clk, reset => reset); --
    end block;
    -- CP-element group 320:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 320: predecessors 
    -- CP-element group 320: marked-predecessors 
    -- CP-element group 320: 	322 
    -- CP-element group 320: 	325 
    -- CP-element group 320: successors 
    -- CP-element group 320: 	322 
    -- CP-element group 320:  members (3) 
      -- CP-element group 320: 	 assign_stmt_97_to_assign_stmt_1138/CONCAT_u32_u64_1055_update_start_
      -- CP-element group 320: 	 assign_stmt_97_to_assign_stmt_1138/CONCAT_u32_u64_1055_Update/$entry
      -- CP-element group 320: 	 assign_stmt_97_to_assign_stmt_1138/CONCAT_u32_u64_1055_Update/cr
      -- 
    cr_1716_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1716_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(320), ack => CONCAT_u32_u64_1055_inst_req_1); -- 
    maxPool4_cp_element_group_320: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_320"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(322) & maxPool4_CP_346_elements(325);
      gj_maxPool4_cp_element_group_320 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(320), clk => clk, reset => reset); --
    end block;
    -- CP-element group 321:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 321: predecessors 
    -- CP-element group 321: 	319 
    -- CP-element group 321: successors 
    -- CP-element group 321: marked-successors 
    -- CP-element group 321: 	53 
    -- CP-element group 321: 	57 
    -- CP-element group 321: 	61 
    -- CP-element group 321: 	65 
    -- CP-element group 321: 	117 
    -- CP-element group 321: 	121 
    -- CP-element group 321: 	125 
    -- CP-element group 321: 	129 
    -- CP-element group 321: 	181 
    -- CP-element group 321: 	185 
    -- CP-element group 321: 	189 
    -- CP-element group 321: 	193 
    -- CP-element group 321: 	245 
    -- CP-element group 321: 	249 
    -- CP-element group 321: 	253 
    -- CP-element group 321: 	257 
    -- CP-element group 321: 	319 
    -- CP-element group 321:  members (3) 
      -- CP-element group 321: 	 assign_stmt_97_to_assign_stmt_1138/CONCAT_u32_u64_1055_sample_completed_
      -- CP-element group 321: 	 assign_stmt_97_to_assign_stmt_1138/CONCAT_u32_u64_1055_Sample/$exit
      -- CP-element group 321: 	 assign_stmt_97_to_assign_stmt_1138/CONCAT_u32_u64_1055_Sample/ra
      -- 
    ra_1712_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 321_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u32_u64_1055_inst_ack_0, ack => maxPool4_CP_346_elements(321)); -- 
    -- CP-element group 322:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 322: predecessors 
    -- CP-element group 322: 	320 
    -- CP-element group 322: successors 
    -- CP-element group 322: 	323 
    -- CP-element group 322: marked-successors 
    -- CP-element group 322: 	320 
    -- CP-element group 322:  members (3) 
      -- CP-element group 322: 	 assign_stmt_97_to_assign_stmt_1138/CONCAT_u32_u64_1055_update_completed_
      -- CP-element group 322: 	 assign_stmt_97_to_assign_stmt_1138/CONCAT_u32_u64_1055_Update/$exit
      -- CP-element group 322: 	 assign_stmt_97_to_assign_stmt_1138/CONCAT_u32_u64_1055_Update/ca
      -- 
    ca_1717_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 322_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u32_u64_1055_inst_ack_1, ack => maxPool4_CP_346_elements(322)); -- 
    -- CP-element group 323:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 323: predecessors 
    -- CP-element group 323: 	318 
    -- CP-element group 323: 	322 
    -- CP-element group 323: marked-predecessors 
    -- CP-element group 323: 	325 
    -- CP-element group 323: 	382 
    -- CP-element group 323: successors 
    -- CP-element group 323: 	325 
    -- CP-element group 323:  members (9) 
      -- CP-element group 323: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1044_Sample/$entry
      -- CP-element group 323: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1044_Sample/ptr_deref_1044_Split/$entry
      -- CP-element group 323: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1044_Sample/ptr_deref_1044_Split/$exit
      -- CP-element group 323: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1044_Sample/ptr_deref_1044_Split/split_req
      -- CP-element group 323: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1044_Sample/ptr_deref_1044_Split/split_ack
      -- CP-element group 323: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1044_Sample/word_access_start/$entry
      -- CP-element group 323: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1044_Sample/word_access_start/word_0/$entry
      -- CP-element group 323: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1044_Sample/word_access_start/word_0/rr
      -- CP-element group 323: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1044_sample_start_
      -- 
    rr_1755_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1755_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(323), ack => ptr_deref_1044_store_0_req_0); -- 
    maxPool4_cp_element_group_323: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 1,3 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_323"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(318) & maxPool4_CP_346_elements(322) & maxPool4_CP_346_elements(325) & maxPool4_CP_346_elements(382);
      gj_maxPool4_cp_element_group_323 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(323), clk => clk, reset => reset); --
    end block;
    -- CP-element group 324:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 324: predecessors 
    -- CP-element group 324: marked-predecessors 
    -- CP-element group 324: 	326 
    -- CP-element group 324: successors 
    -- CP-element group 324: 	326 
    -- CP-element group 324:  members (5) 
      -- CP-element group 324: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1044_Update/$entry
      -- CP-element group 324: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1044_Update/word_access_complete/$entry
      -- CP-element group 324: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1044_Update/word_access_complete/word_0/$entry
      -- CP-element group 324: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1044_Update/word_access_complete/word_0/cr
      -- CP-element group 324: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1044_update_start_
      -- 
    cr_1766_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1766_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(324), ack => ptr_deref_1044_store_0_req_1); -- 
    maxPool4_cp_element_group_324: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_324"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= maxPool4_CP_346_elements(326);
      gj_maxPool4_cp_element_group_324 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(324), clk => clk, reset => reset); --
    end block;
    -- CP-element group 325:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 325: predecessors 
    -- CP-element group 325: 	323 
    -- CP-element group 325: successors 
    -- CP-element group 325: 	388 
    -- CP-element group 325: marked-successors 
    -- CP-element group 325: 	316 
    -- CP-element group 325: 	320 
    -- CP-element group 325: 	323 
    -- CP-element group 325:  members (5) 
      -- CP-element group 325: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1044_Sample/$exit
      -- CP-element group 325: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1044_Sample/word_access_start/$exit
      -- CP-element group 325: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1044_Sample/word_access_start/word_0/$exit
      -- CP-element group 325: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1044_Sample/word_access_start/word_0/ra
      -- CP-element group 325: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1044_sample_completed_
      -- 
    ra_1756_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 325_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1044_store_0_ack_0, ack => maxPool4_CP_346_elements(325)); -- 
    -- CP-element group 326:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 326: predecessors 
    -- CP-element group 326: 	324 
    -- CP-element group 326: successors 
    -- CP-element group 326: 	391 
    -- CP-element group 326: marked-successors 
    -- CP-element group 326: 	324 
    -- CP-element group 326:  members (5) 
      -- CP-element group 326: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1044_update_completed_
      -- CP-element group 326: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1044_Update/$exit
      -- CP-element group 326: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1044_Update/word_access_complete/$exit
      -- CP-element group 326: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1044_Update/word_access_complete/word_0/$exit
      -- CP-element group 326: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1044_Update/word_access_complete/word_0/ca
      -- 
    ca_1767_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 326_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1044_store_0_ack_1, ack => maxPool4_CP_346_elements(326)); -- 
    -- CP-element group 327:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 327: predecessors 
    -- CP-element group 327: 	331 
    -- CP-element group 327: marked-predecessors 
    -- CP-element group 327: 	332 
    -- CP-element group 327: successors 
    -- CP-element group 327: 	332 
    -- CP-element group 327:  members (3) 
      -- CP-element group 327: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_1064_request/req
      -- CP-element group 327: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_1064_request/$entry
      -- CP-element group 327: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_1064_sample_start_
      -- 
    req_1807_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1807_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(327), ack => addr_of_1064_final_reg_req_0); -- 
    maxPool4_cp_element_group_327: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_327"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(331) & maxPool4_CP_346_elements(332);
      gj_maxPool4_cp_element_group_327 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(327), clk => clk, reset => reset); --
    end block;
    -- CP-element group 328:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 328: predecessors 
    -- CP-element group 328: 	1 
    -- CP-element group 328: marked-predecessors 
    -- CP-element group 328: 	333 
    -- CP-element group 328: 	336 
    -- CP-element group 328: successors 
    -- CP-element group 328: 	333 
    -- CP-element group 328:  members (3) 
      -- CP-element group 328: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_1064_complete/$entry
      -- CP-element group 328: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_1064_complete/req
      -- CP-element group 328: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_1064_update_start_
      -- 
    req_1812_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1812_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(328), ack => addr_of_1064_final_reg_req_1); -- 
    maxPool4_cp_element_group_328: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_328"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(1) & maxPool4_CP_346_elements(333) & maxPool4_CP_346_elements(336);
      gj_maxPool4_cp_element_group_328 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(328), clk => clk, reset => reset); --
    end block;
    -- CP-element group 329:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 329: predecessors 
    -- CP-element group 329: 	1 
    -- CP-element group 329: marked-predecessors 
    -- CP-element group 329: 	331 
    -- CP-element group 329: 	332 
    -- CP-element group 329: successors 
    -- CP-element group 329: 	331 
    -- CP-element group 329:  members (3) 
      -- CP-element group 329: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1063_final_index_sum_regn_Update/$entry
      -- CP-element group 329: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1063_final_index_sum_regn_update_start
      -- CP-element group 329: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1063_final_index_sum_regn_Update/req
      -- 
    req_1797_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1797_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(329), ack => array_obj_ref_1063_index_offset_req_1); -- 
    maxPool4_cp_element_group_329: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_329"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(1) & maxPool4_CP_346_elements(331) & maxPool4_CP_346_elements(332);
      gj_maxPool4_cp_element_group_329 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(329), clk => clk, reset => reset); --
    end block;
    -- CP-element group 330:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 330: predecessors 
    -- CP-element group 330: 	1 
    -- CP-element group 330: successors 
    -- CP-element group 330: 	391 
    -- CP-element group 330: marked-successors 
    -- CP-element group 330: 	2 
    -- CP-element group 330:  members (3) 
      -- CP-element group 330: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1063_final_index_sum_regn_sample_complete
      -- CP-element group 330: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1063_final_index_sum_regn_Sample/$exit
      -- CP-element group 330: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1063_final_index_sum_regn_Sample/ack
      -- 
    ack_1793_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 330_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1063_index_offset_ack_0, ack => maxPool4_CP_346_elements(330)); -- 
    -- CP-element group 331:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 331: predecessors 
    -- CP-element group 331: 	329 
    -- CP-element group 331: successors 
    -- CP-element group 331: 	327 
    -- CP-element group 331: marked-successors 
    -- CP-element group 331: 	329 
    -- CP-element group 331:  members (8) 
      -- CP-element group 331: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1063_final_index_sum_regn_Update/$exit
      -- CP-element group 331: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1063_base_plus_offset/$entry
      -- CP-element group 331: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1063_base_plus_offset/$exit
      -- CP-element group 331: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1063_base_plus_offset/sum_rename_req
      -- CP-element group 331: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1063_base_plus_offset/sum_rename_ack
      -- CP-element group 331: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1063_final_index_sum_regn_Update/ack
      -- CP-element group 331: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1063_offset_calculated
      -- CP-element group 331: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1063_root_address_calculated
      -- 
    ack_1798_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 331_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1063_index_offset_ack_1, ack => maxPool4_CP_346_elements(331)); -- 
    -- CP-element group 332:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 332: predecessors 
    -- CP-element group 332: 	327 
    -- CP-element group 332: successors 
    -- CP-element group 332: marked-successors 
    -- CP-element group 332: 	327 
    -- CP-element group 332: 	329 
    -- CP-element group 332:  members (3) 
      -- CP-element group 332: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_1064_request/ack
      -- CP-element group 332: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_1064_request/$exit
      -- CP-element group 332: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_1064_sample_completed_
      -- 
    ack_1808_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 332_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1064_final_reg_ack_0, ack => maxPool4_CP_346_elements(332)); -- 
    -- CP-element group 333:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 333: predecessors 
    -- CP-element group 333: 	328 
    -- CP-element group 333: successors 
    -- CP-element group 333: 	334 
    -- CP-element group 333: marked-successors 
    -- CP-element group 333: 	328 
    -- CP-element group 333:  members (3) 
      -- CP-element group 333: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_1064_complete/$exit
      -- CP-element group 333: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_1064_update_completed_
      -- CP-element group 333: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_1064_complete/ack
      -- 
    ack_1813_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 333_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1064_final_reg_ack_1, ack => maxPool4_CP_346_elements(333)); -- 
    -- CP-element group 334:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 334: predecessors 
    -- CP-element group 334: 	333 
    -- CP-element group 334: marked-predecessors 
    -- CP-element group 334: 	336 
    -- CP-element group 334: successors 
    -- CP-element group 334: 	336 
    -- CP-element group 334:  members (3) 
      -- CP-element group 334: 	 assign_stmt_97_to_assign_stmt_1138/assign_stmt_1068_sample_start_
      -- CP-element group 334: 	 assign_stmt_97_to_assign_stmt_1138/assign_stmt_1068_Sample/$entry
      -- CP-element group 334: 	 assign_stmt_97_to_assign_stmt_1138/assign_stmt_1068_Sample/req
      -- 
    req_1821_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1821_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(334), ack => W_myptr6_1063_delayed_8_0_1066_inst_req_0); -- 
    maxPool4_cp_element_group_334: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_334"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(333) & maxPool4_CP_346_elements(336);
      gj_maxPool4_cp_element_group_334 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(334), clk => clk, reset => reset); --
    end block;
    -- CP-element group 335:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 335: predecessors 
    -- CP-element group 335: marked-predecessors 
    -- CP-element group 335: 	337 
    -- CP-element group 335: 	344 
    -- CP-element group 335: successors 
    -- CP-element group 335: 	337 
    -- CP-element group 335:  members (3) 
      -- CP-element group 335: 	 assign_stmt_97_to_assign_stmt_1138/assign_stmt_1068_update_start_
      -- CP-element group 335: 	 assign_stmt_97_to_assign_stmt_1138/assign_stmt_1068_Update/req
      -- CP-element group 335: 	 assign_stmt_97_to_assign_stmt_1138/assign_stmt_1068_Update/$entry
      -- 
    req_1826_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1826_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(335), ack => W_myptr6_1063_delayed_8_0_1066_inst_req_1); -- 
    maxPool4_cp_element_group_335: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_335"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(337) & maxPool4_CP_346_elements(344);
      gj_maxPool4_cp_element_group_335 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(335), clk => clk, reset => reset); --
    end block;
    -- CP-element group 336:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 336: predecessors 
    -- CP-element group 336: 	334 
    -- CP-element group 336: successors 
    -- CP-element group 336: marked-successors 
    -- CP-element group 336: 	328 
    -- CP-element group 336: 	334 
    -- CP-element group 336:  members (3) 
      -- CP-element group 336: 	 assign_stmt_97_to_assign_stmt_1138/assign_stmt_1068_sample_completed_
      -- CP-element group 336: 	 assign_stmt_97_to_assign_stmt_1138/assign_stmt_1068_Sample/$exit
      -- CP-element group 336: 	 assign_stmt_97_to_assign_stmt_1138/assign_stmt_1068_Sample/ack
      -- 
    ack_1822_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 336_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_myptr6_1063_delayed_8_0_1066_inst_ack_0, ack => maxPool4_CP_346_elements(336)); -- 
    -- CP-element group 337:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 337: predecessors 
    -- CP-element group 337: 	335 
    -- CP-element group 337: successors 
    -- CP-element group 337: 	342 
    -- CP-element group 337: marked-successors 
    -- CP-element group 337: 	335 
    -- CP-element group 337:  members (19) 
      -- CP-element group 337: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1070_base_address_calculated
      -- CP-element group 337: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1070_base_addr_resize/$exit
      -- CP-element group 337: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1070_base_addr_resize/$entry
      -- CP-element group 337: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1070_word_address_calculated
      -- CP-element group 337: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1070_word_addrgen/$entry
      -- CP-element group 337: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1070_word_addrgen/$exit
      -- CP-element group 337: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1070_word_addrgen/root_register_req
      -- CP-element group 337: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1070_base_addr_resize/base_resize_ack
      -- CP-element group 337: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1070_root_address_calculated
      -- CP-element group 337: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1070_base_plus_offset/$entry
      -- CP-element group 337: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1070_base_plus_offset/$exit
      -- CP-element group 337: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1070_base_addr_resize/base_resize_req
      -- CP-element group 337: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1070_base_address_resized
      -- CP-element group 337: 	 assign_stmt_97_to_assign_stmt_1138/assign_stmt_1068_update_completed_
      -- CP-element group 337: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1070_word_addrgen/root_register_ack
      -- CP-element group 337: 	 assign_stmt_97_to_assign_stmt_1138/assign_stmt_1068_Update/ack
      -- CP-element group 337: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1070_base_plus_offset/sum_rename_ack
      -- CP-element group 337: 	 assign_stmt_97_to_assign_stmt_1138/assign_stmt_1068_Update/$exit
      -- CP-element group 337: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1070_base_plus_offset/sum_rename_req
      -- 
    ack_1827_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 337_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_myptr6_1063_delayed_8_0_1066_inst_ack_1, ack => maxPool4_CP_346_elements(337)); -- 
    -- CP-element group 338:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 338: predecessors 
    -- CP-element group 338: 	71 
    -- CP-element group 338: 	75 
    -- CP-element group 338: 	79 
    -- CP-element group 338: 	83 
    -- CP-element group 338: 	135 
    -- CP-element group 338: 	139 
    -- CP-element group 338: 	143 
    -- CP-element group 338: 	147 
    -- CP-element group 338: 	199 
    -- CP-element group 338: 	203 
    -- CP-element group 338: 	207 
    -- CP-element group 338: 	211 
    -- CP-element group 338: 	263 
    -- CP-element group 338: 	267 
    -- CP-element group 338: 	271 
    -- CP-element group 338: 	275 
    -- CP-element group 338: marked-predecessors 
    -- CP-element group 338: 	340 
    -- CP-element group 338: successors 
    -- CP-element group 338: 	340 
    -- CP-element group 338:  members (3) 
      -- CP-element group 338: 	 assign_stmt_97_to_assign_stmt_1138/CONCAT_u32_u64_1081_sample_start_
      -- CP-element group 338: 	 assign_stmt_97_to_assign_stmt_1138/CONCAT_u32_u64_1081_Sample/rr
      -- CP-element group 338: 	 assign_stmt_97_to_assign_stmt_1138/CONCAT_u32_u64_1081_Sample/$entry
      -- 
    rr_1835_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1835_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(338), ack => CONCAT_u32_u64_1081_inst_req_0); -- 
    maxPool4_cp_element_group_338: block -- 
      constant place_capacities: IntegerArray(0 to 16) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_markings: IntegerArray(0 to 16)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 1);
      constant place_delays: IntegerArray(0 to 16) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_338"; 
      signal preds: BooleanArray(1 to 17); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(71) & maxPool4_CP_346_elements(75) & maxPool4_CP_346_elements(79) & maxPool4_CP_346_elements(83) & maxPool4_CP_346_elements(135) & maxPool4_CP_346_elements(139) & maxPool4_CP_346_elements(143) & maxPool4_CP_346_elements(147) & maxPool4_CP_346_elements(199) & maxPool4_CP_346_elements(203) & maxPool4_CP_346_elements(207) & maxPool4_CP_346_elements(211) & maxPool4_CP_346_elements(263) & maxPool4_CP_346_elements(267) & maxPool4_CP_346_elements(271) & maxPool4_CP_346_elements(275) & maxPool4_CP_346_elements(340);
      gj_maxPool4_cp_element_group_338 : generic_join generic map(name => joinName, number_of_predecessors => 17, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(338), clk => clk, reset => reset); --
    end block;
    -- CP-element group 339:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 339: predecessors 
    -- CP-element group 339: marked-predecessors 
    -- CP-element group 339: 	341 
    -- CP-element group 339: 	344 
    -- CP-element group 339: successors 
    -- CP-element group 339: 	341 
    -- CP-element group 339:  members (3) 
      -- CP-element group 339: 	 assign_stmt_97_to_assign_stmt_1138/CONCAT_u32_u64_1081_update_start_
      -- CP-element group 339: 	 assign_stmt_97_to_assign_stmt_1138/CONCAT_u32_u64_1081_Update/cr
      -- CP-element group 339: 	 assign_stmt_97_to_assign_stmt_1138/CONCAT_u32_u64_1081_Update/$entry
      -- 
    cr_1840_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1840_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(339), ack => CONCAT_u32_u64_1081_inst_req_1); -- 
    maxPool4_cp_element_group_339: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_339"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(341) & maxPool4_CP_346_elements(344);
      gj_maxPool4_cp_element_group_339 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(339), clk => clk, reset => reset); --
    end block;
    -- CP-element group 340:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 340: predecessors 
    -- CP-element group 340: 	338 
    -- CP-element group 340: successors 
    -- CP-element group 340: marked-successors 
    -- CP-element group 340: 	69 
    -- CP-element group 340: 	73 
    -- CP-element group 340: 	77 
    -- CP-element group 340: 	81 
    -- CP-element group 340: 	133 
    -- CP-element group 340: 	137 
    -- CP-element group 340: 	141 
    -- CP-element group 340: 	145 
    -- CP-element group 340: 	197 
    -- CP-element group 340: 	201 
    -- CP-element group 340: 	205 
    -- CP-element group 340: 	209 
    -- CP-element group 340: 	261 
    -- CP-element group 340: 	265 
    -- CP-element group 340: 	269 
    -- CP-element group 340: 	273 
    -- CP-element group 340: 	338 
    -- CP-element group 340:  members (3) 
      -- CP-element group 340: 	 assign_stmt_97_to_assign_stmt_1138/CONCAT_u32_u64_1081_sample_completed_
      -- CP-element group 340: 	 assign_stmt_97_to_assign_stmt_1138/CONCAT_u32_u64_1081_Sample/ra
      -- CP-element group 340: 	 assign_stmt_97_to_assign_stmt_1138/CONCAT_u32_u64_1081_Sample/$exit
      -- 
    ra_1836_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 340_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u32_u64_1081_inst_ack_0, ack => maxPool4_CP_346_elements(340)); -- 
    -- CP-element group 341:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 341: predecessors 
    -- CP-element group 341: 	339 
    -- CP-element group 341: successors 
    -- CP-element group 341: 	342 
    -- CP-element group 341: marked-successors 
    -- CP-element group 341: 	339 
    -- CP-element group 341:  members (3) 
      -- CP-element group 341: 	 assign_stmt_97_to_assign_stmt_1138/CONCAT_u32_u64_1081_update_completed_
      -- CP-element group 341: 	 assign_stmt_97_to_assign_stmt_1138/CONCAT_u32_u64_1081_Update/ca
      -- CP-element group 341: 	 assign_stmt_97_to_assign_stmt_1138/CONCAT_u32_u64_1081_Update/$exit
      -- 
    ca_1841_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 341_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u32_u64_1081_inst_ack_1, ack => maxPool4_CP_346_elements(341)); -- 
    -- CP-element group 342:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 342: predecessors 
    -- CP-element group 342: 	337 
    -- CP-element group 342: 	341 
    -- CP-element group 342: 	388 
    -- CP-element group 342: marked-predecessors 
    -- CP-element group 342: 	344 
    -- CP-element group 342: successors 
    -- CP-element group 342: 	344 
    -- CP-element group 342:  members (9) 
      -- CP-element group 342: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1070_Sample/ptr_deref_1070_Split/split_req
      -- CP-element group 342: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1070_Sample/ptr_deref_1070_Split/$exit
      -- CP-element group 342: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1070_Sample/ptr_deref_1070_Split/$entry
      -- CP-element group 342: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1070_Sample/word_access_start/word_0/rr
      -- CP-element group 342: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1070_Sample/word_access_start/word_0/$entry
      -- CP-element group 342: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1070_Sample/$entry
      -- CP-element group 342: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1070_sample_start_
      -- CP-element group 342: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1070_Sample/word_access_start/$entry
      -- CP-element group 342: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1070_Sample/ptr_deref_1070_Split/split_ack
      -- 
    rr_1879_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1879_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(342), ack => ptr_deref_1070_store_0_req_0); -- 
    maxPool4_cp_element_group_342: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_342"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(337) & maxPool4_CP_346_elements(341) & maxPool4_CP_346_elements(388) & maxPool4_CP_346_elements(344);
      gj_maxPool4_cp_element_group_342 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(342), clk => clk, reset => reset); --
    end block;
    -- CP-element group 343:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 343: predecessors 
    -- CP-element group 343: marked-predecessors 
    -- CP-element group 343: 	345 
    -- CP-element group 343: successors 
    -- CP-element group 343: 	345 
    -- CP-element group 343:  members (5) 
      -- CP-element group 343: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1070_Update/word_access_complete/word_0/$entry
      -- CP-element group 343: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1070_Update/word_access_complete/word_0/cr
      -- CP-element group 343: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1070_Update/$entry
      -- CP-element group 343: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1070_update_start_
      -- CP-element group 343: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1070_Update/word_access_complete/$entry
      -- 
    cr_1890_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1890_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(343), ack => ptr_deref_1070_store_0_req_1); -- 
    maxPool4_cp_element_group_343: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_343"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= maxPool4_CP_346_elements(345);
      gj_maxPool4_cp_element_group_343 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(343), clk => clk, reset => reset); --
    end block;
    -- CP-element group 344:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 344: predecessors 
    -- CP-element group 344: 	342 
    -- CP-element group 344: successors 
    -- CP-element group 344: 	389 
    -- CP-element group 344: marked-successors 
    -- CP-element group 344: 	335 
    -- CP-element group 344: 	339 
    -- CP-element group 344: 	342 
    -- CP-element group 344:  members (5) 
      -- CP-element group 344: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1070_Sample/word_access_start/word_0/ra
      -- CP-element group 344: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1070_Sample/$exit
      -- CP-element group 344: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1070_sample_completed_
      -- CP-element group 344: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1070_Sample/word_access_start/$exit
      -- CP-element group 344: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1070_Sample/word_access_start/word_0/$exit
      -- 
    ra_1880_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 344_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1070_store_0_ack_0, ack => maxPool4_CP_346_elements(344)); -- 
    -- CP-element group 345:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 345: predecessors 
    -- CP-element group 345: 	343 
    -- CP-element group 345: successors 
    -- CP-element group 345: 	391 
    -- CP-element group 345: marked-successors 
    -- CP-element group 345: 	343 
    -- CP-element group 345:  members (5) 
      -- CP-element group 345: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1070_Update/word_access_complete/$exit
      -- CP-element group 345: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1070_Update/word_access_complete/word_0/$exit
      -- CP-element group 345: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1070_Update/word_access_complete/word_0/ca
      -- CP-element group 345: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1070_Update/$exit
      -- CP-element group 345: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1070_update_completed_
      -- 
    ca_1891_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 345_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1070_store_0_ack_1, ack => maxPool4_CP_346_elements(345)); -- 
    -- CP-element group 346:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 346: predecessors 
    -- CP-element group 346: 	350 
    -- CP-element group 346: marked-predecessors 
    -- CP-element group 346: 	351 
    -- CP-element group 346: successors 
    -- CP-element group 346: 	351 
    -- CP-element group 346:  members (3) 
      -- CP-element group 346: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_1090_sample_start_
      -- CP-element group 346: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_1090_request/$entry
      -- CP-element group 346: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_1090_request/req
      -- 
    req_1931_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1931_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(346), ack => addr_of_1090_final_reg_req_0); -- 
    maxPool4_cp_element_group_346: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_346"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(350) & maxPool4_CP_346_elements(351);
      gj_maxPool4_cp_element_group_346 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(346), clk => clk, reset => reset); --
    end block;
    -- CP-element group 347:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 347: predecessors 
    -- CP-element group 347: 	1 
    -- CP-element group 347: marked-predecessors 
    -- CP-element group 347: 	352 
    -- CP-element group 347: 	355 
    -- CP-element group 347: successors 
    -- CP-element group 347: 	352 
    -- CP-element group 347:  members (3) 
      -- CP-element group 347: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_1090_update_start_
      -- CP-element group 347: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_1090_complete/$entry
      -- CP-element group 347: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_1090_complete/req
      -- 
    req_1936_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1936_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(347), ack => addr_of_1090_final_reg_req_1); -- 
    maxPool4_cp_element_group_347: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_347"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(1) & maxPool4_CP_346_elements(352) & maxPool4_CP_346_elements(355);
      gj_maxPool4_cp_element_group_347 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(347), clk => clk, reset => reset); --
    end block;
    -- CP-element group 348:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 348: predecessors 
    -- CP-element group 348: 	1 
    -- CP-element group 348: marked-predecessors 
    -- CP-element group 348: 	350 
    -- CP-element group 348: 	351 
    -- CP-element group 348: successors 
    -- CP-element group 348: 	350 
    -- CP-element group 348:  members (3) 
      -- CP-element group 348: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1089_final_index_sum_regn_update_start
      -- CP-element group 348: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1089_final_index_sum_regn_Update/$entry
      -- CP-element group 348: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1089_final_index_sum_regn_Update/req
      -- 
    req_1921_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1921_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(348), ack => array_obj_ref_1089_index_offset_req_1); -- 
    maxPool4_cp_element_group_348: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_348"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(1) & maxPool4_CP_346_elements(350) & maxPool4_CP_346_elements(351);
      gj_maxPool4_cp_element_group_348 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(348), clk => clk, reset => reset); --
    end block;
    -- CP-element group 349:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 349: predecessors 
    -- CP-element group 349: 	1 
    -- CP-element group 349: successors 
    -- CP-element group 349: 	391 
    -- CP-element group 349: marked-successors 
    -- CP-element group 349: 	2 
    -- CP-element group 349:  members (3) 
      -- CP-element group 349: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1089_final_index_sum_regn_sample_complete
      -- CP-element group 349: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1089_final_index_sum_regn_Sample/$exit
      -- CP-element group 349: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1089_final_index_sum_regn_Sample/ack
      -- 
    ack_1917_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 349_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1089_index_offset_ack_0, ack => maxPool4_CP_346_elements(349)); -- 
    -- CP-element group 350:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 350: predecessors 
    -- CP-element group 350: 	348 
    -- CP-element group 350: successors 
    -- CP-element group 350: 	346 
    -- CP-element group 350: marked-successors 
    -- CP-element group 350: 	348 
    -- CP-element group 350:  members (8) 
      -- CP-element group 350: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1089_root_address_calculated
      -- CP-element group 350: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1089_offset_calculated
      -- CP-element group 350: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1089_final_index_sum_regn_Update/$exit
      -- CP-element group 350: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1089_final_index_sum_regn_Update/ack
      -- CP-element group 350: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1089_base_plus_offset/$entry
      -- CP-element group 350: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1089_base_plus_offset/$exit
      -- CP-element group 350: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1089_base_plus_offset/sum_rename_req
      -- CP-element group 350: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1089_base_plus_offset/sum_rename_ack
      -- 
    ack_1922_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 350_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1089_index_offset_ack_1, ack => maxPool4_CP_346_elements(350)); -- 
    -- CP-element group 351:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 351: predecessors 
    -- CP-element group 351: 	346 
    -- CP-element group 351: successors 
    -- CP-element group 351: marked-successors 
    -- CP-element group 351: 	346 
    -- CP-element group 351: 	348 
    -- CP-element group 351:  members (3) 
      -- CP-element group 351: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_1090_sample_completed_
      -- CP-element group 351: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_1090_request/$exit
      -- CP-element group 351: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_1090_request/ack
      -- 
    ack_1932_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 351_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1090_final_reg_ack_0, ack => maxPool4_CP_346_elements(351)); -- 
    -- CP-element group 352:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 352: predecessors 
    -- CP-element group 352: 	347 
    -- CP-element group 352: successors 
    -- CP-element group 352: 	353 
    -- CP-element group 352: marked-successors 
    -- CP-element group 352: 	347 
    -- CP-element group 352:  members (3) 
      -- CP-element group 352: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_1090_update_completed_
      -- CP-element group 352: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_1090_complete/$exit
      -- CP-element group 352: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_1090_complete/ack
      -- 
    ack_1937_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 352_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1090_final_reg_ack_1, ack => maxPool4_CP_346_elements(352)); -- 
    -- CP-element group 353:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 353: predecessors 
    -- CP-element group 353: 	352 
    -- CP-element group 353: marked-predecessors 
    -- CP-element group 353: 	355 
    -- CP-element group 353: successors 
    -- CP-element group 353: 	355 
    -- CP-element group 353:  members (3) 
      -- CP-element group 353: 	 assign_stmt_97_to_assign_stmt_1138/assign_stmt_1094_sample_start_
      -- CP-element group 353: 	 assign_stmt_97_to_assign_stmt_1138/assign_stmt_1094_Sample/$entry
      -- CP-element group 353: 	 assign_stmt_97_to_assign_stmt_1138/assign_stmt_1094_Sample/req
      -- 
    req_1945_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1945_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(353), ack => W_myptr7_1086_delayed_8_0_1092_inst_req_0); -- 
    maxPool4_cp_element_group_353: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_353"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(352) & maxPool4_CP_346_elements(355);
      gj_maxPool4_cp_element_group_353 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(353), clk => clk, reset => reset); --
    end block;
    -- CP-element group 354:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 354: predecessors 
    -- CP-element group 354: marked-predecessors 
    -- CP-element group 354: 	356 
    -- CP-element group 354: 	363 
    -- CP-element group 354: successors 
    -- CP-element group 354: 	356 
    -- CP-element group 354:  members (3) 
      -- CP-element group 354: 	 assign_stmt_97_to_assign_stmt_1138/assign_stmt_1094_update_start_
      -- CP-element group 354: 	 assign_stmt_97_to_assign_stmt_1138/assign_stmt_1094_Update/$entry
      -- CP-element group 354: 	 assign_stmt_97_to_assign_stmt_1138/assign_stmt_1094_Update/req
      -- 
    req_1950_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1950_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(354), ack => W_myptr7_1086_delayed_8_0_1092_inst_req_1); -- 
    maxPool4_cp_element_group_354: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_354"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(356) & maxPool4_CP_346_elements(363);
      gj_maxPool4_cp_element_group_354 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(354), clk => clk, reset => reset); --
    end block;
    -- CP-element group 355:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 355: predecessors 
    -- CP-element group 355: 	353 
    -- CP-element group 355: successors 
    -- CP-element group 355: marked-successors 
    -- CP-element group 355: 	347 
    -- CP-element group 355: 	353 
    -- CP-element group 355:  members (3) 
      -- CP-element group 355: 	 assign_stmt_97_to_assign_stmt_1138/assign_stmt_1094_sample_completed_
      -- CP-element group 355: 	 assign_stmt_97_to_assign_stmt_1138/assign_stmt_1094_Sample/$exit
      -- CP-element group 355: 	 assign_stmt_97_to_assign_stmt_1138/assign_stmt_1094_Sample/ack
      -- 
    ack_1946_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 355_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_myptr7_1086_delayed_8_0_1092_inst_ack_0, ack => maxPool4_CP_346_elements(355)); -- 
    -- CP-element group 356:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 356: predecessors 
    -- CP-element group 356: 	354 
    -- CP-element group 356: successors 
    -- CP-element group 356: 	361 
    -- CP-element group 356: marked-successors 
    -- CP-element group 356: 	354 
    -- CP-element group 356:  members (19) 
      -- CP-element group 356: 	 assign_stmt_97_to_assign_stmt_1138/assign_stmt_1094_update_completed_
      -- CP-element group 356: 	 assign_stmt_97_to_assign_stmt_1138/assign_stmt_1094_Update/$exit
      -- CP-element group 356: 	 assign_stmt_97_to_assign_stmt_1138/assign_stmt_1094_Update/ack
      -- CP-element group 356: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1096_base_address_calculated
      -- CP-element group 356: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1096_word_address_calculated
      -- CP-element group 356: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1096_root_address_calculated
      -- CP-element group 356: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1096_base_address_resized
      -- CP-element group 356: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1096_base_addr_resize/$entry
      -- CP-element group 356: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1096_base_addr_resize/$exit
      -- CP-element group 356: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1096_base_addr_resize/base_resize_req
      -- CP-element group 356: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1096_base_addr_resize/base_resize_ack
      -- CP-element group 356: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1096_base_plus_offset/$entry
      -- CP-element group 356: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1096_base_plus_offset/$exit
      -- CP-element group 356: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1096_base_plus_offset/sum_rename_req
      -- CP-element group 356: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1096_base_plus_offset/sum_rename_ack
      -- CP-element group 356: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1096_word_addrgen/$entry
      -- CP-element group 356: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1096_word_addrgen/$exit
      -- CP-element group 356: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1096_word_addrgen/root_register_req
      -- CP-element group 356: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1096_word_addrgen/root_register_ack
      -- 
    ack_1951_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 356_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_myptr7_1086_delayed_8_0_1092_inst_ack_1, ack => maxPool4_CP_346_elements(356)); -- 
    -- CP-element group 357:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 357: predecessors 
    -- CP-element group 357: 	87 
    -- CP-element group 357: 	91 
    -- CP-element group 357: 	95 
    -- CP-element group 357: 	99 
    -- CP-element group 357: 	151 
    -- CP-element group 357: 	155 
    -- CP-element group 357: 	159 
    -- CP-element group 357: 	163 
    -- CP-element group 357: 	215 
    -- CP-element group 357: 	219 
    -- CP-element group 357: 	223 
    -- CP-element group 357: 	227 
    -- CP-element group 357: 	279 
    -- CP-element group 357: 	283 
    -- CP-element group 357: 	287 
    -- CP-element group 357: 	291 
    -- CP-element group 357: marked-predecessors 
    -- CP-element group 357: 	359 
    -- CP-element group 357: successors 
    -- CP-element group 357: 	359 
    -- CP-element group 357:  members (3) 
      -- CP-element group 357: 	 assign_stmt_97_to_assign_stmt_1138/CONCAT_u32_u64_1107_sample_start_
      -- CP-element group 357: 	 assign_stmt_97_to_assign_stmt_1138/CONCAT_u32_u64_1107_Sample/$entry
      -- CP-element group 357: 	 assign_stmt_97_to_assign_stmt_1138/CONCAT_u32_u64_1107_Sample/rr
      -- 
    rr_1959_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1959_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(357), ack => CONCAT_u32_u64_1107_inst_req_0); -- 
    maxPool4_cp_element_group_357: block -- 
      constant place_capacities: IntegerArray(0 to 16) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_markings: IntegerArray(0 to 16)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 1);
      constant place_delays: IntegerArray(0 to 16) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_357"; 
      signal preds: BooleanArray(1 to 17); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(87) & maxPool4_CP_346_elements(91) & maxPool4_CP_346_elements(95) & maxPool4_CP_346_elements(99) & maxPool4_CP_346_elements(151) & maxPool4_CP_346_elements(155) & maxPool4_CP_346_elements(159) & maxPool4_CP_346_elements(163) & maxPool4_CP_346_elements(215) & maxPool4_CP_346_elements(219) & maxPool4_CP_346_elements(223) & maxPool4_CP_346_elements(227) & maxPool4_CP_346_elements(279) & maxPool4_CP_346_elements(283) & maxPool4_CP_346_elements(287) & maxPool4_CP_346_elements(291) & maxPool4_CP_346_elements(359);
      gj_maxPool4_cp_element_group_357 : generic_join generic map(name => joinName, number_of_predecessors => 17, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(357), clk => clk, reset => reset); --
    end block;
    -- CP-element group 358:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 358: predecessors 
    -- CP-element group 358: marked-predecessors 
    -- CP-element group 358: 	360 
    -- CP-element group 358: 	363 
    -- CP-element group 358: successors 
    -- CP-element group 358: 	360 
    -- CP-element group 358:  members (3) 
      -- CP-element group 358: 	 assign_stmt_97_to_assign_stmt_1138/CONCAT_u32_u64_1107_update_start_
      -- CP-element group 358: 	 assign_stmt_97_to_assign_stmt_1138/CONCAT_u32_u64_1107_Update/$entry
      -- CP-element group 358: 	 assign_stmt_97_to_assign_stmt_1138/CONCAT_u32_u64_1107_Update/cr
      -- 
    cr_1964_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1964_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(358), ack => CONCAT_u32_u64_1107_inst_req_1); -- 
    maxPool4_cp_element_group_358: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_358"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(360) & maxPool4_CP_346_elements(363);
      gj_maxPool4_cp_element_group_358 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(358), clk => clk, reset => reset); --
    end block;
    -- CP-element group 359:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 359: predecessors 
    -- CP-element group 359: 	357 
    -- CP-element group 359: successors 
    -- CP-element group 359: marked-successors 
    -- CP-element group 359: 	85 
    -- CP-element group 359: 	89 
    -- CP-element group 359: 	93 
    -- CP-element group 359: 	97 
    -- CP-element group 359: 	149 
    -- CP-element group 359: 	153 
    -- CP-element group 359: 	157 
    -- CP-element group 359: 	161 
    -- CP-element group 359: 	213 
    -- CP-element group 359: 	217 
    -- CP-element group 359: 	221 
    -- CP-element group 359: 	225 
    -- CP-element group 359: 	277 
    -- CP-element group 359: 	281 
    -- CP-element group 359: 	285 
    -- CP-element group 359: 	289 
    -- CP-element group 359: 	357 
    -- CP-element group 359:  members (3) 
      -- CP-element group 359: 	 assign_stmt_97_to_assign_stmt_1138/CONCAT_u32_u64_1107_sample_completed_
      -- CP-element group 359: 	 assign_stmt_97_to_assign_stmt_1138/CONCAT_u32_u64_1107_Sample/$exit
      -- CP-element group 359: 	 assign_stmt_97_to_assign_stmt_1138/CONCAT_u32_u64_1107_Sample/ra
      -- 
    ra_1960_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 359_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u32_u64_1107_inst_ack_0, ack => maxPool4_CP_346_elements(359)); -- 
    -- CP-element group 360:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 360: predecessors 
    -- CP-element group 360: 	358 
    -- CP-element group 360: successors 
    -- CP-element group 360: 	361 
    -- CP-element group 360: marked-successors 
    -- CP-element group 360: 	358 
    -- CP-element group 360:  members (3) 
      -- CP-element group 360: 	 assign_stmt_97_to_assign_stmt_1138/CONCAT_u32_u64_1107_update_completed_
      -- CP-element group 360: 	 assign_stmt_97_to_assign_stmt_1138/CONCAT_u32_u64_1107_Update/$exit
      -- CP-element group 360: 	 assign_stmt_97_to_assign_stmt_1138/CONCAT_u32_u64_1107_Update/ca
      -- 
    ca_1965_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 360_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u32_u64_1107_inst_ack_1, ack => maxPool4_CP_346_elements(360)); -- 
    -- CP-element group 361:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 361: predecessors 
    -- CP-element group 361: 	356 
    -- CP-element group 361: 	360 
    -- CP-element group 361: 	389 
    -- CP-element group 361: marked-predecessors 
    -- CP-element group 361: 	363 
    -- CP-element group 361: successors 
    -- CP-element group 361: 	363 
    -- CP-element group 361:  members (9) 
      -- CP-element group 361: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1096_sample_start_
      -- CP-element group 361: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1096_Sample/$entry
      -- CP-element group 361: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1096_Sample/ptr_deref_1096_Split/$entry
      -- CP-element group 361: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1096_Sample/ptr_deref_1096_Split/$exit
      -- CP-element group 361: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1096_Sample/ptr_deref_1096_Split/split_req
      -- CP-element group 361: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1096_Sample/ptr_deref_1096_Split/split_ack
      -- CP-element group 361: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1096_Sample/word_access_start/$entry
      -- CP-element group 361: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1096_Sample/word_access_start/word_0/$entry
      -- CP-element group 361: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1096_Sample/word_access_start/word_0/rr
      -- 
    rr_2003_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2003_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(361), ack => ptr_deref_1096_store_0_req_0); -- 
    maxPool4_cp_element_group_361: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_361"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(356) & maxPool4_CP_346_elements(360) & maxPool4_CP_346_elements(389) & maxPool4_CP_346_elements(363);
      gj_maxPool4_cp_element_group_361 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(361), clk => clk, reset => reset); --
    end block;
    -- CP-element group 362:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 362: predecessors 
    -- CP-element group 362: marked-predecessors 
    -- CP-element group 362: 	364 
    -- CP-element group 362: successors 
    -- CP-element group 362: 	364 
    -- CP-element group 362:  members (5) 
      -- CP-element group 362: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1096_update_start_
      -- CP-element group 362: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1096_Update/$entry
      -- CP-element group 362: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1096_Update/word_access_complete/$entry
      -- CP-element group 362: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1096_Update/word_access_complete/word_0/$entry
      -- CP-element group 362: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1096_Update/word_access_complete/word_0/cr
      -- 
    cr_2014_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2014_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(362), ack => ptr_deref_1096_store_0_req_1); -- 
    maxPool4_cp_element_group_362: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_362"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= maxPool4_CP_346_elements(364);
      gj_maxPool4_cp_element_group_362 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(362), clk => clk, reset => reset); --
    end block;
    -- CP-element group 363:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 363: predecessors 
    -- CP-element group 363: 	361 
    -- CP-element group 363: successors 
    -- CP-element group 363: 	390 
    -- CP-element group 363: marked-successors 
    -- CP-element group 363: 	354 
    -- CP-element group 363: 	358 
    -- CP-element group 363: 	361 
    -- CP-element group 363:  members (5) 
      -- CP-element group 363: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1096_sample_completed_
      -- CP-element group 363: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1096_Sample/$exit
      -- CP-element group 363: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1096_Sample/word_access_start/$exit
      -- CP-element group 363: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1096_Sample/word_access_start/word_0/$exit
      -- CP-element group 363: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1096_Sample/word_access_start/word_0/ra
      -- 
    ra_2004_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 363_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1096_store_0_ack_0, ack => maxPool4_CP_346_elements(363)); -- 
    -- CP-element group 364:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 364: predecessors 
    -- CP-element group 364: 	362 
    -- CP-element group 364: successors 
    -- CP-element group 364: 	391 
    -- CP-element group 364: marked-successors 
    -- CP-element group 364: 	362 
    -- CP-element group 364:  members (5) 
      -- CP-element group 364: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1096_update_completed_
      -- CP-element group 364: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1096_Update/$exit
      -- CP-element group 364: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1096_Update/word_access_complete/$exit
      -- CP-element group 364: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1096_Update/word_access_complete/word_0/$exit
      -- CP-element group 364: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1096_Update/word_access_complete/word_0/ca
      -- 
    ca_2015_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 364_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1096_store_0_ack_1, ack => maxPool4_CP_346_elements(364)); -- 
    -- CP-element group 365:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 365: predecessors 
    -- CP-element group 365: 	369 
    -- CP-element group 365: marked-predecessors 
    -- CP-element group 365: 	370 
    -- CP-element group 365: successors 
    -- CP-element group 365: 	370 
    -- CP-element group 365:  members (3) 
      -- CP-element group 365: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_1116_sample_start_
      -- CP-element group 365: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_1116_request/$entry
      -- CP-element group 365: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_1116_request/req
      -- 
    req_2055_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2055_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(365), ack => addr_of_1116_final_reg_req_0); -- 
    maxPool4_cp_element_group_365: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_365"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(369) & maxPool4_CP_346_elements(370);
      gj_maxPool4_cp_element_group_365 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(365), clk => clk, reset => reset); --
    end block;
    -- CP-element group 366:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 366: predecessors 
    -- CP-element group 366: 	1 
    -- CP-element group 366: marked-predecessors 
    -- CP-element group 366: 	371 
    -- CP-element group 366: 	374 
    -- CP-element group 366: successors 
    -- CP-element group 366: 	371 
    -- CP-element group 366:  members (3) 
      -- CP-element group 366: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_1116_update_start_
      -- CP-element group 366: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_1116_complete/$entry
      -- CP-element group 366: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_1116_complete/req
      -- 
    req_2060_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2060_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(366), ack => addr_of_1116_final_reg_req_1); -- 
    maxPool4_cp_element_group_366: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_366"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(1) & maxPool4_CP_346_elements(371) & maxPool4_CP_346_elements(374);
      gj_maxPool4_cp_element_group_366 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(366), clk => clk, reset => reset); --
    end block;
    -- CP-element group 367:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 367: predecessors 
    -- CP-element group 367: 	1 
    -- CP-element group 367: marked-predecessors 
    -- CP-element group 367: 	369 
    -- CP-element group 367: 	370 
    -- CP-element group 367: successors 
    -- CP-element group 367: 	369 
    -- CP-element group 367:  members (3) 
      -- CP-element group 367: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1115_final_index_sum_regn_update_start
      -- CP-element group 367: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1115_final_index_sum_regn_Update/$entry
      -- CP-element group 367: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1115_final_index_sum_regn_Update/req
      -- 
    req_2045_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2045_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(367), ack => array_obj_ref_1115_index_offset_req_1); -- 
    maxPool4_cp_element_group_367: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_367"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(1) & maxPool4_CP_346_elements(369) & maxPool4_CP_346_elements(370);
      gj_maxPool4_cp_element_group_367 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(367), clk => clk, reset => reset); --
    end block;
    -- CP-element group 368:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 368: predecessors 
    -- CP-element group 368: 	1 
    -- CP-element group 368: successors 
    -- CP-element group 368: 	391 
    -- CP-element group 368: marked-successors 
    -- CP-element group 368: 	2 
    -- CP-element group 368:  members (3) 
      -- CP-element group 368: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1115_final_index_sum_regn_sample_complete
      -- CP-element group 368: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1115_final_index_sum_regn_Sample/$exit
      -- CP-element group 368: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1115_final_index_sum_regn_Sample/ack
      -- 
    ack_2041_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 368_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1115_index_offset_ack_0, ack => maxPool4_CP_346_elements(368)); -- 
    -- CP-element group 369:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 369: predecessors 
    -- CP-element group 369: 	367 
    -- CP-element group 369: successors 
    -- CP-element group 369: 	365 
    -- CP-element group 369: marked-successors 
    -- CP-element group 369: 	367 
    -- CP-element group 369:  members (8) 
      -- CP-element group 369: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1115_root_address_calculated
      -- CP-element group 369: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1115_offset_calculated
      -- CP-element group 369: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1115_final_index_sum_regn_Update/$exit
      -- CP-element group 369: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1115_final_index_sum_regn_Update/ack
      -- CP-element group 369: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1115_base_plus_offset/$entry
      -- CP-element group 369: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1115_base_plus_offset/$exit
      -- CP-element group 369: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1115_base_plus_offset/sum_rename_req
      -- CP-element group 369: 	 assign_stmt_97_to_assign_stmt_1138/array_obj_ref_1115_base_plus_offset/sum_rename_ack
      -- 
    ack_2046_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 369_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1115_index_offset_ack_1, ack => maxPool4_CP_346_elements(369)); -- 
    -- CP-element group 370:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 370: predecessors 
    -- CP-element group 370: 	365 
    -- CP-element group 370: successors 
    -- CP-element group 370: marked-successors 
    -- CP-element group 370: 	365 
    -- CP-element group 370: 	367 
    -- CP-element group 370:  members (3) 
      -- CP-element group 370: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_1116_sample_completed_
      -- CP-element group 370: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_1116_request/$exit
      -- CP-element group 370: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_1116_request/ack
      -- 
    ack_2056_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 370_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1116_final_reg_ack_0, ack => maxPool4_CP_346_elements(370)); -- 
    -- CP-element group 371:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 371: predecessors 
    -- CP-element group 371: 	366 
    -- CP-element group 371: successors 
    -- CP-element group 371: 	372 
    -- CP-element group 371: marked-successors 
    -- CP-element group 371: 	366 
    -- CP-element group 371:  members (3) 
      -- CP-element group 371: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_1116_update_completed_
      -- CP-element group 371: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_1116_complete/$exit
      -- CP-element group 371: 	 assign_stmt_97_to_assign_stmt_1138/addr_of_1116_complete/ack
      -- 
    ack_2061_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 371_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1116_final_reg_ack_1, ack => maxPool4_CP_346_elements(371)); -- 
    -- CP-element group 372:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 372: predecessors 
    -- CP-element group 372: 	371 
    -- CP-element group 372: marked-predecessors 
    -- CP-element group 372: 	374 
    -- CP-element group 372: successors 
    -- CP-element group 372: 	374 
    -- CP-element group 372:  members (3) 
      -- CP-element group 372: 	 assign_stmt_97_to_assign_stmt_1138/assign_stmt_1120_sample_start_
      -- CP-element group 372: 	 assign_stmt_97_to_assign_stmt_1138/assign_stmt_1120_Sample/$entry
      -- CP-element group 372: 	 assign_stmt_97_to_assign_stmt_1138/assign_stmt_1120_Sample/req
      -- 
    req_2069_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2069_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(372), ack => W_myptr8_1109_delayed_8_0_1118_inst_req_0); -- 
    maxPool4_cp_element_group_372: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_372"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(371) & maxPool4_CP_346_elements(374);
      gj_maxPool4_cp_element_group_372 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(372), clk => clk, reset => reset); --
    end block;
    -- CP-element group 373:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 373: predecessors 
    -- CP-element group 373: marked-predecessors 
    -- CP-element group 373: 	375 
    -- CP-element group 373: 	382 
    -- CP-element group 373: successors 
    -- CP-element group 373: 	375 
    -- CP-element group 373:  members (3) 
      -- CP-element group 373: 	 assign_stmt_97_to_assign_stmt_1138/assign_stmt_1120_update_start_
      -- CP-element group 373: 	 assign_stmt_97_to_assign_stmt_1138/assign_stmt_1120_Update/$entry
      -- CP-element group 373: 	 assign_stmt_97_to_assign_stmt_1138/assign_stmt_1120_Update/req
      -- 
    req_2074_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2074_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(373), ack => W_myptr8_1109_delayed_8_0_1118_inst_req_1); -- 
    maxPool4_cp_element_group_373: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_373"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(375) & maxPool4_CP_346_elements(382);
      gj_maxPool4_cp_element_group_373 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(373), clk => clk, reset => reset); --
    end block;
    -- CP-element group 374:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 374: predecessors 
    -- CP-element group 374: 	372 
    -- CP-element group 374: successors 
    -- CP-element group 374: marked-successors 
    -- CP-element group 374: 	366 
    -- CP-element group 374: 	372 
    -- CP-element group 374:  members (3) 
      -- CP-element group 374: 	 assign_stmt_97_to_assign_stmt_1138/assign_stmt_1120_sample_completed_
      -- CP-element group 374: 	 assign_stmt_97_to_assign_stmt_1138/assign_stmt_1120_Sample/$exit
      -- CP-element group 374: 	 assign_stmt_97_to_assign_stmt_1138/assign_stmt_1120_Sample/ack
      -- 
    ack_2070_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 374_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_myptr8_1109_delayed_8_0_1118_inst_ack_0, ack => maxPool4_CP_346_elements(374)); -- 
    -- CP-element group 375:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 375: predecessors 
    -- CP-element group 375: 	373 
    -- CP-element group 375: successors 
    -- CP-element group 375: 	380 
    -- CP-element group 375: marked-successors 
    -- CP-element group 375: 	373 
    -- CP-element group 375:  members (19) 
      -- CP-element group 375: 	 assign_stmt_97_to_assign_stmt_1138/assign_stmt_1120_update_completed_
      -- CP-element group 375: 	 assign_stmt_97_to_assign_stmt_1138/assign_stmt_1120_Update/$exit
      -- CP-element group 375: 	 assign_stmt_97_to_assign_stmt_1138/assign_stmt_1120_Update/ack
      -- CP-element group 375: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1122_base_address_calculated
      -- CP-element group 375: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1122_word_address_calculated
      -- CP-element group 375: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1122_root_address_calculated
      -- CP-element group 375: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1122_base_address_resized
      -- CP-element group 375: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1122_base_addr_resize/$entry
      -- CP-element group 375: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1122_base_addr_resize/$exit
      -- CP-element group 375: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1122_base_addr_resize/base_resize_req
      -- CP-element group 375: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1122_base_addr_resize/base_resize_ack
      -- CP-element group 375: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1122_base_plus_offset/$entry
      -- CP-element group 375: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1122_base_plus_offset/$exit
      -- CP-element group 375: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1122_base_plus_offset/sum_rename_req
      -- CP-element group 375: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1122_base_plus_offset/sum_rename_ack
      -- CP-element group 375: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1122_word_addrgen/$entry
      -- CP-element group 375: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1122_word_addrgen/$exit
      -- CP-element group 375: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1122_word_addrgen/root_register_req
      -- CP-element group 375: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1122_word_addrgen/root_register_ack
      -- 
    ack_2075_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 375_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_myptr8_1109_delayed_8_0_1118_inst_ack_1, ack => maxPool4_CP_346_elements(375)); -- 
    -- CP-element group 376:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 376: predecessors 
    -- CP-element group 376: 	103 
    -- CP-element group 376: 	107 
    -- CP-element group 376: 	111 
    -- CP-element group 376: 	115 
    -- CP-element group 376: 	167 
    -- CP-element group 376: 	171 
    -- CP-element group 376: 	175 
    -- CP-element group 376: 	179 
    -- CP-element group 376: 	231 
    -- CP-element group 376: 	235 
    -- CP-element group 376: 	239 
    -- CP-element group 376: 	243 
    -- CP-element group 376: 	295 
    -- CP-element group 376: 	299 
    -- CP-element group 376: 	303 
    -- CP-element group 376: 	307 
    -- CP-element group 376: marked-predecessors 
    -- CP-element group 376: 	378 
    -- CP-element group 376: successors 
    -- CP-element group 376: 	378 
    -- CP-element group 376:  members (3) 
      -- CP-element group 376: 	 assign_stmt_97_to_assign_stmt_1138/CONCAT_u32_u64_1133_sample_start_
      -- CP-element group 376: 	 assign_stmt_97_to_assign_stmt_1138/CONCAT_u32_u64_1133_Sample/$entry
      -- CP-element group 376: 	 assign_stmt_97_to_assign_stmt_1138/CONCAT_u32_u64_1133_Sample/rr
      -- 
    rr_2083_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2083_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(376), ack => CONCAT_u32_u64_1133_inst_req_0); -- 
    maxPool4_cp_element_group_376: block -- 
      constant place_capacities: IntegerArray(0 to 16) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_markings: IntegerArray(0 to 16)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 1);
      constant place_delays: IntegerArray(0 to 16) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_376"; 
      signal preds: BooleanArray(1 to 17); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(103) & maxPool4_CP_346_elements(107) & maxPool4_CP_346_elements(111) & maxPool4_CP_346_elements(115) & maxPool4_CP_346_elements(167) & maxPool4_CP_346_elements(171) & maxPool4_CP_346_elements(175) & maxPool4_CP_346_elements(179) & maxPool4_CP_346_elements(231) & maxPool4_CP_346_elements(235) & maxPool4_CP_346_elements(239) & maxPool4_CP_346_elements(243) & maxPool4_CP_346_elements(295) & maxPool4_CP_346_elements(299) & maxPool4_CP_346_elements(303) & maxPool4_CP_346_elements(307) & maxPool4_CP_346_elements(378);
      gj_maxPool4_cp_element_group_376 : generic_join generic map(name => joinName, number_of_predecessors => 17, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(376), clk => clk, reset => reset); --
    end block;
    -- CP-element group 377:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 377: predecessors 
    -- CP-element group 377: marked-predecessors 
    -- CP-element group 377: 	379 
    -- CP-element group 377: 	382 
    -- CP-element group 377: successors 
    -- CP-element group 377: 	379 
    -- CP-element group 377:  members (3) 
      -- CP-element group 377: 	 assign_stmt_97_to_assign_stmt_1138/CONCAT_u32_u64_1133_update_start_
      -- CP-element group 377: 	 assign_stmt_97_to_assign_stmt_1138/CONCAT_u32_u64_1133_Update/$entry
      -- CP-element group 377: 	 assign_stmt_97_to_assign_stmt_1138/CONCAT_u32_u64_1133_Update/cr
      -- 
    cr_2088_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2088_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(377), ack => CONCAT_u32_u64_1133_inst_req_1); -- 
    maxPool4_cp_element_group_377: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_377"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(379) & maxPool4_CP_346_elements(382);
      gj_maxPool4_cp_element_group_377 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(377), clk => clk, reset => reset); --
    end block;
    -- CP-element group 378:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 378: predecessors 
    -- CP-element group 378: 	376 
    -- CP-element group 378: successors 
    -- CP-element group 378: marked-successors 
    -- CP-element group 378: 	101 
    -- CP-element group 378: 	105 
    -- CP-element group 378: 	109 
    -- CP-element group 378: 	113 
    -- CP-element group 378: 	165 
    -- CP-element group 378: 	169 
    -- CP-element group 378: 	173 
    -- CP-element group 378: 	177 
    -- CP-element group 378: 	229 
    -- CP-element group 378: 	233 
    -- CP-element group 378: 	237 
    -- CP-element group 378: 	241 
    -- CP-element group 378: 	293 
    -- CP-element group 378: 	297 
    -- CP-element group 378: 	301 
    -- CP-element group 378: 	305 
    -- CP-element group 378: 	376 
    -- CP-element group 378:  members (3) 
      -- CP-element group 378: 	 assign_stmt_97_to_assign_stmt_1138/CONCAT_u32_u64_1133_sample_completed_
      -- CP-element group 378: 	 assign_stmt_97_to_assign_stmt_1138/CONCAT_u32_u64_1133_Sample/$exit
      -- CP-element group 378: 	 assign_stmt_97_to_assign_stmt_1138/CONCAT_u32_u64_1133_Sample/ra
      -- 
    ra_2084_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 378_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u32_u64_1133_inst_ack_0, ack => maxPool4_CP_346_elements(378)); -- 
    -- CP-element group 379:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 379: predecessors 
    -- CP-element group 379: 	377 
    -- CP-element group 379: successors 
    -- CP-element group 379: 	380 
    -- CP-element group 379: marked-successors 
    -- CP-element group 379: 	377 
    -- CP-element group 379:  members (3) 
      -- CP-element group 379: 	 assign_stmt_97_to_assign_stmt_1138/CONCAT_u32_u64_1133_update_completed_
      -- CP-element group 379: 	 assign_stmt_97_to_assign_stmt_1138/CONCAT_u32_u64_1133_Update/$exit
      -- CP-element group 379: 	 assign_stmt_97_to_assign_stmt_1138/CONCAT_u32_u64_1133_Update/ca
      -- 
    ca_2089_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 379_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u32_u64_1133_inst_ack_1, ack => maxPool4_CP_346_elements(379)); -- 
    -- CP-element group 380:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 380: predecessors 
    -- CP-element group 380: 	375 
    -- CP-element group 380: 	379 
    -- CP-element group 380: 	390 
    -- CP-element group 380: marked-predecessors 
    -- CP-element group 380: 	382 
    -- CP-element group 380: successors 
    -- CP-element group 380: 	382 
    -- CP-element group 380:  members (9) 
      -- CP-element group 380: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1122_sample_start_
      -- CP-element group 380: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1122_Sample/$entry
      -- CP-element group 380: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1122_Sample/ptr_deref_1122_Split/$entry
      -- CP-element group 380: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1122_Sample/ptr_deref_1122_Split/$exit
      -- CP-element group 380: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1122_Sample/ptr_deref_1122_Split/split_req
      -- CP-element group 380: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1122_Sample/ptr_deref_1122_Split/split_ack
      -- CP-element group 380: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1122_Sample/word_access_start/$entry
      -- CP-element group 380: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1122_Sample/word_access_start/word_0/$entry
      -- CP-element group 380: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1122_Sample/word_access_start/word_0/rr
      -- 
    rr_2127_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2127_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(380), ack => ptr_deref_1122_store_0_req_0); -- 
    maxPool4_cp_element_group_380: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_380"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(375) & maxPool4_CP_346_elements(379) & maxPool4_CP_346_elements(390) & maxPool4_CP_346_elements(382);
      gj_maxPool4_cp_element_group_380 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(380), clk => clk, reset => reset); --
    end block;
    -- CP-element group 381:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 381: predecessors 
    -- CP-element group 381: marked-predecessors 
    -- CP-element group 381: 	383 
    -- CP-element group 381: successors 
    -- CP-element group 381: 	383 
    -- CP-element group 381:  members (5) 
      -- CP-element group 381: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1122_update_start_
      -- CP-element group 381: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1122_Update/$entry
      -- CP-element group 381: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1122_Update/word_access_complete/$entry
      -- CP-element group 381: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1122_Update/word_access_complete/word_0/$entry
      -- CP-element group 381: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1122_Update/word_access_complete/word_0/cr
      -- 
    cr_2138_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2138_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(381), ack => ptr_deref_1122_store_0_req_1); -- 
    maxPool4_cp_element_group_381: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_381"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= maxPool4_CP_346_elements(383);
      gj_maxPool4_cp_element_group_381 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(381), clk => clk, reset => reset); --
    end block;
    -- CP-element group 382:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 382: predecessors 
    -- CP-element group 382: 	380 
    -- CP-element group 382: successors 
    -- CP-element group 382: 	391 
    -- CP-element group 382: marked-successors 
    -- CP-element group 382: 	323 
    -- CP-element group 382: 	373 
    -- CP-element group 382: 	377 
    -- CP-element group 382: 	380 
    -- CP-element group 382:  members (6) 
      -- CP-element group 382: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1122_sample_completed_
      -- CP-element group 382: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1122_Sample/$exit
      -- CP-element group 382: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1122_Sample/word_access_start/$exit
      -- CP-element group 382: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1122_Sample/word_access_start/word_0/$exit
      -- CP-element group 382: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1122_Sample/word_access_start/word_0/ra
      -- CP-element group 382: 	 assign_stmt_97_to_assign_stmt_1138/ring_reenable_memory_space_0
      -- 
    ra_2128_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 382_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1122_store_0_ack_0, ack => maxPool4_CP_346_elements(382)); -- 
    -- CP-element group 383:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 383: predecessors 
    -- CP-element group 383: 	381 
    -- CP-element group 383: successors 
    -- CP-element group 383: 	391 
    -- CP-element group 383: marked-successors 
    -- CP-element group 383: 	381 
    -- CP-element group 383:  members (5) 
      -- CP-element group 383: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1122_update_completed_
      -- CP-element group 383: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1122_Update/$exit
      -- CP-element group 383: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1122_Update/word_access_complete/$exit
      -- CP-element group 383: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1122_Update/word_access_complete/word_0/$exit
      -- CP-element group 383: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1122_Update/word_access_complete/word_0/ca
      -- 
    ca_2139_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 383_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1122_store_0_ack_1, ack => maxPool4_CP_346_elements(383)); -- 
    -- CP-element group 384:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 384: predecessors 
    -- CP-element group 384: 	55 
    -- CP-element group 384: 	119 
    -- CP-element group 384: 	183 
    -- CP-element group 384: 	247 
    -- CP-element group 384: marked-predecessors 
    -- CP-element group 384: 	386 
    -- CP-element group 384: successors 
    -- CP-element group 384: 	386 
    -- CP-element group 384:  members (3) 
      -- CP-element group 384: 	 assign_stmt_97_to_assign_stmt_1138/type_cast_1137_sample_start_
      -- CP-element group 384: 	 assign_stmt_97_to_assign_stmt_1138/type_cast_1137_Sample/$entry
      -- CP-element group 384: 	 assign_stmt_97_to_assign_stmt_1138/type_cast_1137_Sample/rr
      -- 
    rr_2147_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2147_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(384), ack => type_cast_1137_inst_req_0); -- 
    maxPool4_cp_element_group_384: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_384"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(55) & maxPool4_CP_346_elements(119) & maxPool4_CP_346_elements(183) & maxPool4_CP_346_elements(247) & maxPool4_CP_346_elements(386);
      gj_maxPool4_cp_element_group_384 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(384), clk => clk, reset => reset); --
    end block;
    -- CP-element group 385:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 385: predecessors 
    -- CP-element group 385: 	7 
    -- CP-element group 385: marked-predecessors 
    -- CP-element group 385: 	387 
    -- CP-element group 385: successors 
    -- CP-element group 385: 	387 
    -- CP-element group 385:  members (3) 
      -- CP-element group 385: 	 assign_stmt_97_to_assign_stmt_1138/type_cast_1137_update_start_
      -- CP-element group 385: 	 assign_stmt_97_to_assign_stmt_1138/type_cast_1137_Update/$entry
      -- CP-element group 385: 	 assign_stmt_97_to_assign_stmt_1138/type_cast_1137_Update/cr
      -- 
    cr_2152_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2152_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => maxPool4_CP_346_elements(385), ack => type_cast_1137_inst_req_1); -- 
    maxPool4_cp_element_group_385: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_385"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(7) & maxPool4_CP_346_elements(387);
      gj_maxPool4_cp_element_group_385 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(385), clk => clk, reset => reset); --
    end block;
    -- CP-element group 386:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 386: predecessors 
    -- CP-element group 386: 	384 
    -- CP-element group 386: successors 
    -- CP-element group 386: marked-successors 
    -- CP-element group 386: 	53 
    -- CP-element group 386: 	117 
    -- CP-element group 386: 	181 
    -- CP-element group 386: 	245 
    -- CP-element group 386: 	384 
    -- CP-element group 386:  members (3) 
      -- CP-element group 386: 	 assign_stmt_97_to_assign_stmt_1138/type_cast_1137_sample_completed_
      -- CP-element group 386: 	 assign_stmt_97_to_assign_stmt_1138/type_cast_1137_Sample/$exit
      -- CP-element group 386: 	 assign_stmt_97_to_assign_stmt_1138/type_cast_1137_Sample/ra
      -- 
    ra_2148_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 386_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1137_inst_ack_0, ack => maxPool4_CP_346_elements(386)); -- 
    -- CP-element group 387:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 387: predecessors 
    -- CP-element group 387: 	385 
    -- CP-element group 387: successors 
    -- CP-element group 387: 	391 
    -- CP-element group 387: marked-successors 
    -- CP-element group 387: 	385 
    -- CP-element group 387:  members (3) 
      -- CP-element group 387: 	 assign_stmt_97_to_assign_stmt_1138/type_cast_1137_update_completed_
      -- CP-element group 387: 	 assign_stmt_97_to_assign_stmt_1138/type_cast_1137_Update/$exit
      -- CP-element group 387: 	 assign_stmt_97_to_assign_stmt_1138/type_cast_1137_Update/ca
      -- 
    ca_2153_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 387_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1137_inst_ack_1, ack => maxPool4_CP_346_elements(387)); -- 
    -- CP-element group 388:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 388: predecessors 
    -- CP-element group 388: 	325 
    -- CP-element group 388: successors 
    -- CP-element group 388: 	342 
    -- CP-element group 388:  members (1) 
      -- CP-element group 388: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1044_ptr_deref_1070_delay
      -- 
    -- Element group maxPool4_CP_346_elements(388) is a control-delay.
    cp_element_388_delay: control_delay_element  generic map(name => " 388_delay", delay_value => 1)  port map(req => maxPool4_CP_346_elements(325), ack => maxPool4_CP_346_elements(388), clk => clk, reset =>reset);
    -- CP-element group 389:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 389: predecessors 
    -- CP-element group 389: 	344 
    -- CP-element group 389: successors 
    -- CP-element group 389: 	361 
    -- CP-element group 389:  members (1) 
      -- CP-element group 389: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1070_ptr_deref_1096_delay
      -- 
    -- Element group maxPool4_CP_346_elements(389) is a control-delay.
    cp_element_389_delay: control_delay_element  generic map(name => " 389_delay", delay_value => 1)  port map(req => maxPool4_CP_346_elements(344), ack => maxPool4_CP_346_elements(389), clk => clk, reset =>reset);
    -- CP-element group 390:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 390: predecessors 
    -- CP-element group 390: 	363 
    -- CP-element group 390: successors 
    -- CP-element group 390: 	380 
    -- CP-element group 390:  members (1) 
      -- CP-element group 390: 	 assign_stmt_97_to_assign_stmt_1138/ptr_deref_1096_ptr_deref_1122_delay
      -- 
    -- Element group maxPool4_CP_346_elements(390) is a control-delay.
    cp_element_390_delay: control_delay_element  generic map(name => " 390_delay", delay_value => 1)  port map(req => maxPool4_CP_346_elements(363), ack => maxPool4_CP_346_elements(390), clk => clk, reset =>reset);
    -- CP-element group 391:  join  transition  bypass  pipeline-parent 
    -- CP-element group 391: predecessors 
    -- CP-element group 391: 	11 
    -- CP-element group 391: 	18 
    -- CP-element group 391: 	25 
    -- CP-element group 391: 	32 
    -- CP-element group 391: 	311 
    -- CP-element group 391: 	326 
    -- CP-element group 391: 	330 
    -- CP-element group 391: 	345 
    -- CP-element group 391: 	349 
    -- CP-element group 391: 	364 
    -- CP-element group 391: 	368 
    -- CP-element group 391: 	382 
    -- CP-element group 391: 	383 
    -- CP-element group 391: 	387 
    -- CP-element group 391: successors 
    -- CP-element group 391: 	398 
    -- CP-element group 391:  members (1) 
      -- CP-element group 391: 	 assign_stmt_97_to_assign_stmt_1138/$exit
      -- 
    maxPool4_cp_element_group_391: block -- 
      constant place_capacities: IntegerArray(0 to 13) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 15,8 => 15,9 => 15,10 => 15,11 => 15,12 => 15,13 => 15);
      constant place_markings: IntegerArray(0 to 13)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0);
      constant place_delays: IntegerArray(0 to 13) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0);
      constant joinName: string(1 to 29) := "maxPool4_cp_element_group_391"; 
      signal preds: BooleanArray(1 to 14); -- 
    begin -- 
      preds <= maxPool4_CP_346_elements(11) & maxPool4_CP_346_elements(18) & maxPool4_CP_346_elements(25) & maxPool4_CP_346_elements(32) & maxPool4_CP_346_elements(311) & maxPool4_CP_346_elements(326) & maxPool4_CP_346_elements(330) & maxPool4_CP_346_elements(345) & maxPool4_CP_346_elements(349) & maxPool4_CP_346_elements(364) & maxPool4_CP_346_elements(368) & maxPool4_CP_346_elements(382) & maxPool4_CP_346_elements(383) & maxPool4_CP_346_elements(387);
      gj_maxPool4_cp_element_group_391 : generic_join generic map(name => joinName, number_of_predecessors => 14, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => maxPool4_CP_346_elements(391), clk => clk, reset => reset); --
    end block;
    -- CP-element group 392:  place  bypass  pipeline-parent 
    -- CP-element group 392: predecessors 
    -- CP-element group 392: 	2 
    -- CP-element group 392: successors 
    -- CP-element group 392:  members (1) 
      -- CP-element group 392: 	 addr_update_enable
      -- 
    maxPool4_CP_346_elements(392) <= maxPool4_CP_346_elements(2);
    -- CP-element group 393:  place  bypass  pipeline-parent 
    -- CP-element group 393: predecessors 
    -- CP-element group 393: 	3 
    -- CP-element group 393: successors 
    -- CP-element group 393:  members (1) 
      -- CP-element group 393: 	 addr1_update_enable
      -- 
    maxPool4_CP_346_elements(393) <= maxPool4_CP_346_elements(3);
    -- CP-element group 394:  place  bypass  pipeline-parent 
    -- CP-element group 394: predecessors 
    -- CP-element group 394: 	4 
    -- CP-element group 394: successors 
    -- CP-element group 394:  members (1) 
      -- CP-element group 394: 	 addr2_update_enable
      -- 
    maxPool4_CP_346_elements(394) <= maxPool4_CP_346_elements(4);
    -- CP-element group 395:  place  bypass  pipeline-parent 
    -- CP-element group 395: predecessors 
    -- CP-element group 395: 	5 
    -- CP-element group 395: successors 
    -- CP-element group 395:  members (1) 
      -- CP-element group 395: 	 addr3_update_enable
      -- 
    maxPool4_CP_346_elements(395) <= maxPool4_CP_346_elements(5);
    -- CP-element group 396:  place  bypass  pipeline-parent 
    -- CP-element group 396: predecessors 
    -- CP-element group 396: 	6 
    -- CP-element group 396: successors 
    -- CP-element group 396:  members (1) 
      -- CP-element group 396: 	 addr4_update_enable
      -- 
    maxPool4_CP_346_elements(396) <= maxPool4_CP_346_elements(6);
    -- CP-element group 397:  place  bypass  pipeline-parent 
    -- CP-element group 397: predecessors 
    -- CP-element group 397: successors 
    -- CP-element group 397: 	7 
    -- CP-element group 397:  members (1) 
      -- CP-element group 397: 	 output_update_enable
      -- 
    -- CP-element group 398:  transition  bypass  pipeline-parent 
    -- CP-element group 398: predecessors 
    -- CP-element group 398: 	391 
    -- CP-element group 398: successors 
    -- CP-element group 398:  members (1) 
      -- CP-element group 398: 	 $exit
      -- 
    maxPool4_CP_346_elements(398) <= maxPool4_CP_346_elements(391);
    --  hookup: inputs to control-path 
    maxPool4_CP_346_elements(397) <= output_update_enable;
    -- hookup: output from control-path 
    addr_update_enable <= maxPool4_CP_346_elements(392);
    addr1_update_enable <= maxPool4_CP_346_elements(393);
    addr2_update_enable <= maxPool4_CP_346_elements(394);
    addr3_update_enable <= maxPool4_CP_346_elements(395);
    addr4_update_enable <= maxPool4_CP_346_elements(396);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u32_u32_1062_resized : std_logic_vector(13 downto 0);
    signal ADD_u32_u32_1062_scaled : std_logic_vector(13 downto 0);
    signal ADD_u32_u32_1062_wire : std_logic_vector(31 downto 0);
    signal ADD_u32_u32_1088_resized : std_logic_vector(13 downto 0);
    signal ADD_u32_u32_1088_scaled : std_logic_vector(13 downto 0);
    signal ADD_u32_u32_1088_wire : std_logic_vector(31 downto 0);
    signal ADD_u32_u32_1114_resized : std_logic_vector(13 downto 0);
    signal ADD_u32_u32_1114_scaled : std_logic_vector(13 downto 0);
    signal ADD_u32_u32_1114_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u16_u32_1049_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u16_u32_1054_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u16_u32_1075_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u16_u32_1080_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u16_u32_1101_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u16_u32_1106_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u16_u32_1127_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u16_u32_1132_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u32_u64_1055_wire : std_logic_vector(63 downto 0);
    signal CONCAT_u32_u64_1081_wire : std_logic_vector(63 downto 0);
    signal CONCAT_u32_u64_1107_wire : std_logic_vector(63 downto 0);
    signal CONCAT_u32_u64_1133_wire : std_logic_vector(63 downto 0);
    signal R_addr1_94_resized : std_logic_vector(13 downto 0);
    signal R_addr1_94_scaled : std_logic_vector(13 downto 0);
    signal R_addr2_101_resized : std_logic_vector(13 downto 0);
    signal R_addr2_101_scaled : std_logic_vector(13 downto 0);
    signal R_addr3_108_resized : std_logic_vector(13 downto 0);
    signal R_addr3_108_scaled : std_logic_vector(13 downto 0);
    signal R_addr4_115_resized : std_logic_vector(13 downto 0);
    signal R_addr4_115_scaled : std_logic_vector(13 downto 0);
    signal R_addr_1036_resized : std_logic_vector(13 downto 0);
    signal R_addr_1036_scaled : std_logic_vector(13 downto 0);
    signal SGT_i16_u1_1004_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_1012_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_1020_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_1028_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_652_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_660_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_668_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_676_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_684_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_692_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_700_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_708_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_716_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_724_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_732_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_740_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_748_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_756_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_764_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_772_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_780_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_788_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_796_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_804_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_812_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_820_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_828_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_836_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_844_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_852_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_860_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_868_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_876_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_884_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_892_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_900_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_908_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_916_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_924_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_932_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_940_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_948_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_956_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_964_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_972_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_980_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_988_wire : std_logic_vector(0 downto 0);
    signal SGT_i16_u1_996_wire : std_logic_vector(0 downto 0);
    signal a110_432 : std_logic_vector(15 downto 0);
    signal a111_436 : std_logic_vector(15 downto 0);
    signal a112_440 : std_logic_vector(15 downto 0);
    signal a113_444 : std_logic_vector(15 downto 0);
    signal a114_448 : std_logic_vector(15 downto 0);
    signal a115_452 : std_logic_vector(15 downto 0);
    signal a116_456 : std_logic_vector(15 downto 0);
    signal a11_396 : std_logic_vector(15 downto 0);
    signal a12_400 : std_logic_vector(15 downto 0);
    signal a13_404 : std_logic_vector(15 downto 0);
    signal a14_408 : std_logic_vector(15 downto 0);
    signal a15_412 : std_logic_vector(15 downto 0);
    signal a16_416 : std_logic_vector(15 downto 0);
    signal a17_420 : std_logic_vector(15 downto 0);
    signal a18_424 : std_logic_vector(15 downto 0);
    signal a19_428 : std_logic_vector(15 downto 0);
    signal a210_496 : std_logic_vector(15 downto 0);
    signal a211_500 : std_logic_vector(15 downto 0);
    signal a212_504 : std_logic_vector(15 downto 0);
    signal a213_508 : std_logic_vector(15 downto 0);
    signal a214_512 : std_logic_vector(15 downto 0);
    signal a215_516 : std_logic_vector(15 downto 0);
    signal a216_520 : std_logic_vector(15 downto 0);
    signal a21_460 : std_logic_vector(15 downto 0);
    signal a22_464 : std_logic_vector(15 downto 0);
    signal a23_468 : std_logic_vector(15 downto 0);
    signal a24_472 : std_logic_vector(15 downto 0);
    signal a25_476 : std_logic_vector(15 downto 0);
    signal a26_480 : std_logic_vector(15 downto 0);
    signal a27_484 : std_logic_vector(15 downto 0);
    signal a28_488 : std_logic_vector(15 downto 0);
    signal a29_492 : std_logic_vector(15 downto 0);
    signal a310_560 : std_logic_vector(15 downto 0);
    signal a311_564 : std_logic_vector(15 downto 0);
    signal a312_568 : std_logic_vector(15 downto 0);
    signal a313_572 : std_logic_vector(15 downto 0);
    signal a314_576 : std_logic_vector(15 downto 0);
    signal a315_580 : std_logic_vector(15 downto 0);
    signal a316_584 : std_logic_vector(15 downto 0);
    signal a31_524 : std_logic_vector(15 downto 0);
    signal a32_528 : std_logic_vector(15 downto 0);
    signal a33_532 : std_logic_vector(15 downto 0);
    signal a34_536 : std_logic_vector(15 downto 0);
    signal a35_540 : std_logic_vector(15 downto 0);
    signal a36_544 : std_logic_vector(15 downto 0);
    signal a37_548 : std_logic_vector(15 downto 0);
    signal a38_552 : std_logic_vector(15 downto 0);
    signal a39_556 : std_logic_vector(15 downto 0);
    signal a410_624 : std_logic_vector(15 downto 0);
    signal a411_628 : std_logic_vector(15 downto 0);
    signal a412_632 : std_logic_vector(15 downto 0);
    signal a413_636 : std_logic_vector(15 downto 0);
    signal a414_640 : std_logic_vector(15 downto 0);
    signal a415_644 : std_logic_vector(15 downto 0);
    signal a416_648 : std_logic_vector(15 downto 0);
    signal a41_588 : std_logic_vector(15 downto 0);
    signal a42_592 : std_logic_vector(15 downto 0);
    signal a43_596 : std_logic_vector(15 downto 0);
    signal a44_600 : std_logic_vector(15 downto 0);
    signal a45_604 : std_logic_vector(15 downto 0);
    signal a46_608 : std_logic_vector(15 downto 0);
    signal a47_612 : std_logic_vector(15 downto 0);
    signal a48_616 : std_logic_vector(15 downto 0);
    signal a49_620 : std_logic_vector(15 downto 0);
    signal array_obj_ref_102_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_102_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_102_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_102_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_102_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_102_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1037_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1037_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1037_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1037_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1037_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1037_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1063_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1063_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1063_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1063_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1063_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1063_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1089_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1089_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1089_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1089_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1089_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1089_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_109_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_109_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_109_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_109_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_109_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_109_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1115_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1115_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1115_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1115_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1115_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1115_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_116_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_116_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_116_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_116_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_116_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_116_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_95_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_95_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_95_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_95_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_95_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_95_root_address : std_logic_vector(13 downto 0);
    signal c1_122 : std_logic_vector(255 downto 0);
    signal c2_126 : std_logic_vector(255 downto 0);
    signal c3_130 : std_logic_vector(255 downto 0);
    signal c4_134 : std_logic_vector(255 downto 0);
    signal konst_1061_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1087_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1113_wire_constant : std_logic_vector(31 downto 0);
    signal myptr1_97 : std_logic_vector(31 downto 0);
    signal myptr2_104 : std_logic_vector(31 downto 0);
    signal myptr3_111 : std_logic_vector(31 downto 0);
    signal myptr4_118 : std_logic_vector(31 downto 0);
    signal myptr5_1039 : std_logic_vector(31 downto 0);
    signal myptr5_1040_delayed_8_0_1042 : std_logic_vector(31 downto 0);
    signal myptr6_1063_delayed_8_0_1068 : std_logic_vector(31 downto 0);
    signal myptr6_1065 : std_logic_vector(31 downto 0);
    signal myptr7_1086_delayed_8_0_1094 : std_logic_vector(31 downto 0);
    signal myptr7_1091 : std_logic_vector(31 downto 0);
    signal myptr8_1109_delayed_8_0_1120 : std_logic_vector(31 downto 0);
    signal myptr8_1117 : std_logic_vector(31 downto 0);
    signal out10_888 : std_logic_vector(15 downto 0);
    signal out11_912 : std_logic_vector(15 downto 0);
    signal out12_936 : std_logic_vector(15 downto 0);
    signal out13_960 : std_logic_vector(15 downto 0);
    signal out14_984 : std_logic_vector(15 downto 0);
    signal out15_1008 : std_logic_vector(15 downto 0);
    signal out16_1032 : std_logic_vector(15 downto 0);
    signal out1_672 : std_logic_vector(15 downto 0);
    signal out2_696 : std_logic_vector(15 downto 0);
    signal out3_720 : std_logic_vector(15 downto 0);
    signal out4_744 : std_logic_vector(15 downto 0);
    signal out5_768 : std_logic_vector(15 downto 0);
    signal out6_792 : std_logic_vector(15 downto 0);
    signal out7_816 : std_logic_vector(15 downto 0);
    signal out8_840 : std_logic_vector(15 downto 0);
    signal out9_864 : std_logic_vector(15 downto 0);
    signal ptr_deref_1044_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1044_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1044_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1044_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1044_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1044_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1070_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1070_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1070_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1070_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1070_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1070_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1096_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1096_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1096_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1096_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1096_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1096_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1122_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1122_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1122_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1122_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1122_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1122_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_121_data_0 : std_logic_vector(255 downto 0);
    signal ptr_deref_121_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_121_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_121_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_121_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_125_data_0 : std_logic_vector(255 downto 0);
    signal ptr_deref_125_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_125_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_125_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_125_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_129_data_0 : std_logic_vector(255 downto 0);
    signal ptr_deref_129_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_129_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_129_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_129_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_133_data_0 : std_logic_vector(255 downto 0);
    signal ptr_deref_133_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_133_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_133_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_133_word_offset_0 : std_logic_vector(13 downto 0);
    signal sliced_v110_175 : std_logic_vector(15 downto 0);
    signal sliced_v111_179 : std_logic_vector(15 downto 0);
    signal sliced_v112_183 : std_logic_vector(15 downto 0);
    signal sliced_v113_187 : std_logic_vector(15 downto 0);
    signal sliced_v114_191 : std_logic_vector(15 downto 0);
    signal sliced_v115_195 : std_logic_vector(15 downto 0);
    signal sliced_v116_199 : std_logic_vector(15 downto 0);
    signal sliced_v11_139 : std_logic_vector(15 downto 0);
    signal sliced_v12_143 : std_logic_vector(15 downto 0);
    signal sliced_v13_147 : std_logic_vector(15 downto 0);
    signal sliced_v14_151 : std_logic_vector(15 downto 0);
    signal sliced_v15_155 : std_logic_vector(15 downto 0);
    signal sliced_v16_159 : std_logic_vector(15 downto 0);
    signal sliced_v17_163 : std_logic_vector(15 downto 0);
    signal sliced_v18_167 : std_logic_vector(15 downto 0);
    signal sliced_v19_171 : std_logic_vector(15 downto 0);
    signal sliced_v210_239 : std_logic_vector(15 downto 0);
    signal sliced_v211_243 : std_logic_vector(15 downto 0);
    signal sliced_v212_247 : std_logic_vector(15 downto 0);
    signal sliced_v213_251 : std_logic_vector(15 downto 0);
    signal sliced_v214_255 : std_logic_vector(15 downto 0);
    signal sliced_v215_259 : std_logic_vector(15 downto 0);
    signal sliced_v216_263 : std_logic_vector(15 downto 0);
    signal sliced_v21_203 : std_logic_vector(15 downto 0);
    signal sliced_v22_207 : std_logic_vector(15 downto 0);
    signal sliced_v23_211 : std_logic_vector(15 downto 0);
    signal sliced_v24_215 : std_logic_vector(15 downto 0);
    signal sliced_v25_219 : std_logic_vector(15 downto 0);
    signal sliced_v26_223 : std_logic_vector(15 downto 0);
    signal sliced_v27_227 : std_logic_vector(15 downto 0);
    signal sliced_v28_231 : std_logic_vector(15 downto 0);
    signal sliced_v29_235 : std_logic_vector(15 downto 0);
    signal sliced_v310_303 : std_logic_vector(15 downto 0);
    signal sliced_v311_307 : std_logic_vector(15 downto 0);
    signal sliced_v312_311 : std_logic_vector(15 downto 0);
    signal sliced_v313_315 : std_logic_vector(15 downto 0);
    signal sliced_v314_319 : std_logic_vector(15 downto 0);
    signal sliced_v315_323 : std_logic_vector(15 downto 0);
    signal sliced_v316_327 : std_logic_vector(15 downto 0);
    signal sliced_v31_267 : std_logic_vector(15 downto 0);
    signal sliced_v32_271 : std_logic_vector(15 downto 0);
    signal sliced_v33_275 : std_logic_vector(15 downto 0);
    signal sliced_v34_279 : std_logic_vector(15 downto 0);
    signal sliced_v35_283 : std_logic_vector(15 downto 0);
    signal sliced_v36_287 : std_logic_vector(15 downto 0);
    signal sliced_v37_291 : std_logic_vector(15 downto 0);
    signal sliced_v38_295 : std_logic_vector(15 downto 0);
    signal sliced_v39_299 : std_logic_vector(15 downto 0);
    signal sliced_v410_367 : std_logic_vector(15 downto 0);
    signal sliced_v411_371 : std_logic_vector(15 downto 0);
    signal sliced_v412_375 : std_logic_vector(15 downto 0);
    signal sliced_v413_379 : std_logic_vector(15 downto 0);
    signal sliced_v414_383 : std_logic_vector(15 downto 0);
    signal sliced_v415_387 : std_logic_vector(15 downto 0);
    signal sliced_v416_391 : std_logic_vector(15 downto 0);
    signal sliced_v41_331 : std_logic_vector(15 downto 0);
    signal sliced_v42_335 : std_logic_vector(15 downto 0);
    signal sliced_v43_339 : std_logic_vector(15 downto 0);
    signal sliced_v44_343 : std_logic_vector(15 downto 0);
    signal sliced_v45_347 : std_logic_vector(15 downto 0);
    signal sliced_v46_351 : std_logic_vector(15 downto 0);
    signal sliced_v47_355 : std_logic_vector(15 downto 0);
    signal sliced_v48_359 : std_logic_vector(15 downto 0);
    signal sliced_v49_363 : std_logic_vector(15 downto 0);
    signal t101_872 : std_logic_vector(15 downto 0);
    signal t102_880 : std_logic_vector(15 downto 0);
    signal t111_896 : std_logic_vector(15 downto 0);
    signal t112_904 : std_logic_vector(15 downto 0);
    signal t11_656 : std_logic_vector(15 downto 0);
    signal t121_920 : std_logic_vector(15 downto 0);
    signal t122_928 : std_logic_vector(15 downto 0);
    signal t12_664 : std_logic_vector(15 downto 0);
    signal t131_944 : std_logic_vector(15 downto 0);
    signal t132_952 : std_logic_vector(15 downto 0);
    signal t141_968 : std_logic_vector(15 downto 0);
    signal t142_976 : std_logic_vector(15 downto 0);
    signal t151_992 : std_logic_vector(15 downto 0);
    signal t152_1000 : std_logic_vector(15 downto 0);
    signal t161_1016 : std_logic_vector(15 downto 0);
    signal t162_1024 : std_logic_vector(15 downto 0);
    signal t21_680 : std_logic_vector(15 downto 0);
    signal t22_688 : std_logic_vector(15 downto 0);
    signal t31_704 : std_logic_vector(15 downto 0);
    signal t32_712 : std_logic_vector(15 downto 0);
    signal t41_728 : std_logic_vector(15 downto 0);
    signal t42_736 : std_logic_vector(15 downto 0);
    signal t51_752 : std_logic_vector(15 downto 0);
    signal t52_760 : std_logic_vector(15 downto 0);
    signal t61_776 : std_logic_vector(15 downto 0);
    signal t62_784 : std_logic_vector(15 downto 0);
    signal t71_800 : std_logic_vector(15 downto 0);
    signal t72_808 : std_logic_vector(15 downto 0);
    signal t81_824 : std_logic_vector(15 downto 0);
    signal t82_832 : std_logic_vector(15 downto 0);
    signal t91_848 : std_logic_vector(15 downto 0);
    signal t92_856 : std_logic_vector(15 downto 0);
    signal type_cast_1046_wire : std_logic_vector(15 downto 0);
    signal type_cast_1048_wire : std_logic_vector(15 downto 0);
    signal type_cast_1051_wire : std_logic_vector(15 downto 0);
    signal type_cast_1053_wire : std_logic_vector(15 downto 0);
    signal type_cast_1072_wire : std_logic_vector(15 downto 0);
    signal type_cast_1074_wire : std_logic_vector(15 downto 0);
    signal type_cast_1077_wire : std_logic_vector(15 downto 0);
    signal type_cast_1079_wire : std_logic_vector(15 downto 0);
    signal type_cast_1098_wire : std_logic_vector(15 downto 0);
    signal type_cast_1100_wire : std_logic_vector(15 downto 0);
    signal type_cast_1103_wire : std_logic_vector(15 downto 0);
    signal type_cast_1105_wire : std_logic_vector(15 downto 0);
    signal type_cast_1124_wire : std_logic_vector(15 downto 0);
    signal type_cast_1126_wire : std_logic_vector(15 downto 0);
    signal type_cast_1129_wire : std_logic_vector(15 downto 0);
    signal type_cast_1131_wire : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_102_constant_part_of_offset <= "00000000000000";
    array_obj_ref_102_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_102_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_102_resized_base_address <= "00000000000000";
    array_obj_ref_1037_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1037_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1037_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1037_resized_base_address <= "00000000000000";
    array_obj_ref_1063_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1063_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1063_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1063_resized_base_address <= "00000000000000";
    array_obj_ref_1089_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1089_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1089_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1089_resized_base_address <= "00000000000000";
    array_obj_ref_109_constant_part_of_offset <= "00000000000000";
    array_obj_ref_109_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_109_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_109_resized_base_address <= "00000000000000";
    array_obj_ref_1115_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1115_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1115_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1115_resized_base_address <= "00000000000000";
    array_obj_ref_116_constant_part_of_offset <= "00000000000000";
    array_obj_ref_116_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_116_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_116_resized_base_address <= "00000000000000";
    array_obj_ref_95_constant_part_of_offset <= "00000000000000";
    array_obj_ref_95_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_95_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_95_resized_base_address <= "00000000000000";
    konst_1061_wire_constant <= "00000000000000000000000000000001";
    konst_1087_wire_constant <= "00000000000000000000000000000010";
    konst_1113_wire_constant <= "00000000000000000000000000000011";
    ptr_deref_1044_word_offset_0 <= "00000000000000";
    ptr_deref_1070_word_offset_0 <= "00000000000000";
    ptr_deref_1096_word_offset_0 <= "00000000000000";
    ptr_deref_1122_word_offset_0 <= "00000000000000";
    ptr_deref_121_word_offset_0 <= "00000000000000";
    ptr_deref_125_word_offset_0 <= "00000000000000";
    ptr_deref_129_word_offset_0 <= "00000000000000";
    ptr_deref_133_word_offset_0 <= "00000000000000";
    -- flow-through select operator MUX_1007_inst
    out15_1008 <= t151_992 when (SGT_i16_u1_1004_wire(0) /=  '0') else t152_1000;
    -- flow-through select operator MUX_1015_inst
    t161_1016 <= a116_456 when (SGT_i16_u1_1012_wire(0) /=  '0') else a216_520;
    -- flow-through select operator MUX_1023_inst
    t162_1024 <= a316_584 when (SGT_i16_u1_1020_wire(0) /=  '0') else a416_648;
    -- flow-through select operator MUX_1031_inst
    out16_1032 <= t161_1016 when (SGT_i16_u1_1028_wire(0) /=  '0') else t162_1024;
    -- flow-through select operator MUX_655_inst
    t11_656 <= a11_396 when (SGT_i16_u1_652_wire(0) /=  '0') else a21_460;
    -- flow-through select operator MUX_663_inst
    t12_664 <= a31_524 when (SGT_i16_u1_660_wire(0) /=  '0') else a41_588;
    -- flow-through select operator MUX_671_inst
    out1_672 <= t11_656 when (SGT_i16_u1_668_wire(0) /=  '0') else t12_664;
    -- flow-through select operator MUX_679_inst
    t21_680 <= a12_400 when (SGT_i16_u1_676_wire(0) /=  '0') else a22_464;
    -- flow-through select operator MUX_687_inst
    t22_688 <= a32_528 when (SGT_i16_u1_684_wire(0) /=  '0') else a42_592;
    -- flow-through select operator MUX_695_inst
    out2_696 <= t21_680 when (SGT_i16_u1_692_wire(0) /=  '0') else t22_688;
    -- flow-through select operator MUX_703_inst
    t31_704 <= a13_404 when (SGT_i16_u1_700_wire(0) /=  '0') else a23_468;
    -- flow-through select operator MUX_711_inst
    t32_712 <= a33_532 when (SGT_i16_u1_708_wire(0) /=  '0') else a43_596;
    -- flow-through select operator MUX_719_inst
    out3_720 <= t31_704 when (SGT_i16_u1_716_wire(0) /=  '0') else t32_712;
    -- flow-through select operator MUX_727_inst
    t41_728 <= a14_408 when (SGT_i16_u1_724_wire(0) /=  '0') else a24_472;
    -- flow-through select operator MUX_735_inst
    t42_736 <= a34_536 when (SGT_i16_u1_732_wire(0) /=  '0') else a44_600;
    -- flow-through select operator MUX_743_inst
    out4_744 <= t41_728 when (SGT_i16_u1_740_wire(0) /=  '0') else t42_736;
    -- flow-through select operator MUX_751_inst
    t51_752 <= a15_412 when (SGT_i16_u1_748_wire(0) /=  '0') else a25_476;
    -- flow-through select operator MUX_759_inst
    t52_760 <= a35_540 when (SGT_i16_u1_756_wire(0) /=  '0') else a45_604;
    -- flow-through select operator MUX_767_inst
    out5_768 <= t51_752 when (SGT_i16_u1_764_wire(0) /=  '0') else t52_760;
    -- flow-through select operator MUX_775_inst
    t61_776 <= a16_416 when (SGT_i16_u1_772_wire(0) /=  '0') else a26_480;
    -- flow-through select operator MUX_783_inst
    t62_784 <= a36_544 when (SGT_i16_u1_780_wire(0) /=  '0') else a46_608;
    -- flow-through select operator MUX_791_inst
    out6_792 <= t61_776 when (SGT_i16_u1_788_wire(0) /=  '0') else t62_784;
    -- flow-through select operator MUX_799_inst
    t71_800 <= a17_420 when (SGT_i16_u1_796_wire(0) /=  '0') else a27_484;
    -- flow-through select operator MUX_807_inst
    t72_808 <= a37_548 when (SGT_i16_u1_804_wire(0) /=  '0') else a47_612;
    -- flow-through select operator MUX_815_inst
    out7_816 <= t71_800 when (SGT_i16_u1_812_wire(0) /=  '0') else t72_808;
    -- flow-through select operator MUX_823_inst
    t81_824 <= a18_424 when (SGT_i16_u1_820_wire(0) /=  '0') else a28_488;
    -- flow-through select operator MUX_831_inst
    t82_832 <= a38_552 when (SGT_i16_u1_828_wire(0) /=  '0') else a48_616;
    -- flow-through select operator MUX_839_inst
    out8_840 <= t81_824 when (SGT_i16_u1_836_wire(0) /=  '0') else t82_832;
    -- flow-through select operator MUX_847_inst
    t91_848 <= a19_428 when (SGT_i16_u1_844_wire(0) /=  '0') else a29_492;
    -- flow-through select operator MUX_855_inst
    t92_856 <= a39_556 when (SGT_i16_u1_852_wire(0) /=  '0') else a49_620;
    -- flow-through select operator MUX_863_inst
    out9_864 <= t91_848 when (SGT_i16_u1_860_wire(0) /=  '0') else t92_856;
    -- flow-through select operator MUX_871_inst
    t101_872 <= a110_432 when (SGT_i16_u1_868_wire(0) /=  '0') else a210_496;
    -- flow-through select operator MUX_879_inst
    t102_880 <= a310_560 when (SGT_i16_u1_876_wire(0) /=  '0') else a410_624;
    -- flow-through select operator MUX_887_inst
    out10_888 <= t101_872 when (SGT_i16_u1_884_wire(0) /=  '0') else t102_880;
    -- flow-through select operator MUX_895_inst
    t111_896 <= a111_436 when (SGT_i16_u1_892_wire(0) /=  '0') else a211_500;
    -- flow-through select operator MUX_903_inst
    t112_904 <= a311_564 when (SGT_i16_u1_900_wire(0) /=  '0') else a411_628;
    -- flow-through select operator MUX_911_inst
    out11_912 <= t111_896 when (SGT_i16_u1_908_wire(0) /=  '0') else t112_904;
    -- flow-through select operator MUX_919_inst
    t121_920 <= a112_440 when (SGT_i16_u1_916_wire(0) /=  '0') else a212_504;
    -- flow-through select operator MUX_927_inst
    t122_928 <= a312_568 when (SGT_i16_u1_924_wire(0) /=  '0') else a412_632;
    -- flow-through select operator MUX_935_inst
    out12_936 <= t121_920 when (SGT_i16_u1_932_wire(0) /=  '0') else t122_928;
    -- flow-through select operator MUX_943_inst
    t131_944 <= a113_444 when (SGT_i16_u1_940_wire(0) /=  '0') else a213_508;
    -- flow-through select operator MUX_951_inst
    t132_952 <= a313_572 when (SGT_i16_u1_948_wire(0) /=  '0') else a413_636;
    -- flow-through select operator MUX_959_inst
    out13_960 <= t131_944 when (SGT_i16_u1_956_wire(0) /=  '0') else t132_952;
    -- flow-through select operator MUX_967_inst
    t141_968 <= a114_448 when (SGT_i16_u1_964_wire(0) /=  '0') else a214_512;
    -- flow-through select operator MUX_975_inst
    t142_976 <= a314_576 when (SGT_i16_u1_972_wire(0) /=  '0') else a414_640;
    -- flow-through select operator MUX_983_inst
    out14_984 <= t141_968 when (SGT_i16_u1_980_wire(0) /=  '0') else t142_976;
    -- flow-through select operator MUX_991_inst
    t151_992 <= a115_452 when (SGT_i16_u1_988_wire(0) /=  '0') else a215_516;
    -- flow-through select operator MUX_999_inst
    t152_1000 <= a315_580 when (SGT_i16_u1_996_wire(0) /=  '0') else a415_644;
    slice_138_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_138_inst_req_0;
      slice_138_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_138_inst_req_1;
      slice_138_inst_ack_1<= update_ack(0);
      slice_138_inst: SliceSplitProtocol generic map(name => "slice_138_inst", in_data_width => 256, high_index => 255, low_index => 240, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_122, dout => sliced_v11_139, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_142_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_142_inst_req_0;
      slice_142_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_142_inst_req_1;
      slice_142_inst_ack_1<= update_ack(0);
      slice_142_inst: SliceSplitProtocol generic map(name => "slice_142_inst", in_data_width => 256, high_index => 239, low_index => 224, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_122, dout => sliced_v12_143, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_146_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_146_inst_req_0;
      slice_146_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_146_inst_req_1;
      slice_146_inst_ack_1<= update_ack(0);
      slice_146_inst: SliceSplitProtocol generic map(name => "slice_146_inst", in_data_width => 256, high_index => 223, low_index => 208, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_122, dout => sliced_v13_147, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_150_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_150_inst_req_0;
      slice_150_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_150_inst_req_1;
      slice_150_inst_ack_1<= update_ack(0);
      slice_150_inst: SliceSplitProtocol generic map(name => "slice_150_inst", in_data_width => 256, high_index => 207, low_index => 192, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_122, dout => sliced_v14_151, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_154_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_154_inst_req_0;
      slice_154_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_154_inst_req_1;
      slice_154_inst_ack_1<= update_ack(0);
      slice_154_inst: SliceSplitProtocol generic map(name => "slice_154_inst", in_data_width => 256, high_index => 191, low_index => 176, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_122, dout => sliced_v15_155, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_158_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_158_inst_req_0;
      slice_158_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_158_inst_req_1;
      slice_158_inst_ack_1<= update_ack(0);
      slice_158_inst: SliceSplitProtocol generic map(name => "slice_158_inst", in_data_width => 256, high_index => 175, low_index => 160, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_122, dout => sliced_v16_159, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_162_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_162_inst_req_0;
      slice_162_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_162_inst_req_1;
      slice_162_inst_ack_1<= update_ack(0);
      slice_162_inst: SliceSplitProtocol generic map(name => "slice_162_inst", in_data_width => 256, high_index => 159, low_index => 144, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_122, dout => sliced_v17_163, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_166_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_166_inst_req_0;
      slice_166_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_166_inst_req_1;
      slice_166_inst_ack_1<= update_ack(0);
      slice_166_inst: SliceSplitProtocol generic map(name => "slice_166_inst", in_data_width => 256, high_index => 143, low_index => 128, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_122, dout => sliced_v18_167, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_170_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_170_inst_req_0;
      slice_170_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_170_inst_req_1;
      slice_170_inst_ack_1<= update_ack(0);
      slice_170_inst: SliceSplitProtocol generic map(name => "slice_170_inst", in_data_width => 256, high_index => 127, low_index => 112, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_122, dout => sliced_v19_171, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_174_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_174_inst_req_0;
      slice_174_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_174_inst_req_1;
      slice_174_inst_ack_1<= update_ack(0);
      slice_174_inst: SliceSplitProtocol generic map(name => "slice_174_inst", in_data_width => 256, high_index => 111, low_index => 96, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_122, dout => sliced_v110_175, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_178_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_178_inst_req_0;
      slice_178_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_178_inst_req_1;
      slice_178_inst_ack_1<= update_ack(0);
      slice_178_inst: SliceSplitProtocol generic map(name => "slice_178_inst", in_data_width => 256, high_index => 95, low_index => 80, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_122, dout => sliced_v111_179, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_182_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_182_inst_req_0;
      slice_182_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_182_inst_req_1;
      slice_182_inst_ack_1<= update_ack(0);
      slice_182_inst: SliceSplitProtocol generic map(name => "slice_182_inst", in_data_width => 256, high_index => 79, low_index => 64, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_122, dout => sliced_v112_183, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_186_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_186_inst_req_0;
      slice_186_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_186_inst_req_1;
      slice_186_inst_ack_1<= update_ack(0);
      slice_186_inst: SliceSplitProtocol generic map(name => "slice_186_inst", in_data_width => 256, high_index => 63, low_index => 48, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_122, dout => sliced_v113_187, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_190_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_190_inst_req_0;
      slice_190_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_190_inst_req_1;
      slice_190_inst_ack_1<= update_ack(0);
      slice_190_inst: SliceSplitProtocol generic map(name => "slice_190_inst", in_data_width => 256, high_index => 47, low_index => 32, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_122, dout => sliced_v114_191, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_194_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_194_inst_req_0;
      slice_194_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_194_inst_req_1;
      slice_194_inst_ack_1<= update_ack(0);
      slice_194_inst: SliceSplitProtocol generic map(name => "slice_194_inst", in_data_width => 256, high_index => 31, low_index => 16, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_122, dout => sliced_v115_195, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_198_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_198_inst_req_0;
      slice_198_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_198_inst_req_1;
      slice_198_inst_ack_1<= update_ack(0);
      slice_198_inst: SliceSplitProtocol generic map(name => "slice_198_inst", in_data_width => 256, high_index => 15, low_index => 0, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c1_122, dout => sliced_v116_199, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_202_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_202_inst_req_0;
      slice_202_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_202_inst_req_1;
      slice_202_inst_ack_1<= update_ack(0);
      slice_202_inst: SliceSplitProtocol generic map(name => "slice_202_inst", in_data_width => 256, high_index => 255, low_index => 240, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_126, dout => sliced_v21_203, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_206_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_206_inst_req_0;
      slice_206_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_206_inst_req_1;
      slice_206_inst_ack_1<= update_ack(0);
      slice_206_inst: SliceSplitProtocol generic map(name => "slice_206_inst", in_data_width => 256, high_index => 239, low_index => 224, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_126, dout => sliced_v22_207, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_210_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_210_inst_req_0;
      slice_210_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_210_inst_req_1;
      slice_210_inst_ack_1<= update_ack(0);
      slice_210_inst: SliceSplitProtocol generic map(name => "slice_210_inst", in_data_width => 256, high_index => 223, low_index => 208, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_126, dout => sliced_v23_211, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_214_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_214_inst_req_0;
      slice_214_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_214_inst_req_1;
      slice_214_inst_ack_1<= update_ack(0);
      slice_214_inst: SliceSplitProtocol generic map(name => "slice_214_inst", in_data_width => 256, high_index => 207, low_index => 192, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_126, dout => sliced_v24_215, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_218_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_218_inst_req_0;
      slice_218_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_218_inst_req_1;
      slice_218_inst_ack_1<= update_ack(0);
      slice_218_inst: SliceSplitProtocol generic map(name => "slice_218_inst", in_data_width => 256, high_index => 191, low_index => 176, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_126, dout => sliced_v25_219, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_222_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_222_inst_req_0;
      slice_222_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_222_inst_req_1;
      slice_222_inst_ack_1<= update_ack(0);
      slice_222_inst: SliceSplitProtocol generic map(name => "slice_222_inst", in_data_width => 256, high_index => 175, low_index => 160, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_126, dout => sliced_v26_223, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_226_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_226_inst_req_0;
      slice_226_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_226_inst_req_1;
      slice_226_inst_ack_1<= update_ack(0);
      slice_226_inst: SliceSplitProtocol generic map(name => "slice_226_inst", in_data_width => 256, high_index => 159, low_index => 144, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_126, dout => sliced_v27_227, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_230_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_230_inst_req_0;
      slice_230_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_230_inst_req_1;
      slice_230_inst_ack_1<= update_ack(0);
      slice_230_inst: SliceSplitProtocol generic map(name => "slice_230_inst", in_data_width => 256, high_index => 143, low_index => 128, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_126, dout => sliced_v28_231, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_234_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_234_inst_req_0;
      slice_234_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_234_inst_req_1;
      slice_234_inst_ack_1<= update_ack(0);
      slice_234_inst: SliceSplitProtocol generic map(name => "slice_234_inst", in_data_width => 256, high_index => 127, low_index => 112, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_126, dout => sliced_v29_235, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_238_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_238_inst_req_0;
      slice_238_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_238_inst_req_1;
      slice_238_inst_ack_1<= update_ack(0);
      slice_238_inst: SliceSplitProtocol generic map(name => "slice_238_inst", in_data_width => 256, high_index => 111, low_index => 96, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_126, dout => sliced_v210_239, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_242_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_242_inst_req_0;
      slice_242_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_242_inst_req_1;
      slice_242_inst_ack_1<= update_ack(0);
      slice_242_inst: SliceSplitProtocol generic map(name => "slice_242_inst", in_data_width => 256, high_index => 95, low_index => 80, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_126, dout => sliced_v211_243, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_246_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_246_inst_req_0;
      slice_246_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_246_inst_req_1;
      slice_246_inst_ack_1<= update_ack(0);
      slice_246_inst: SliceSplitProtocol generic map(name => "slice_246_inst", in_data_width => 256, high_index => 79, low_index => 64, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_126, dout => sliced_v212_247, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_250_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_250_inst_req_0;
      slice_250_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_250_inst_req_1;
      slice_250_inst_ack_1<= update_ack(0);
      slice_250_inst: SliceSplitProtocol generic map(name => "slice_250_inst", in_data_width => 256, high_index => 63, low_index => 48, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_126, dout => sliced_v213_251, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_254_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_254_inst_req_0;
      slice_254_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_254_inst_req_1;
      slice_254_inst_ack_1<= update_ack(0);
      slice_254_inst: SliceSplitProtocol generic map(name => "slice_254_inst", in_data_width => 256, high_index => 47, low_index => 32, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_126, dout => sliced_v214_255, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_258_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_258_inst_req_0;
      slice_258_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_258_inst_req_1;
      slice_258_inst_ack_1<= update_ack(0);
      slice_258_inst: SliceSplitProtocol generic map(name => "slice_258_inst", in_data_width => 256, high_index => 31, low_index => 16, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_126, dout => sliced_v215_259, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_262_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_262_inst_req_0;
      slice_262_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_262_inst_req_1;
      slice_262_inst_ack_1<= update_ack(0);
      slice_262_inst: SliceSplitProtocol generic map(name => "slice_262_inst", in_data_width => 256, high_index => 15, low_index => 0, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c2_126, dout => sliced_v216_263, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_266_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_266_inst_req_0;
      slice_266_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_266_inst_req_1;
      slice_266_inst_ack_1<= update_ack(0);
      slice_266_inst: SliceSplitProtocol generic map(name => "slice_266_inst", in_data_width => 256, high_index => 255, low_index => 240, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_130, dout => sliced_v31_267, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_270_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_270_inst_req_0;
      slice_270_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_270_inst_req_1;
      slice_270_inst_ack_1<= update_ack(0);
      slice_270_inst: SliceSplitProtocol generic map(name => "slice_270_inst", in_data_width => 256, high_index => 239, low_index => 224, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_130, dout => sliced_v32_271, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_274_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_274_inst_req_0;
      slice_274_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_274_inst_req_1;
      slice_274_inst_ack_1<= update_ack(0);
      slice_274_inst: SliceSplitProtocol generic map(name => "slice_274_inst", in_data_width => 256, high_index => 223, low_index => 208, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_130, dout => sliced_v33_275, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_278_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_278_inst_req_0;
      slice_278_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_278_inst_req_1;
      slice_278_inst_ack_1<= update_ack(0);
      slice_278_inst: SliceSplitProtocol generic map(name => "slice_278_inst", in_data_width => 256, high_index => 207, low_index => 192, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_130, dout => sliced_v34_279, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_282_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_282_inst_req_0;
      slice_282_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_282_inst_req_1;
      slice_282_inst_ack_1<= update_ack(0);
      slice_282_inst: SliceSplitProtocol generic map(name => "slice_282_inst", in_data_width => 256, high_index => 191, low_index => 176, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_130, dout => sliced_v35_283, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_286_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_286_inst_req_0;
      slice_286_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_286_inst_req_1;
      slice_286_inst_ack_1<= update_ack(0);
      slice_286_inst: SliceSplitProtocol generic map(name => "slice_286_inst", in_data_width => 256, high_index => 175, low_index => 160, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_130, dout => sliced_v36_287, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_290_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_290_inst_req_0;
      slice_290_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_290_inst_req_1;
      slice_290_inst_ack_1<= update_ack(0);
      slice_290_inst: SliceSplitProtocol generic map(name => "slice_290_inst", in_data_width => 256, high_index => 159, low_index => 144, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_130, dout => sliced_v37_291, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_294_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_294_inst_req_0;
      slice_294_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_294_inst_req_1;
      slice_294_inst_ack_1<= update_ack(0);
      slice_294_inst: SliceSplitProtocol generic map(name => "slice_294_inst", in_data_width => 256, high_index => 143, low_index => 128, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_130, dout => sliced_v38_295, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_298_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_298_inst_req_0;
      slice_298_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_298_inst_req_1;
      slice_298_inst_ack_1<= update_ack(0);
      slice_298_inst: SliceSplitProtocol generic map(name => "slice_298_inst", in_data_width => 256, high_index => 127, low_index => 112, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_130, dout => sliced_v39_299, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_302_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_302_inst_req_0;
      slice_302_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_302_inst_req_1;
      slice_302_inst_ack_1<= update_ack(0);
      slice_302_inst: SliceSplitProtocol generic map(name => "slice_302_inst", in_data_width => 256, high_index => 111, low_index => 96, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_130, dout => sliced_v310_303, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_306_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_306_inst_req_0;
      slice_306_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_306_inst_req_1;
      slice_306_inst_ack_1<= update_ack(0);
      slice_306_inst: SliceSplitProtocol generic map(name => "slice_306_inst", in_data_width => 256, high_index => 95, low_index => 80, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_130, dout => sliced_v311_307, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_310_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_310_inst_req_0;
      slice_310_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_310_inst_req_1;
      slice_310_inst_ack_1<= update_ack(0);
      slice_310_inst: SliceSplitProtocol generic map(name => "slice_310_inst", in_data_width => 256, high_index => 79, low_index => 64, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_130, dout => sliced_v312_311, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_314_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_314_inst_req_0;
      slice_314_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_314_inst_req_1;
      slice_314_inst_ack_1<= update_ack(0);
      slice_314_inst: SliceSplitProtocol generic map(name => "slice_314_inst", in_data_width => 256, high_index => 63, low_index => 48, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_130, dout => sliced_v313_315, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_318_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_318_inst_req_0;
      slice_318_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_318_inst_req_1;
      slice_318_inst_ack_1<= update_ack(0);
      slice_318_inst: SliceSplitProtocol generic map(name => "slice_318_inst", in_data_width => 256, high_index => 47, low_index => 32, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_130, dout => sliced_v314_319, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_322_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_322_inst_req_0;
      slice_322_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_322_inst_req_1;
      slice_322_inst_ack_1<= update_ack(0);
      slice_322_inst: SliceSplitProtocol generic map(name => "slice_322_inst", in_data_width => 256, high_index => 31, low_index => 16, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_130, dout => sliced_v315_323, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_326_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_326_inst_req_0;
      slice_326_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_326_inst_req_1;
      slice_326_inst_ack_1<= update_ack(0);
      slice_326_inst: SliceSplitProtocol generic map(name => "slice_326_inst", in_data_width => 256, high_index => 15, low_index => 0, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c3_130, dout => sliced_v316_327, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_330_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_330_inst_req_0;
      slice_330_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_330_inst_req_1;
      slice_330_inst_ack_1<= update_ack(0);
      slice_330_inst: SliceSplitProtocol generic map(name => "slice_330_inst", in_data_width => 256, high_index => 255, low_index => 240, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_134, dout => sliced_v41_331, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_334_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_334_inst_req_0;
      slice_334_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_334_inst_req_1;
      slice_334_inst_ack_1<= update_ack(0);
      slice_334_inst: SliceSplitProtocol generic map(name => "slice_334_inst", in_data_width => 256, high_index => 239, low_index => 224, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_134, dout => sliced_v42_335, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_338_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_338_inst_req_0;
      slice_338_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_338_inst_req_1;
      slice_338_inst_ack_1<= update_ack(0);
      slice_338_inst: SliceSplitProtocol generic map(name => "slice_338_inst", in_data_width => 256, high_index => 223, low_index => 208, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_134, dout => sliced_v43_339, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_342_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_342_inst_req_0;
      slice_342_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_342_inst_req_1;
      slice_342_inst_ack_1<= update_ack(0);
      slice_342_inst: SliceSplitProtocol generic map(name => "slice_342_inst", in_data_width => 256, high_index => 207, low_index => 192, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_134, dout => sliced_v44_343, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_346_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_346_inst_req_0;
      slice_346_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_346_inst_req_1;
      slice_346_inst_ack_1<= update_ack(0);
      slice_346_inst: SliceSplitProtocol generic map(name => "slice_346_inst", in_data_width => 256, high_index => 191, low_index => 176, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_134, dout => sliced_v45_347, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_350_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_350_inst_req_0;
      slice_350_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_350_inst_req_1;
      slice_350_inst_ack_1<= update_ack(0);
      slice_350_inst: SliceSplitProtocol generic map(name => "slice_350_inst", in_data_width => 256, high_index => 175, low_index => 160, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_134, dout => sliced_v46_351, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_354_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_354_inst_req_0;
      slice_354_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_354_inst_req_1;
      slice_354_inst_ack_1<= update_ack(0);
      slice_354_inst: SliceSplitProtocol generic map(name => "slice_354_inst", in_data_width => 256, high_index => 159, low_index => 144, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_134, dout => sliced_v47_355, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_358_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_358_inst_req_0;
      slice_358_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_358_inst_req_1;
      slice_358_inst_ack_1<= update_ack(0);
      slice_358_inst: SliceSplitProtocol generic map(name => "slice_358_inst", in_data_width => 256, high_index => 143, low_index => 128, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_134, dout => sliced_v48_359, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_362_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_362_inst_req_0;
      slice_362_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_362_inst_req_1;
      slice_362_inst_ack_1<= update_ack(0);
      slice_362_inst: SliceSplitProtocol generic map(name => "slice_362_inst", in_data_width => 256, high_index => 127, low_index => 112, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_134, dout => sliced_v49_363, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_366_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_366_inst_req_0;
      slice_366_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_366_inst_req_1;
      slice_366_inst_ack_1<= update_ack(0);
      slice_366_inst: SliceSplitProtocol generic map(name => "slice_366_inst", in_data_width => 256, high_index => 111, low_index => 96, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_134, dout => sliced_v410_367, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_370_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_370_inst_req_0;
      slice_370_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_370_inst_req_1;
      slice_370_inst_ack_1<= update_ack(0);
      slice_370_inst: SliceSplitProtocol generic map(name => "slice_370_inst", in_data_width => 256, high_index => 95, low_index => 80, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_134, dout => sliced_v411_371, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_374_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_374_inst_req_0;
      slice_374_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_374_inst_req_1;
      slice_374_inst_ack_1<= update_ack(0);
      slice_374_inst: SliceSplitProtocol generic map(name => "slice_374_inst", in_data_width => 256, high_index => 79, low_index => 64, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_134, dout => sliced_v412_375, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_378_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_378_inst_req_0;
      slice_378_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_378_inst_req_1;
      slice_378_inst_ack_1<= update_ack(0);
      slice_378_inst: SliceSplitProtocol generic map(name => "slice_378_inst", in_data_width => 256, high_index => 63, low_index => 48, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_134, dout => sliced_v413_379, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_382_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_382_inst_req_0;
      slice_382_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_382_inst_req_1;
      slice_382_inst_ack_1<= update_ack(0);
      slice_382_inst: SliceSplitProtocol generic map(name => "slice_382_inst", in_data_width => 256, high_index => 47, low_index => 32, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_134, dout => sliced_v414_383, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_386_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_386_inst_req_0;
      slice_386_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_386_inst_req_1;
      slice_386_inst_ack_1<= update_ack(0);
      slice_386_inst: SliceSplitProtocol generic map(name => "slice_386_inst", in_data_width => 256, high_index => 31, low_index => 16, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_134, dout => sliced_v415_387, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_390_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_390_inst_req_0;
      slice_390_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_390_inst_req_1;
      slice_390_inst_ack_1<= update_ack(0);
      slice_390_inst: SliceSplitProtocol generic map(name => "slice_390_inst", in_data_width => 256, high_index => 15, low_index => 0, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => c4_134, dout => sliced_v416_391, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    W_myptr5_1040_delayed_8_0_1040_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_myptr5_1040_delayed_8_0_1040_inst_req_0;
      W_myptr5_1040_delayed_8_0_1040_inst_ack_0<= wack(0);
      rreq(0) <= W_myptr5_1040_delayed_8_0_1040_inst_req_1;
      W_myptr5_1040_delayed_8_0_1040_inst_ack_1<= rack(0);
      W_myptr5_1040_delayed_8_0_1040_inst : InterlockBuffer generic map ( -- 
        name => "W_myptr5_1040_delayed_8_0_1040_inst",
        buffer_size => 8,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => myptr5_1039,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => myptr5_1040_delayed_8_0_1042,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_myptr6_1063_delayed_8_0_1066_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_myptr6_1063_delayed_8_0_1066_inst_req_0;
      W_myptr6_1063_delayed_8_0_1066_inst_ack_0<= wack(0);
      rreq(0) <= W_myptr6_1063_delayed_8_0_1066_inst_req_1;
      W_myptr6_1063_delayed_8_0_1066_inst_ack_1<= rack(0);
      W_myptr6_1063_delayed_8_0_1066_inst : InterlockBuffer generic map ( -- 
        name => "W_myptr6_1063_delayed_8_0_1066_inst",
        buffer_size => 8,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => myptr6_1065,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => myptr6_1063_delayed_8_0_1068,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_myptr7_1086_delayed_8_0_1092_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_myptr7_1086_delayed_8_0_1092_inst_req_0;
      W_myptr7_1086_delayed_8_0_1092_inst_ack_0<= wack(0);
      rreq(0) <= W_myptr7_1086_delayed_8_0_1092_inst_req_1;
      W_myptr7_1086_delayed_8_0_1092_inst_ack_1<= rack(0);
      W_myptr7_1086_delayed_8_0_1092_inst : InterlockBuffer generic map ( -- 
        name => "W_myptr7_1086_delayed_8_0_1092_inst",
        buffer_size => 8,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => myptr7_1091,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => myptr7_1086_delayed_8_0_1094,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_myptr8_1109_delayed_8_0_1118_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_myptr8_1109_delayed_8_0_1118_inst_req_0;
      W_myptr8_1109_delayed_8_0_1118_inst_ack_0<= wack(0);
      rreq(0) <= W_myptr8_1109_delayed_8_0_1118_inst_req_1;
      W_myptr8_1109_delayed_8_0_1118_inst_ack_1<= rack(0);
      W_myptr8_1109_delayed_8_0_1118_inst : InterlockBuffer generic map ( -- 
        name => "W_myptr8_1109_delayed_8_0_1118_inst",
        buffer_size => 8,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => myptr8_1117,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => myptr8_1109_delayed_8_0_1120,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1038_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1038_final_reg_req_0;
      addr_of_1038_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1038_final_reg_req_1;
      addr_of_1038_final_reg_ack_1<= rack(0);
      addr_of_1038_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1038_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1037_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => myptr5_1039,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_103_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_103_final_reg_req_0;
      addr_of_103_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_103_final_reg_req_1;
      addr_of_103_final_reg_ack_1<= rack(0);
      addr_of_103_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_103_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_102_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => myptr2_104,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1064_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1064_final_reg_req_0;
      addr_of_1064_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1064_final_reg_req_1;
      addr_of_1064_final_reg_ack_1<= rack(0);
      addr_of_1064_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1064_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1063_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => myptr6_1065,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1090_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1090_final_reg_req_0;
      addr_of_1090_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1090_final_reg_req_1;
      addr_of_1090_final_reg_ack_1<= rack(0);
      addr_of_1090_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1090_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1089_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => myptr7_1091,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_110_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_110_final_reg_req_0;
      addr_of_110_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_110_final_reg_req_1;
      addr_of_110_final_reg_ack_1<= rack(0);
      addr_of_110_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_110_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_109_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => myptr3_111,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1116_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1116_final_reg_req_0;
      addr_of_1116_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1116_final_reg_req_1;
      addr_of_1116_final_reg_ack_1<= rack(0);
      addr_of_1116_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1116_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1115_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => myptr8_1117,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_117_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_117_final_reg_req_0;
      addr_of_117_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_117_final_reg_req_1;
      addr_of_117_final_reg_ack_1<= rack(0);
      addr_of_117_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_117_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_116_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => myptr4_118,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_96_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_96_final_reg_req_0;
      addr_of_96_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_96_final_reg_req_1;
      addr_of_96_final_reg_ack_1<= rack(0);
      addr_of_96_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_96_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_95_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => myptr1_97,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1046_inst
    process(out1_672) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out1_672(15 downto 0);
      type_cast_1046_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1048_inst
    process(out2_696) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out2_696(15 downto 0);
      type_cast_1048_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1051_inst
    process(out3_720) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out3_720(15 downto 0);
      type_cast_1051_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1053_inst
    process(out4_744) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out4_744(15 downto 0);
      type_cast_1053_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1072_inst
    process(out5_768) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out5_768(15 downto 0);
      type_cast_1072_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1074_inst
    process(out6_792) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out6_792(15 downto 0);
      type_cast_1074_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1077_inst
    process(out7_816) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out7_816(15 downto 0);
      type_cast_1077_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1079_inst
    process(out8_840) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out8_840(15 downto 0);
      type_cast_1079_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1098_inst
    process(out9_864) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out9_864(15 downto 0);
      type_cast_1098_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1100_inst
    process(out10_888) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out10_888(15 downto 0);
      type_cast_1100_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1103_inst
    process(out11_912) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out11_912(15 downto 0);
      type_cast_1103_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1105_inst
    process(out12_936) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out12_936(15 downto 0);
      type_cast_1105_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1124_inst
    process(out13_960) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out13_960(15 downto 0);
      type_cast_1124_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1126_inst
    process(out14_984) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out14_984(15 downto 0);
      type_cast_1126_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1129_inst
    process(out15_1008) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out15_1008(15 downto 0);
      type_cast_1129_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1131_inst
    process(out16_1032) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := out16_1032(15 downto 0);
      type_cast_1131_wire <= tmp_var; -- 
    end process;
    type_cast_1137_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1137_inst_req_0;
      type_cast_1137_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1137_inst_req_1;
      type_cast_1137_inst_ack_1<= rack(0);
      type_cast_1137_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1137_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => out1_672,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => output_buffer,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_395_inst
    process(sliced_v11_139) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v11_139(15 downto 0);
      a11_396 <= tmp_var; -- 
    end process;
    -- interlock type_cast_399_inst
    process(sliced_v12_143) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v12_143(15 downto 0);
      a12_400 <= tmp_var; -- 
    end process;
    -- interlock type_cast_403_inst
    process(sliced_v13_147) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v13_147(15 downto 0);
      a13_404 <= tmp_var; -- 
    end process;
    -- interlock type_cast_407_inst
    process(sliced_v14_151) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v14_151(15 downto 0);
      a14_408 <= tmp_var; -- 
    end process;
    -- interlock type_cast_411_inst
    process(sliced_v15_155) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v15_155(15 downto 0);
      a15_412 <= tmp_var; -- 
    end process;
    -- interlock type_cast_415_inst
    process(sliced_v16_159) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v16_159(15 downto 0);
      a16_416 <= tmp_var; -- 
    end process;
    -- interlock type_cast_419_inst
    process(sliced_v17_163) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v17_163(15 downto 0);
      a17_420 <= tmp_var; -- 
    end process;
    -- interlock type_cast_423_inst
    process(sliced_v18_167) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v18_167(15 downto 0);
      a18_424 <= tmp_var; -- 
    end process;
    -- interlock type_cast_427_inst
    process(sliced_v19_171) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v19_171(15 downto 0);
      a19_428 <= tmp_var; -- 
    end process;
    -- interlock type_cast_431_inst
    process(sliced_v110_175) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v110_175(15 downto 0);
      a110_432 <= tmp_var; -- 
    end process;
    -- interlock type_cast_435_inst
    process(sliced_v111_179) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v111_179(15 downto 0);
      a111_436 <= tmp_var; -- 
    end process;
    -- interlock type_cast_439_inst
    process(sliced_v112_183) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v112_183(15 downto 0);
      a112_440 <= tmp_var; -- 
    end process;
    -- interlock type_cast_443_inst
    process(sliced_v113_187) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v113_187(15 downto 0);
      a113_444 <= tmp_var; -- 
    end process;
    -- interlock type_cast_447_inst
    process(sliced_v114_191) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v114_191(15 downto 0);
      a114_448 <= tmp_var; -- 
    end process;
    -- interlock type_cast_451_inst
    process(sliced_v115_195) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v115_195(15 downto 0);
      a115_452 <= tmp_var; -- 
    end process;
    -- interlock type_cast_455_inst
    process(sliced_v116_199) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v116_199(15 downto 0);
      a116_456 <= tmp_var; -- 
    end process;
    -- interlock type_cast_459_inst
    process(sliced_v21_203) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v21_203(15 downto 0);
      a21_460 <= tmp_var; -- 
    end process;
    -- interlock type_cast_463_inst
    process(sliced_v22_207) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v22_207(15 downto 0);
      a22_464 <= tmp_var; -- 
    end process;
    -- interlock type_cast_467_inst
    process(sliced_v23_211) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v23_211(15 downto 0);
      a23_468 <= tmp_var; -- 
    end process;
    -- interlock type_cast_471_inst
    process(sliced_v24_215) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v24_215(15 downto 0);
      a24_472 <= tmp_var; -- 
    end process;
    -- interlock type_cast_475_inst
    process(sliced_v25_219) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v25_219(15 downto 0);
      a25_476 <= tmp_var; -- 
    end process;
    -- interlock type_cast_479_inst
    process(sliced_v26_223) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v26_223(15 downto 0);
      a26_480 <= tmp_var; -- 
    end process;
    -- interlock type_cast_483_inst
    process(sliced_v27_227) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v27_227(15 downto 0);
      a27_484 <= tmp_var; -- 
    end process;
    -- interlock type_cast_487_inst
    process(sliced_v28_231) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v28_231(15 downto 0);
      a28_488 <= tmp_var; -- 
    end process;
    -- interlock type_cast_491_inst
    process(sliced_v29_235) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v29_235(15 downto 0);
      a29_492 <= tmp_var; -- 
    end process;
    -- interlock type_cast_495_inst
    process(sliced_v210_239) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v210_239(15 downto 0);
      a210_496 <= tmp_var; -- 
    end process;
    -- interlock type_cast_499_inst
    process(sliced_v211_243) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v211_243(15 downto 0);
      a211_500 <= tmp_var; -- 
    end process;
    -- interlock type_cast_503_inst
    process(sliced_v212_247) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v212_247(15 downto 0);
      a212_504 <= tmp_var; -- 
    end process;
    -- interlock type_cast_507_inst
    process(sliced_v213_251) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v213_251(15 downto 0);
      a213_508 <= tmp_var; -- 
    end process;
    -- interlock type_cast_511_inst
    process(sliced_v214_255) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v214_255(15 downto 0);
      a214_512 <= tmp_var; -- 
    end process;
    -- interlock type_cast_515_inst
    process(sliced_v215_259) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v215_259(15 downto 0);
      a215_516 <= tmp_var; -- 
    end process;
    -- interlock type_cast_519_inst
    process(sliced_v216_263) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v216_263(15 downto 0);
      a216_520 <= tmp_var; -- 
    end process;
    -- interlock type_cast_523_inst
    process(sliced_v31_267) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v31_267(15 downto 0);
      a31_524 <= tmp_var; -- 
    end process;
    -- interlock type_cast_527_inst
    process(sliced_v32_271) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v32_271(15 downto 0);
      a32_528 <= tmp_var; -- 
    end process;
    -- interlock type_cast_531_inst
    process(sliced_v33_275) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v33_275(15 downto 0);
      a33_532 <= tmp_var; -- 
    end process;
    -- interlock type_cast_535_inst
    process(sliced_v34_279) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v34_279(15 downto 0);
      a34_536 <= tmp_var; -- 
    end process;
    -- interlock type_cast_539_inst
    process(sliced_v35_283) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v35_283(15 downto 0);
      a35_540 <= tmp_var; -- 
    end process;
    -- interlock type_cast_543_inst
    process(sliced_v36_287) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v36_287(15 downto 0);
      a36_544 <= tmp_var; -- 
    end process;
    -- interlock type_cast_547_inst
    process(sliced_v37_291) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v37_291(15 downto 0);
      a37_548 <= tmp_var; -- 
    end process;
    -- interlock type_cast_551_inst
    process(sliced_v38_295) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v38_295(15 downto 0);
      a38_552 <= tmp_var; -- 
    end process;
    -- interlock type_cast_555_inst
    process(sliced_v39_299) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v39_299(15 downto 0);
      a39_556 <= tmp_var; -- 
    end process;
    -- interlock type_cast_559_inst
    process(sliced_v310_303) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v310_303(15 downto 0);
      a310_560 <= tmp_var; -- 
    end process;
    -- interlock type_cast_563_inst
    process(sliced_v311_307) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v311_307(15 downto 0);
      a311_564 <= tmp_var; -- 
    end process;
    -- interlock type_cast_567_inst
    process(sliced_v312_311) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v312_311(15 downto 0);
      a312_568 <= tmp_var; -- 
    end process;
    -- interlock type_cast_571_inst
    process(sliced_v313_315) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v313_315(15 downto 0);
      a313_572 <= tmp_var; -- 
    end process;
    -- interlock type_cast_575_inst
    process(sliced_v314_319) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v314_319(15 downto 0);
      a314_576 <= tmp_var; -- 
    end process;
    -- interlock type_cast_579_inst
    process(sliced_v315_323) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v315_323(15 downto 0);
      a315_580 <= tmp_var; -- 
    end process;
    -- interlock type_cast_583_inst
    process(sliced_v316_327) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v316_327(15 downto 0);
      a316_584 <= tmp_var; -- 
    end process;
    -- interlock type_cast_587_inst
    process(sliced_v41_331) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v41_331(15 downto 0);
      a41_588 <= tmp_var; -- 
    end process;
    -- interlock type_cast_591_inst
    process(sliced_v42_335) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v42_335(15 downto 0);
      a42_592 <= tmp_var; -- 
    end process;
    -- interlock type_cast_595_inst
    process(sliced_v43_339) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v43_339(15 downto 0);
      a43_596 <= tmp_var; -- 
    end process;
    -- interlock type_cast_599_inst
    process(sliced_v44_343) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v44_343(15 downto 0);
      a44_600 <= tmp_var; -- 
    end process;
    -- interlock type_cast_603_inst
    process(sliced_v45_347) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v45_347(15 downto 0);
      a45_604 <= tmp_var; -- 
    end process;
    -- interlock type_cast_607_inst
    process(sliced_v46_351) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v46_351(15 downto 0);
      a46_608 <= tmp_var; -- 
    end process;
    -- interlock type_cast_611_inst
    process(sliced_v47_355) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v47_355(15 downto 0);
      a47_612 <= tmp_var; -- 
    end process;
    -- interlock type_cast_615_inst
    process(sliced_v48_359) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v48_359(15 downto 0);
      a48_616 <= tmp_var; -- 
    end process;
    -- interlock type_cast_619_inst
    process(sliced_v49_363) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v49_363(15 downto 0);
      a49_620 <= tmp_var; -- 
    end process;
    -- interlock type_cast_623_inst
    process(sliced_v410_367) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v410_367(15 downto 0);
      a410_624 <= tmp_var; -- 
    end process;
    -- interlock type_cast_627_inst
    process(sliced_v411_371) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v411_371(15 downto 0);
      a411_628 <= tmp_var; -- 
    end process;
    -- interlock type_cast_631_inst
    process(sliced_v412_375) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v412_375(15 downto 0);
      a412_632 <= tmp_var; -- 
    end process;
    -- interlock type_cast_635_inst
    process(sliced_v413_379) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v413_379(15 downto 0);
      a413_636 <= tmp_var; -- 
    end process;
    -- interlock type_cast_639_inst
    process(sliced_v414_383) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v414_383(15 downto 0);
      a414_640 <= tmp_var; -- 
    end process;
    -- interlock type_cast_643_inst
    process(sliced_v415_387) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v415_387(15 downto 0);
      a415_644 <= tmp_var; -- 
    end process;
    -- interlock type_cast_647_inst
    process(sliced_v416_391) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := sliced_v416_391(15 downto 0);
      a416_648 <= tmp_var; -- 
    end process;
    -- equivalence array_obj_ref_102_index_1_rename
    process(R_addr2_101_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr2_101_resized;
      ov(13 downto 0) := iv;
      R_addr2_101_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_102_index_1_resize
    process(addr2_buffer) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := addr2_buffer;
      ov := iv(13 downto 0);
      R_addr2_101_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_102_root_address_inst
    process(array_obj_ref_102_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_102_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_102_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1037_index_1_rename
    process(R_addr_1036_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr_1036_resized;
      ov(13 downto 0) := iv;
      R_addr_1036_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1037_index_1_resize
    process(addr_buffer) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := addr_buffer;
      ov := iv(13 downto 0);
      R_addr_1036_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1037_root_address_inst
    process(array_obj_ref_1037_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1037_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1037_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1063_index_1_rename
    process(ADD_u32_u32_1062_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ADD_u32_u32_1062_resized;
      ov(13 downto 0) := iv;
      ADD_u32_u32_1062_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1063_index_1_resize
    process(ADD_u32_u32_1062_wire) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ADD_u32_u32_1062_wire;
      ov := iv(13 downto 0);
      ADD_u32_u32_1062_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1063_root_address_inst
    process(array_obj_ref_1063_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1063_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1063_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1089_index_1_rename
    process(ADD_u32_u32_1088_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ADD_u32_u32_1088_resized;
      ov(13 downto 0) := iv;
      ADD_u32_u32_1088_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1089_index_1_resize
    process(ADD_u32_u32_1088_wire) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ADD_u32_u32_1088_wire;
      ov := iv(13 downto 0);
      ADD_u32_u32_1088_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1089_root_address_inst
    process(array_obj_ref_1089_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1089_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1089_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_109_index_1_rename
    process(R_addr3_108_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr3_108_resized;
      ov(13 downto 0) := iv;
      R_addr3_108_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_109_index_1_resize
    process(addr3_buffer) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := addr3_buffer;
      ov := iv(13 downto 0);
      R_addr3_108_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_109_root_address_inst
    process(array_obj_ref_109_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_109_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_109_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1115_index_1_rename
    process(ADD_u32_u32_1114_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ADD_u32_u32_1114_resized;
      ov(13 downto 0) := iv;
      ADD_u32_u32_1114_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1115_index_1_resize
    process(ADD_u32_u32_1114_wire) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ADD_u32_u32_1114_wire;
      ov := iv(13 downto 0);
      ADD_u32_u32_1114_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1115_root_address_inst
    process(array_obj_ref_1115_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1115_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1115_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_116_index_1_rename
    process(R_addr4_115_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr4_115_resized;
      ov(13 downto 0) := iv;
      R_addr4_115_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_116_index_1_resize
    process(addr4_buffer) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := addr4_buffer;
      ov := iv(13 downto 0);
      R_addr4_115_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_116_root_address_inst
    process(array_obj_ref_116_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_116_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_116_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_95_index_1_rename
    process(R_addr1_94_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_addr1_94_resized;
      ov(13 downto 0) := iv;
      R_addr1_94_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_95_index_1_resize
    process(addr1_buffer) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := addr1_buffer;
      ov := iv(13 downto 0);
      R_addr1_94_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_95_root_address_inst
    process(array_obj_ref_95_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_95_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_95_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1044_addr_0
    process(ptr_deref_1044_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1044_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1044_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1044_base_resize
    process(myptr5_1040_delayed_8_0_1042) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := myptr5_1040_delayed_8_0_1042;
      ov := iv(13 downto 0);
      ptr_deref_1044_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1044_gather_scatter
    process(CONCAT_u32_u64_1055_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := CONCAT_u32_u64_1055_wire;
      ov(63 downto 0) := iv;
      ptr_deref_1044_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1044_root_address_inst
    process(ptr_deref_1044_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1044_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1044_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1070_addr_0
    process(ptr_deref_1070_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1070_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1070_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1070_base_resize
    process(myptr6_1063_delayed_8_0_1068) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := myptr6_1063_delayed_8_0_1068;
      ov := iv(13 downto 0);
      ptr_deref_1070_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1070_gather_scatter
    process(CONCAT_u32_u64_1081_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := CONCAT_u32_u64_1081_wire;
      ov(63 downto 0) := iv;
      ptr_deref_1070_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1070_root_address_inst
    process(ptr_deref_1070_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1070_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1070_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1096_addr_0
    process(ptr_deref_1096_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1096_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1096_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1096_base_resize
    process(myptr7_1086_delayed_8_0_1094) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := myptr7_1086_delayed_8_0_1094;
      ov := iv(13 downto 0);
      ptr_deref_1096_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1096_gather_scatter
    process(CONCAT_u32_u64_1107_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := CONCAT_u32_u64_1107_wire;
      ov(63 downto 0) := iv;
      ptr_deref_1096_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1096_root_address_inst
    process(ptr_deref_1096_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1096_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1096_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1122_addr_0
    process(ptr_deref_1122_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1122_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1122_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1122_base_resize
    process(myptr8_1109_delayed_8_0_1120) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := myptr8_1109_delayed_8_0_1120;
      ov := iv(13 downto 0);
      ptr_deref_1122_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1122_gather_scatter
    process(CONCAT_u32_u64_1133_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := CONCAT_u32_u64_1133_wire;
      ov(63 downto 0) := iv;
      ptr_deref_1122_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1122_root_address_inst
    process(ptr_deref_1122_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1122_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1122_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_121_addr_0
    process(ptr_deref_121_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_121_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_121_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_121_base_resize
    process(myptr1_97) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := myptr1_97;
      ov := iv(13 downto 0);
      ptr_deref_121_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_121_gather_scatter
    process(ptr_deref_121_data_0) --
      variable iv : std_logic_vector(255 downto 0);
      variable ov : std_logic_vector(255 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_121_data_0;
      ov(255 downto 0) := iv;
      c1_122 <= ov(255 downto 0);
      --
    end process;
    -- equivalence ptr_deref_121_root_address_inst
    process(ptr_deref_121_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_121_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_121_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_125_addr_0
    process(ptr_deref_125_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_125_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_125_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_125_base_resize
    process(myptr2_104) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := myptr2_104;
      ov := iv(13 downto 0);
      ptr_deref_125_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_125_gather_scatter
    process(ptr_deref_125_data_0) --
      variable iv : std_logic_vector(255 downto 0);
      variable ov : std_logic_vector(255 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_125_data_0;
      ov(255 downto 0) := iv;
      c2_126 <= ov(255 downto 0);
      --
    end process;
    -- equivalence ptr_deref_125_root_address_inst
    process(ptr_deref_125_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_125_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_125_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_129_addr_0
    process(ptr_deref_129_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_129_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_129_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_129_base_resize
    process(myptr3_111) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := myptr3_111;
      ov := iv(13 downto 0);
      ptr_deref_129_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_129_gather_scatter
    process(ptr_deref_129_data_0) --
      variable iv : std_logic_vector(255 downto 0);
      variable ov : std_logic_vector(255 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_129_data_0;
      ov(255 downto 0) := iv;
      c3_130 <= ov(255 downto 0);
      --
    end process;
    -- equivalence ptr_deref_129_root_address_inst
    process(ptr_deref_129_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_129_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_129_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_133_addr_0
    process(ptr_deref_133_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_133_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_133_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_133_base_resize
    process(myptr4_118) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := myptr4_118;
      ov := iv(13 downto 0);
      ptr_deref_133_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_133_gather_scatter
    process(ptr_deref_133_data_0) --
      variable iv : std_logic_vector(255 downto 0);
      variable ov : std_logic_vector(255 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_133_data_0;
      ov(255 downto 0) := iv;
      c4_134 <= ov(255 downto 0);
      --
    end process;
    -- equivalence ptr_deref_133_root_address_inst
    process(ptr_deref_133_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_133_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_133_root_address <= ov(13 downto 0);
      --
    end process;
    -- binary operator ADD_u32_u32_1062_inst
    process(addr_buffer) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(addr_buffer, konst_1061_wire_constant, tmp_var);
      ADD_u32_u32_1062_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1088_inst
    process(addr_buffer) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(addr_buffer, konst_1087_wire_constant, tmp_var);
      ADD_u32_u32_1088_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1114_inst
    process(addr_buffer) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(addr_buffer, konst_1113_wire_constant, tmp_var);
      ADD_u32_u32_1114_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u16_u32_1049_inst
    process(type_cast_1046_wire, type_cast_1048_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_1046_wire, type_cast_1048_wire, tmp_var);
      CONCAT_u16_u32_1049_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u16_u32_1054_inst
    process(type_cast_1051_wire, type_cast_1053_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_1051_wire, type_cast_1053_wire, tmp_var);
      CONCAT_u16_u32_1054_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u16_u32_1075_inst
    process(type_cast_1072_wire, type_cast_1074_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_1072_wire, type_cast_1074_wire, tmp_var);
      CONCAT_u16_u32_1075_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u16_u32_1080_inst
    process(type_cast_1077_wire, type_cast_1079_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_1077_wire, type_cast_1079_wire, tmp_var);
      CONCAT_u16_u32_1080_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u16_u32_1101_inst
    process(type_cast_1098_wire, type_cast_1100_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_1098_wire, type_cast_1100_wire, tmp_var);
      CONCAT_u16_u32_1101_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u16_u32_1106_inst
    process(type_cast_1103_wire, type_cast_1105_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_1103_wire, type_cast_1105_wire, tmp_var);
      CONCAT_u16_u32_1106_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u16_u32_1127_inst
    process(type_cast_1124_wire, type_cast_1126_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_1124_wire, type_cast_1126_wire, tmp_var);
      CONCAT_u16_u32_1127_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u16_u32_1132_inst
    process(type_cast_1129_wire, type_cast_1131_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_1129_wire, type_cast_1131_wire, tmp_var);
      CONCAT_u16_u32_1132_wire <= tmp_var; --
    end process;
    -- shared split operator group (11) : CONCAT_u32_u64_1055_inst 
    ApConcat_group_11: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= CONCAT_u16_u32_1049_wire & CONCAT_u16_u32_1054_wire;
      CONCAT_u32_u64_1055_wire <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u32_u64_1055_inst_req_0;
      CONCAT_u32_u64_1055_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u32_u64_1055_inst_req_1;
      CONCAT_u32_u64_1055_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_11_gI: SplitGuardInterface generic map(name => "ApConcat_group_11_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_11",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 11
    -- shared split operator group (12) : CONCAT_u32_u64_1081_inst 
    ApConcat_group_12: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= CONCAT_u16_u32_1075_wire & CONCAT_u16_u32_1080_wire;
      CONCAT_u32_u64_1081_wire <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u32_u64_1081_inst_req_0;
      CONCAT_u32_u64_1081_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u32_u64_1081_inst_req_1;
      CONCAT_u32_u64_1081_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_12_gI: SplitGuardInterface generic map(name => "ApConcat_group_12_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_12",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 12
    -- shared split operator group (13) : CONCAT_u32_u64_1107_inst 
    ApConcat_group_13: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= CONCAT_u16_u32_1101_wire & CONCAT_u16_u32_1106_wire;
      CONCAT_u32_u64_1107_wire <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u32_u64_1107_inst_req_0;
      CONCAT_u32_u64_1107_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u32_u64_1107_inst_req_1;
      CONCAT_u32_u64_1107_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_13_gI: SplitGuardInterface generic map(name => "ApConcat_group_13_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_13",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 13
    -- shared split operator group (14) : CONCAT_u32_u64_1133_inst 
    ApConcat_group_14: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= CONCAT_u16_u32_1127_wire & CONCAT_u16_u32_1132_wire;
      CONCAT_u32_u64_1133_wire <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u32_u64_1133_inst_req_0;
      CONCAT_u32_u64_1133_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u32_u64_1133_inst_req_1;
      CONCAT_u32_u64_1133_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_14_gI: SplitGuardInterface generic map(name => "ApConcat_group_14_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_14",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 14
    -- binary operator SGT_i16_u1_1004_inst
    process(t151_992, t152_1000) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t151_992, t152_1000, tmp_var);
      SGT_i16_u1_1004_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_1012_inst
    process(a116_456, a216_520) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a116_456, a216_520, tmp_var);
      SGT_i16_u1_1012_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_1020_inst
    process(a316_584, a416_648) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a316_584, a416_648, tmp_var);
      SGT_i16_u1_1020_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_1028_inst
    process(t161_1016, t162_1024) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t161_1016, t162_1024, tmp_var);
      SGT_i16_u1_1028_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_652_inst
    process(a11_396, a21_460) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a11_396, a21_460, tmp_var);
      SGT_i16_u1_652_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_660_inst
    process(a31_524, a41_588) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a31_524, a41_588, tmp_var);
      SGT_i16_u1_660_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_668_inst
    process(t11_656, t12_664) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t11_656, t12_664, tmp_var);
      SGT_i16_u1_668_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_676_inst
    process(a12_400, a22_464) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a12_400, a22_464, tmp_var);
      SGT_i16_u1_676_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_684_inst
    process(a32_528, a42_592) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a32_528, a42_592, tmp_var);
      SGT_i16_u1_684_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_692_inst
    process(t21_680, t22_688) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t21_680, t22_688, tmp_var);
      SGT_i16_u1_692_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_700_inst
    process(a13_404, a23_468) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a13_404, a23_468, tmp_var);
      SGT_i16_u1_700_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_708_inst
    process(a33_532, a43_596) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a33_532, a43_596, tmp_var);
      SGT_i16_u1_708_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_716_inst
    process(t31_704, t32_712) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t31_704, t32_712, tmp_var);
      SGT_i16_u1_716_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_724_inst
    process(a14_408, a24_472) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a14_408, a24_472, tmp_var);
      SGT_i16_u1_724_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_732_inst
    process(a34_536, a44_600) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a34_536, a44_600, tmp_var);
      SGT_i16_u1_732_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_740_inst
    process(t41_728, t42_736) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t41_728, t42_736, tmp_var);
      SGT_i16_u1_740_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_748_inst
    process(a15_412, a25_476) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a15_412, a25_476, tmp_var);
      SGT_i16_u1_748_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_756_inst
    process(a35_540, a45_604) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a35_540, a45_604, tmp_var);
      SGT_i16_u1_756_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_764_inst
    process(t51_752, t52_760) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t51_752, t52_760, tmp_var);
      SGT_i16_u1_764_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_772_inst
    process(a16_416, a26_480) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a16_416, a26_480, tmp_var);
      SGT_i16_u1_772_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_780_inst
    process(a36_544, a46_608) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a36_544, a46_608, tmp_var);
      SGT_i16_u1_780_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_788_inst
    process(t61_776, t62_784) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t61_776, t62_784, tmp_var);
      SGT_i16_u1_788_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_796_inst
    process(a17_420, a27_484) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a17_420, a27_484, tmp_var);
      SGT_i16_u1_796_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_804_inst
    process(a37_548, a47_612) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a37_548, a47_612, tmp_var);
      SGT_i16_u1_804_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_812_inst
    process(t71_800, t72_808) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t71_800, t72_808, tmp_var);
      SGT_i16_u1_812_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_820_inst
    process(a18_424, a28_488) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a18_424, a28_488, tmp_var);
      SGT_i16_u1_820_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_828_inst
    process(a38_552, a48_616) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a38_552, a48_616, tmp_var);
      SGT_i16_u1_828_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_836_inst
    process(t81_824, t82_832) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t81_824, t82_832, tmp_var);
      SGT_i16_u1_836_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_844_inst
    process(a19_428, a29_492) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a19_428, a29_492, tmp_var);
      SGT_i16_u1_844_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_852_inst
    process(a39_556, a49_620) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a39_556, a49_620, tmp_var);
      SGT_i16_u1_852_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_860_inst
    process(t91_848, t92_856) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t91_848, t92_856, tmp_var);
      SGT_i16_u1_860_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_868_inst
    process(a110_432, a210_496) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a110_432, a210_496, tmp_var);
      SGT_i16_u1_868_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_876_inst
    process(a310_560, a410_624) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a310_560, a410_624, tmp_var);
      SGT_i16_u1_876_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_884_inst
    process(t101_872, t102_880) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t101_872, t102_880, tmp_var);
      SGT_i16_u1_884_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_892_inst
    process(a111_436, a211_500) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a111_436, a211_500, tmp_var);
      SGT_i16_u1_892_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_900_inst
    process(a311_564, a411_628) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a311_564, a411_628, tmp_var);
      SGT_i16_u1_900_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_908_inst
    process(t111_896, t112_904) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t111_896, t112_904, tmp_var);
      SGT_i16_u1_908_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_916_inst
    process(a112_440, a212_504) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a112_440, a212_504, tmp_var);
      SGT_i16_u1_916_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_924_inst
    process(a312_568, a412_632) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a312_568, a412_632, tmp_var);
      SGT_i16_u1_924_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_932_inst
    process(t121_920, t122_928) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t121_920, t122_928, tmp_var);
      SGT_i16_u1_932_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_940_inst
    process(a113_444, a213_508) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a113_444, a213_508, tmp_var);
      SGT_i16_u1_940_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_948_inst
    process(a313_572, a413_636) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a313_572, a413_636, tmp_var);
      SGT_i16_u1_948_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_956_inst
    process(t131_944, t132_952) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t131_944, t132_952, tmp_var);
      SGT_i16_u1_956_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_964_inst
    process(a114_448, a214_512) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a114_448, a214_512, tmp_var);
      SGT_i16_u1_964_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_972_inst
    process(a314_576, a414_640) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a314_576, a414_640, tmp_var);
      SGT_i16_u1_972_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_980_inst
    process(t141_968, t142_976) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(t141_968, t142_976, tmp_var);
      SGT_i16_u1_980_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_988_inst
    process(a115_452, a215_516) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a115_452, a215_516, tmp_var);
      SGT_i16_u1_988_wire <= tmp_var; --
    end process;
    -- binary operator SGT_i16_u1_996_inst
    process(a315_580, a415_644) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntSgt_proc(a315_580, a415_644, tmp_var);
      SGT_i16_u1_996_wire <= tmp_var; --
    end process;
    -- shared split operator group (63) : array_obj_ref_102_index_offset 
    ApIntAdd_group_63: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_addr2_101_scaled;
      array_obj_ref_102_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_102_index_offset_req_0;
      array_obj_ref_102_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_102_index_offset_req_1;
      array_obj_ref_102_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_63_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_63_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_63",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 63
    -- shared split operator group (64) : array_obj_ref_1037_index_offset 
    ApIntAdd_group_64: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_addr_1036_scaled;
      array_obj_ref_1037_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1037_index_offset_req_0;
      array_obj_ref_1037_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1037_index_offset_req_1;
      array_obj_ref_1037_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_64_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_64_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_64",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 64
    -- shared split operator group (65) : array_obj_ref_1063_index_offset 
    ApIntAdd_group_65: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ADD_u32_u32_1062_scaled;
      array_obj_ref_1063_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1063_index_offset_req_0;
      array_obj_ref_1063_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1063_index_offset_req_1;
      array_obj_ref_1063_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_65_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_65_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_65",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 65
    -- shared split operator group (66) : array_obj_ref_1089_index_offset 
    ApIntAdd_group_66: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ADD_u32_u32_1088_scaled;
      array_obj_ref_1089_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1089_index_offset_req_0;
      array_obj_ref_1089_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1089_index_offset_req_1;
      array_obj_ref_1089_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_66_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_66_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_66",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 66
    -- shared split operator group (67) : array_obj_ref_109_index_offset 
    ApIntAdd_group_67: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_addr3_108_scaled;
      array_obj_ref_109_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_109_index_offset_req_0;
      array_obj_ref_109_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_109_index_offset_req_1;
      array_obj_ref_109_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_67_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_67_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_67",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 67
    -- shared split operator group (68) : array_obj_ref_1115_index_offset 
    ApIntAdd_group_68: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ADD_u32_u32_1114_scaled;
      array_obj_ref_1115_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1115_index_offset_req_0;
      array_obj_ref_1115_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1115_index_offset_req_1;
      array_obj_ref_1115_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_68_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_68_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_68",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 68
    -- shared split operator group (69) : array_obj_ref_116_index_offset 
    ApIntAdd_group_69: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_addr4_115_scaled;
      array_obj_ref_116_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_116_index_offset_req_0;
      array_obj_ref_116_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_116_index_offset_req_1;
      array_obj_ref_116_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_69_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_69_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_69",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 69
    -- shared split operator group (70) : array_obj_ref_95_index_offset 
    ApIntAdd_group_70: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_addr1_94_scaled;
      array_obj_ref_95_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_95_index_offset_req_0;
      array_obj_ref_95_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_95_index_offset_req_1;
      array_obj_ref_95_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_70_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_70_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_70",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 70
    -- shared load operator group (0) : ptr_deref_121_load_0 ptr_deref_125_load_0 ptr_deref_129_load_0 ptr_deref_133_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(55 downto 0);
      signal data_out: std_logic_vector(1023 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 3 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 3 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 3 downto 0);
      signal guard_vector : std_logic_vector( 3 downto 0);
      constant inBUFs : IntegerArray(3 downto 0) := (3 => 2, 2 => 2, 1 => 2, 0 => 2);
      constant outBUFs : IntegerArray(3 downto 0) := (3 => 2, 2 => 2, 1 => 2, 0 => 2);
      constant guardFlags : BooleanArray(3 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false);
      constant guardBuffering: IntegerArray(3 downto 0)  := (0 => 6, 1 => 6, 2 => 6, 3 => 6);
      -- 
    begin -- 
      reqL_unguarded(3) <= ptr_deref_121_load_0_req_0;
      reqL_unguarded(2) <= ptr_deref_125_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_129_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_133_load_0_req_0;
      ptr_deref_121_load_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_125_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_129_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_133_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(3) <= ptr_deref_121_load_0_req_1;
      reqR_unguarded(2) <= ptr_deref_125_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_129_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_133_load_0_req_1;
      ptr_deref_121_load_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_125_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_129_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_133_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 4, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_121_word_address_0 & ptr_deref_125_word_address_0 & ptr_deref_129_word_address_0 & ptr_deref_133_word_address_0;
      ptr_deref_121_data_0 <= data_out(1023 downto 768);
      ptr_deref_125_data_0 <= data_out(767 downto 512);
      ptr_deref_129_data_0 <= data_out(511 downto 256);
      ptr_deref_133_data_0 <= data_out(255 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 4,
        tag_length => 3,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 256,
        num_reqs => 4,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(255 downto 0),
          mtag => memory_space_1_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_1044_store_0 ptr_deref_1070_store_0 ptr_deref_1096_store_0 ptr_deref_1122_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(55 downto 0);
      signal data_in: std_logic_vector(255 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 3 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 3 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 3 downto 0);
      signal guard_vector : std_logic_vector( 3 downto 0);
      constant inBUFs : IntegerArray(3 downto 0) := (3 => 2, 2 => 2, 1 => 2, 0 => 2);
      constant outBUFs : IntegerArray(3 downto 0) := (3 => 15, 2 => 15, 1 => 15, 0 => 15);
      constant guardFlags : BooleanArray(3 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false);
      constant guardBuffering: IntegerArray(3 downto 0)  := (0 => 6, 1 => 6, 2 => 6, 3 => 6);
      -- 
    begin -- 
      reqL_unguarded(3) <= ptr_deref_1044_store_0_req_0;
      reqL_unguarded(2) <= ptr_deref_1070_store_0_req_0;
      reqL_unguarded(1) <= ptr_deref_1096_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1122_store_0_req_0;
      ptr_deref_1044_store_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_1070_store_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_1096_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1122_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(3) <= ptr_deref_1044_store_0_req_1;
      reqR_unguarded(2) <= ptr_deref_1070_store_0_req_1;
      reqR_unguarded(1) <= ptr_deref_1096_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1122_store_0_req_1;
      ptr_deref_1044_store_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_1070_store_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_1096_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1122_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      StoreGroup0_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_2: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_3: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 4, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1044_word_address_0 & ptr_deref_1070_word_address_0 & ptr_deref_1096_word_address_0 & ptr_deref_1122_word_address_0;
      data_in <= ptr_deref_1044_data_0 & ptr_deref_1070_data_0 & ptr_deref_1096_data_0 & ptr_deref_1122_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 4,
        tag_length => 3,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(13 downto 0),
          mdata => memory_space_0_sr_data(63 downto 0),
          mtag => memory_space_0_sr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 4,
          detailed_buffering_per_output => outBUFs,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end maxPool4_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity sendB is -- 
  generic (tag_length : integer); 
  port ( -- 
    size : in  std_logic_vector(31 downto 0);
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
    maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity sendB;
architecture sendB_arch of sendB is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 32)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal size_buffer :  std_logic_vector(31 downto 0);
  signal size_update_enable: Boolean;
  -- output port buffer signals
  signal sendB_CP_2164_start: Boolean;
  signal sendB_CP_2164_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal addr_of_1206_final_reg_ack_0 : boolean;
  signal type_cast_1176_inst_req_1 : boolean;
  signal if_stmt_1149_branch_ack_0 : boolean;
  signal array_obj_ref_1205_index_offset_req_0 : boolean;
  signal type_cast_1176_inst_req_0 : boolean;
  signal type_cast_1176_inst_ack_0 : boolean;
  signal addr_of_1206_final_reg_ack_1 : boolean;
  signal type_cast_1176_inst_ack_1 : boolean;
  signal if_stmt_1149_branch_ack_1 : boolean;
  signal array_obj_ref_1205_index_offset_ack_1 : boolean;
  signal array_obj_ref_1205_index_offset_req_1 : boolean;
  signal addr_of_1206_final_reg_req_1 : boolean;
  signal array_obj_ref_1205_index_offset_ack_0 : boolean;
  signal ptr_deref_1210_load_0_ack_1 : boolean;
  signal ptr_deref_1210_load_0_req_1 : boolean;
  signal ptr_deref_1210_load_0_req_0 : boolean;
  signal if_stmt_1149_branch_req_0 : boolean;
  signal type_cast_1256_inst_req_1 : boolean;
  signal type_cast_1256_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1258_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1258_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1258_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1258_inst_ack_0 : boolean;
  signal ptr_deref_1210_load_0_ack_0 : boolean;
  signal addr_of_1206_final_reg_req_0 : boolean;
  signal type_cast_1256_inst_ack_0 : boolean;
  signal type_cast_1256_inst_ack_1 : boolean;
  signal type_cast_1263_inst_req_0 : boolean;
  signal type_cast_1263_inst_ack_0 : boolean;
  signal type_cast_1263_inst_req_1 : boolean;
  signal type_cast_1263_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1265_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1265_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1265_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1265_inst_ack_1 : boolean;
  signal type_cast_1270_inst_req_0 : boolean;
  signal type_cast_1270_inst_ack_0 : boolean;
  signal type_cast_1270_inst_req_1 : boolean;
  signal type_cast_1270_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1272_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1272_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1272_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1272_inst_ack_1 : boolean;
  signal type_cast_1277_inst_req_0 : boolean;
  signal type_cast_1277_inst_ack_0 : boolean;
  signal type_cast_1277_inst_req_1 : boolean;
  signal type_cast_1277_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1279_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1279_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1279_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1279_inst_ack_1 : boolean;
  signal type_cast_1284_inst_req_0 : boolean;
  signal type_cast_1284_inst_ack_0 : boolean;
  signal type_cast_1284_inst_req_1 : boolean;
  signal type_cast_1284_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1286_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1286_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1286_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1286_inst_ack_1 : boolean;
  signal type_cast_1291_inst_req_0 : boolean;
  signal type_cast_1291_inst_ack_0 : boolean;
  signal type_cast_1291_inst_req_1 : boolean;
  signal type_cast_1291_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1293_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1293_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1293_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1293_inst_ack_1 : boolean;
  signal type_cast_1298_inst_req_0 : boolean;
  signal type_cast_1298_inst_ack_0 : boolean;
  signal type_cast_1298_inst_req_1 : boolean;
  signal type_cast_1298_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1300_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1300_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1300_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1300_inst_ack_1 : boolean;
  signal type_cast_1305_inst_req_0 : boolean;
  signal type_cast_1305_inst_ack_0 : boolean;
  signal type_cast_1305_inst_req_1 : boolean;
  signal type_cast_1305_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1307_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1307_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1307_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1307_inst_ack_1 : boolean;
  signal if_stmt_1321_branch_req_0 : boolean;
  signal if_stmt_1321_branch_ack_1 : boolean;
  signal if_stmt_1321_branch_ack_0 : boolean;
  signal phi_stmt_1193_req_0 : boolean;
  signal type_cast_1199_inst_req_0 : boolean;
  signal type_cast_1199_inst_ack_0 : boolean;
  signal type_cast_1199_inst_req_1 : boolean;
  signal type_cast_1199_inst_ack_1 : boolean;
  signal phi_stmt_1193_req_1 : boolean;
  signal phi_stmt_1193_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "sendB_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 32) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(31 downto 0) <= size;
  size_buffer <= in_buffer_data_out(31 downto 0);
  in_buffer_data_in(tag_length + 31 downto 32) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 31 downto 32);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  sendB_CP_2164_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "sendB_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendB_CP_2164_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= sendB_CP_2164_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendB_CP_2164_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  sendB_CP_2164: Block -- control-path 
    signal sendB_CP_2164_elements: BooleanArray(59 downto 0);
    -- 
  begin -- 
    sendB_CP_2164_elements(0) <= sendB_CP_2164_start;
    sendB_CP_2164_symbol <= sendB_CP_2164_elements(59);
    -- CP-element group 0:  branch  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (15) 
      -- CP-element group 0: 	 branch_block_stmt_1142/$entry
      -- CP-element group 0: 	 branch_block_stmt_1142/if_stmt_1149_else_link/$entry
      -- CP-element group 0: 	 branch_block_stmt_1142/R_cmp76_1150_place
      -- CP-element group 0: 	 branch_block_stmt_1142/assign_stmt_1148/$exit
      -- CP-element group 0: 	 branch_block_stmt_1142/assign_stmt_1148__exit__
      -- CP-element group 0: 	 branch_block_stmt_1142/if_stmt_1149__entry__
      -- CP-element group 0: 	 branch_block_stmt_1142/if_stmt_1149_dead_link/$entry
      -- CP-element group 0: 	 branch_block_stmt_1142/if_stmt_1149_if_link/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1142/assign_stmt_1148__entry__
      -- CP-element group 0: 	 branch_block_stmt_1142/branch_block_stmt_1142__entry__
      -- CP-element group 0: 	 branch_block_stmt_1142/if_stmt_1149_eval_test/$entry
      -- CP-element group 0: 	 branch_block_stmt_1142/if_stmt_1149_eval_test/$exit
      -- CP-element group 0: 	 branch_block_stmt_1142/if_stmt_1149_eval_test/branch_req
      -- CP-element group 0: 	 branch_block_stmt_1142/assign_stmt_1148/$entry
      -- 
    branch_req_2202_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2202_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2164_elements(0), ack => if_stmt_1149_branch_req_0); -- 
    -- CP-element group 1:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	4 
    -- CP-element group 1: 	3 
    -- CP-element group 1:  members (18) 
      -- CP-element group 1: 	 branch_block_stmt_1142/assign_stmt_1161_to_assign_stmt_1190/type_cast_1176_Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1142/assign_stmt_1161_to_assign_stmt_1190/type_cast_1176_Update/cr
      -- CP-element group 1: 	 branch_block_stmt_1142/entry_bbx_xnph
      -- CP-element group 1: 	 branch_block_stmt_1142/assign_stmt_1161_to_assign_stmt_1190/type_cast_1176_Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_1142/assign_stmt_1161_to_assign_stmt_1190/type_cast_1176_sample_start_
      -- CP-element group 1: 	 branch_block_stmt_1142/assign_stmt_1161_to_assign_stmt_1190/$entry
      -- CP-element group 1: 	 branch_block_stmt_1142/assign_stmt_1161_to_assign_stmt_1190/type_cast_1176_update_start_
      -- CP-element group 1: 	 branch_block_stmt_1142/assign_stmt_1161_to_assign_stmt_1190/type_cast_1176_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1142/if_stmt_1149_if_link/if_choice_transition
      -- CP-element group 1: 	 branch_block_stmt_1142/merge_stmt_1155__exit__
      -- CP-element group 1: 	 branch_block_stmt_1142/if_stmt_1149_if_link/$exit
      -- CP-element group 1: 	 branch_block_stmt_1142/assign_stmt_1161_to_assign_stmt_1190__entry__
      -- CP-element group 1: 	 branch_block_stmt_1142/entry_bbx_xnph_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_1142/entry_bbx_xnph_PhiReq/$exit
      -- CP-element group 1: 	 branch_block_stmt_1142/merge_stmt_1155_PhiReqMerge
      -- CP-element group 1: 	 branch_block_stmt_1142/merge_stmt_1155_PhiAck/$entry
      -- CP-element group 1: 	 branch_block_stmt_1142/merge_stmt_1155_PhiAck/$exit
      -- CP-element group 1: 	 branch_block_stmt_1142/merge_stmt_1155_PhiAck/dummy
      -- 
    if_choice_transition_2207_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1149_branch_ack_1, ack => sendB_CP_2164_elements(1)); -- 
    cr_2229_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2229_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2164_elements(1), ack => type_cast_1176_inst_req_1); -- 
    rr_2224_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2224_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2164_elements(1), ack => type_cast_1176_inst_req_0); -- 
    -- CP-element group 2:  transition  place  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	59 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 branch_block_stmt_1142/if_stmt_1149_else_link/$exit
      -- CP-element group 2: 	 branch_block_stmt_1142/if_stmt_1149_else_link/else_choice_transition
      -- CP-element group 2: 	 branch_block_stmt_1142/entry_forx_xend
      -- CP-element group 2: 	 branch_block_stmt_1142/entry_forx_xend_PhiReq/$entry
      -- CP-element group 2: 	 branch_block_stmt_1142/entry_forx_xend_PhiReq/$exit
      -- 
    else_choice_transition_2211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1149_branch_ack_0, ack => sendB_CP_2164_elements(2)); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	1 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_1142/assign_stmt_1161_to_assign_stmt_1190/type_cast_1176_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_1142/assign_stmt_1161_to_assign_stmt_1190/type_cast_1176_Sample/ra
      -- CP-element group 3: 	 branch_block_stmt_1142/assign_stmt_1161_to_assign_stmt_1190/type_cast_1176_sample_completed_
      -- 
    ra_2225_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1176_inst_ack_0, ack => sendB_CP_2164_elements(3)); -- 
    -- CP-element group 4:  transition  place  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	1 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	53 
    -- CP-element group 4:  members (9) 
      -- CP-element group 4: 	 branch_block_stmt_1142/assign_stmt_1161_to_assign_stmt_1190/type_cast_1176_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_1142/assign_stmt_1161_to_assign_stmt_1190__exit__
      -- CP-element group 4: 	 branch_block_stmt_1142/assign_stmt_1161_to_assign_stmt_1190/type_cast_1176_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_1142/assign_stmt_1161_to_assign_stmt_1190/type_cast_1176_Update/ca
      -- CP-element group 4: 	 branch_block_stmt_1142/assign_stmt_1161_to_assign_stmt_1190/$exit
      -- CP-element group 4: 	 branch_block_stmt_1142/bbx_xnph_forx_xbody
      -- CP-element group 4: 	 branch_block_stmt_1142/bbx_xnph_forx_xbody_PhiReq/$entry
      -- CP-element group 4: 	 branch_block_stmt_1142/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1193/$entry
      -- CP-element group 4: 	 branch_block_stmt_1142/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1193/phi_stmt_1193_sources/$entry
      -- 
    ca_2230_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1176_inst_ack_1, ack => sendB_CP_2164_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	58 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	50 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/array_obj_ref_1205_final_index_sum_regn_sample_complete
      -- CP-element group 5: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/array_obj_ref_1205_final_index_sum_regn_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/array_obj_ref_1205_final_index_sum_regn_Sample/ack
      -- 
    ack_2259_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1205_index_offset_ack_0, ack => sendB_CP_2164_elements(5)); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	58 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (11) 
      -- CP-element group 6: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/array_obj_ref_1205_base_plus_offset/sum_rename_req
      -- CP-element group 6: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/array_obj_ref_1205_base_plus_offset/$exit
      -- CP-element group 6: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/array_obj_ref_1205_base_plus_offset/$entry
      -- CP-element group 6: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/addr_of_1206_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/array_obj_ref_1205_final_index_sum_regn_Update/ack
      -- CP-element group 6: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/array_obj_ref_1205_base_plus_offset/sum_rename_ack
      -- CP-element group 6: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/array_obj_ref_1205_final_index_sum_regn_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/array_obj_ref_1205_offset_calculated
      -- CP-element group 6: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/array_obj_ref_1205_root_address_calculated
      -- CP-element group 6: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/addr_of_1206_request/$entry
      -- CP-element group 6: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/addr_of_1206_request/req
      -- 
    ack_2264_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1205_index_offset_ack_1, ack => sendB_CP_2164_elements(6)); -- 
    req_2273_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2273_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2164_elements(6), ack => addr_of_1206_final_reg_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/addr_of_1206_request/ack
      -- CP-element group 7: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/addr_of_1206_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/addr_of_1206_request/$exit
      -- 
    ack_2274_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1206_final_reg_ack_0, ack => sendB_CP_2164_elements(7)); -- 
    -- CP-element group 8:  join  fork  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	58 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (24) 
      -- CP-element group 8: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/ptr_deref_1210_base_addr_resize/$exit
      -- CP-element group 8: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/ptr_deref_1210_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/ptr_deref_1210_word_address_calculated
      -- CP-element group 8: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/ptr_deref_1210_base_plus_offset/$exit
      -- CP-element group 8: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/addr_of_1206_complete/ack
      -- CP-element group 8: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/ptr_deref_1210_base_plus_offset/sum_rename_ack
      -- CP-element group 8: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/ptr_deref_1210_base_address_calculated
      -- CP-element group 8: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/addr_of_1206_complete/$exit
      -- CP-element group 8: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/ptr_deref_1210_base_addr_resize/$entry
      -- CP-element group 8: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/ptr_deref_1210_word_addrgen/root_register_ack
      -- CP-element group 8: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/ptr_deref_1210_word_addrgen/root_register_req
      -- CP-element group 8: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/addr_of_1206_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/ptr_deref_1210_base_plus_offset/sum_rename_req
      -- CP-element group 8: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/ptr_deref_1210_root_address_calculated
      -- CP-element group 8: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/ptr_deref_1210_word_addrgen/$entry
      -- CP-element group 8: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/ptr_deref_1210_base_address_resized
      -- CP-element group 8: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/ptr_deref_1210_base_addr_resize/base_resize_ack
      -- CP-element group 8: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/ptr_deref_1210_word_addrgen/$exit
      -- CP-element group 8: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/ptr_deref_1210_base_addr_resize/base_resize_req
      -- CP-element group 8: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/ptr_deref_1210_Sample/word_access_start/word_0/$entry
      -- CP-element group 8: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/ptr_deref_1210_Sample/word_access_start/word_0/rr
      -- CP-element group 8: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/ptr_deref_1210_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/ptr_deref_1210_Sample/word_access_start/$entry
      -- CP-element group 8: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/ptr_deref_1210_base_plus_offset/$entry
      -- 
    ack_2279_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1206_final_reg_ack_1, ack => sendB_CP_2164_elements(8)); -- 
    rr_2312_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2312_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2164_elements(8), ack => ptr_deref_1210_load_0_req_0); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (5) 
      -- CP-element group 9: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/ptr_deref_1210_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/ptr_deref_1210_Sample/word_access_start/$exit
      -- CP-element group 9: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/ptr_deref_1210_Sample/word_access_start/word_0/$exit
      -- CP-element group 9: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/ptr_deref_1210_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/ptr_deref_1210_Sample/word_access_start/word_0/ra
      -- 
    ra_2313_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1210_load_0_ack_0, ack => sendB_CP_2164_elements(9)); -- 
    -- CP-element group 10:  fork  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	58 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10: 	15 
    -- CP-element group 10: 	20 
    -- CP-element group 10: 	25 
    -- CP-element group 10: 	30 
    -- CP-element group 10: 	35 
    -- CP-element group 10: 	40 
    -- CP-element group 10: 	45 
    -- CP-element group 10:  members (33) 
      -- CP-element group 10: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/ptr_deref_1210_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/ptr_deref_1210_Update/word_access_complete/$exit
      -- CP-element group 10: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/ptr_deref_1210_Update/word_access_complete/word_0/ca
      -- CP-element group 10: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/ptr_deref_1210_Update/ptr_deref_1210_Merge/merge_req
      -- CP-element group 10: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1256_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/ptr_deref_1210_Update/ptr_deref_1210_Merge/$entry
      -- CP-element group 10: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/ptr_deref_1210_Update/ptr_deref_1210_Merge/$exit
      -- CP-element group 10: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1256_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1256_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/ptr_deref_1210_Update/word_access_complete/word_0/$exit
      -- CP-element group 10: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/ptr_deref_1210_Update/ptr_deref_1210_Merge/merge_ack
      -- CP-element group 10: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/ptr_deref_1210_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1263_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1263_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1263_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1270_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1270_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1270_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1277_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1277_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1277_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1284_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1284_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1284_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1291_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1291_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1291_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1298_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1298_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1298_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1305_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1305_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1305_Sample/rr
      -- 
    ca_2324_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1210_load_0_ack_1, ack => sendB_CP_2164_elements(10)); -- 
    rr_2337_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2337_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2164_elements(10), ack => type_cast_1256_inst_req_0); -- 
    rr_2365_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2365_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2164_elements(10), ack => type_cast_1263_inst_req_0); -- 
    rr_2393_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2393_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2164_elements(10), ack => type_cast_1270_inst_req_0); -- 
    rr_2421_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2421_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2164_elements(10), ack => type_cast_1277_inst_req_0); -- 
    rr_2449_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2449_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2164_elements(10), ack => type_cast_1284_inst_req_0); -- 
    rr_2477_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2477_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2164_elements(10), ack => type_cast_1291_inst_req_0); -- 
    rr_2505_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2505_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2164_elements(10), ack => type_cast_1298_inst_req_0); -- 
    rr_2533_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2533_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2164_elements(10), ack => type_cast_1305_inst_req_0); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1256_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1256_Sample/ra
      -- CP-element group 11: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1256_sample_completed_
      -- 
    ra_2338_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1256_inst_ack_0, ack => sendB_CP_2164_elements(11)); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	58 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1256_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1258_sample_start_
      -- CP-element group 12: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1258_Sample/req
      -- CP-element group 12: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1256_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1256_Update/ca
      -- CP-element group 12: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1258_Sample/$entry
      -- 
    ca_2343_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1256_inst_ack_1, ack => sendB_CP_2164_elements(12)); -- 
    req_2351_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2351_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2164_elements(12), ack => WPIPE_maxpool_output_pipe_1258_inst_req_0); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1258_Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1258_Update/req
      -- CP-element group 13: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1258_Sample/ack
      -- CP-element group 13: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1258_update_start_
      -- CP-element group 13: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1258_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1258_sample_completed_
      -- 
    ack_2352_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1258_inst_ack_0, ack => sendB_CP_2164_elements(13)); -- 
    req_2356_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2356_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2164_elements(13), ack => WPIPE_maxpool_output_pipe_1258_inst_req_1); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	17 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1258_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1258_Update/ack
      -- CP-element group 14: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1258_update_completed_
      -- 
    ack_2357_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1258_inst_ack_1, ack => sendB_CP_2164_elements(14)); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	10 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1263_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1263_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1263_Sample/ra
      -- 
    ra_2366_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1263_inst_ack_0, ack => sendB_CP_2164_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	58 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1263_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1263_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1263_Update/ca
      -- 
    ca_2371_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1263_inst_ack_1, ack => sendB_CP_2164_elements(16)); -- 
    -- CP-element group 17:  join  transition  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	14 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1265_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1265_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1265_Sample/req
      -- 
    req_2379_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2379_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2164_elements(17), ack => WPIPE_maxpool_output_pipe_1265_inst_req_0); -- 
    sendB_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_2164_elements(14) & sendB_CP_2164_elements(16);
      gj_sendB_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2164_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1265_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1265_update_start_
      -- CP-element group 18: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1265_Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1265_Sample/ack
      -- CP-element group 18: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1265_Update/$entry
      -- CP-element group 18: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1265_Update/req
      -- 
    ack_2380_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1265_inst_ack_0, ack => sendB_CP_2164_elements(18)); -- 
    req_2384_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2384_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2164_elements(18), ack => WPIPE_maxpool_output_pipe_1265_inst_req_1); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	22 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1265_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1265_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1265_Update/ack
      -- 
    ack_2385_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1265_inst_ack_1, ack => sendB_CP_2164_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	10 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1270_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1270_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1270_Sample/ra
      -- 
    ra_2394_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1270_inst_ack_0, ack => sendB_CP_2164_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	58 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1270_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1270_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1270_Update/ca
      -- 
    ca_2399_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1270_inst_ack_1, ack => sendB_CP_2164_elements(21)); -- 
    -- CP-element group 22:  join  transition  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	19 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1272_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1272_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1272_Sample/req
      -- 
    req_2407_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2407_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2164_elements(22), ack => WPIPE_maxpool_output_pipe_1272_inst_req_0); -- 
    sendB_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_2164_elements(19) & sendB_CP_2164_elements(21);
      gj_sendB_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2164_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  transition  input  output  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23:  members (6) 
      -- CP-element group 23: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1272_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1272_update_start_
      -- CP-element group 23: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1272_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1272_Sample/ack
      -- CP-element group 23: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1272_Update/$entry
      -- CP-element group 23: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1272_Update/req
      -- 
    ack_2408_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1272_inst_ack_0, ack => sendB_CP_2164_elements(23)); -- 
    req_2412_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2412_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2164_elements(23), ack => WPIPE_maxpool_output_pipe_1272_inst_req_1); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	27 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1272_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1272_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1272_Update/ack
      -- 
    ack_2413_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1272_inst_ack_1, ack => sendB_CP_2164_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	10 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1277_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1277_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1277_Sample/ra
      -- 
    ra_2422_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1277_inst_ack_0, ack => sendB_CP_2164_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	58 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1277_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1277_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1277_Update/ca
      -- 
    ca_2427_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1277_inst_ack_1, ack => sendB_CP_2164_elements(26)); -- 
    -- CP-element group 27:  join  transition  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	24 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1279_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1279_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1279_Sample/req
      -- 
    req_2435_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2435_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2164_elements(27), ack => WPIPE_maxpool_output_pipe_1279_inst_req_0); -- 
    sendB_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_2164_elements(24) & sendB_CP_2164_elements(26);
      gj_sendB_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2164_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  transition  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (6) 
      -- CP-element group 28: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1279_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1279_update_start_
      -- CP-element group 28: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1279_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1279_Sample/ack
      -- CP-element group 28: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1279_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1279_Update/req
      -- 
    ack_2436_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1279_inst_ack_0, ack => sendB_CP_2164_elements(28)); -- 
    req_2440_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2440_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2164_elements(28), ack => WPIPE_maxpool_output_pipe_1279_inst_req_1); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	32 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1279_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1279_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1279_Update/ack
      -- 
    ack_2441_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1279_inst_ack_1, ack => sendB_CP_2164_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	10 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1284_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1284_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1284_Sample/ra
      -- 
    ra_2450_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1284_inst_ack_0, ack => sendB_CP_2164_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	58 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1284_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1284_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1284_Update/ca
      -- 
    ca_2455_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1284_inst_ack_1, ack => sendB_CP_2164_elements(31)); -- 
    -- CP-element group 32:  join  transition  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	29 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1286_sample_start_
      -- CP-element group 32: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1286_Sample/$entry
      -- CP-element group 32: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1286_Sample/req
      -- 
    req_2463_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2463_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2164_elements(32), ack => WPIPE_maxpool_output_pipe_1286_inst_req_0); -- 
    sendB_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_2164_elements(29) & sendB_CP_2164_elements(31);
      gj_sendB_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2164_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (6) 
      -- CP-element group 33: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1286_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1286_update_start_
      -- CP-element group 33: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1286_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1286_Sample/ack
      -- CP-element group 33: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1286_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1286_Update/req
      -- 
    ack_2464_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1286_inst_ack_0, ack => sendB_CP_2164_elements(33)); -- 
    req_2468_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2468_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2164_elements(33), ack => WPIPE_maxpool_output_pipe_1286_inst_req_1); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	37 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1286_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1286_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1286_Update/ack
      -- 
    ack_2469_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1286_inst_ack_1, ack => sendB_CP_2164_elements(34)); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	10 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1291_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1291_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1291_Sample/ra
      -- 
    ra_2478_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1291_inst_ack_0, ack => sendB_CP_2164_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	58 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	37 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1291_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1291_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1291_Update/ca
      -- 
    ca_2483_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1291_inst_ack_1, ack => sendB_CP_2164_elements(36)); -- 
    -- CP-element group 37:  join  transition  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: 	36 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1293_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1293_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1293_Sample/req
      -- 
    req_2491_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2491_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2164_elements(37), ack => WPIPE_maxpool_output_pipe_1293_inst_req_0); -- 
    sendB_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_2164_elements(34) & sendB_CP_2164_elements(36);
      gj_sendB_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2164_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (6) 
      -- CP-element group 38: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1293_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1293_update_start_
      -- CP-element group 38: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1293_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1293_Sample/ack
      -- CP-element group 38: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1293_Update/$entry
      -- CP-element group 38: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1293_Update/req
      -- 
    ack_2492_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1293_inst_ack_0, ack => sendB_CP_2164_elements(38)); -- 
    req_2496_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2496_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2164_elements(38), ack => WPIPE_maxpool_output_pipe_1293_inst_req_1); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	42 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1293_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1293_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1293_Update/ack
      -- 
    ack_2497_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1293_inst_ack_1, ack => sendB_CP_2164_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	10 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1298_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1298_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1298_Sample/ra
      -- 
    ra_2506_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1298_inst_ack_0, ack => sendB_CP_2164_elements(40)); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	58 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1298_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1298_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1298_Update/ca
      -- 
    ca_2511_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1298_inst_ack_1, ack => sendB_CP_2164_elements(41)); -- 
    -- CP-element group 42:  join  transition  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	39 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1300_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1300_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1300_Sample/req
      -- 
    req_2519_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2519_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2164_elements(42), ack => WPIPE_maxpool_output_pipe_1300_inst_req_0); -- 
    sendB_cp_element_group_42: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_42"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_2164_elements(39) & sendB_CP_2164_elements(41);
      gj_sendB_cp_element_group_42 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2164_elements(42), clk => clk, reset => reset); --
    end block;
    -- CP-element group 43:  transition  input  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (6) 
      -- CP-element group 43: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1300_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1300_update_start_
      -- CP-element group 43: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1300_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1300_Sample/ack
      -- CP-element group 43: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1300_Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1300_Update/req
      -- 
    ack_2520_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1300_inst_ack_0, ack => sendB_CP_2164_elements(43)); -- 
    req_2524_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2524_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2164_elements(43), ack => WPIPE_maxpool_output_pipe_1300_inst_req_1); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	47 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1300_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1300_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1300_Update/ack
      -- 
    ack_2525_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1300_inst_ack_1, ack => sendB_CP_2164_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	10 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1305_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1305_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1305_Sample/ra
      -- 
    ra_2534_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1305_inst_ack_0, ack => sendB_CP_2164_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	58 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1305_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1305_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1305_Update/ca
      -- 
    ca_2539_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1305_inst_ack_1, ack => sendB_CP_2164_elements(46)); -- 
    -- CP-element group 47:  join  transition  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	44 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1307_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1307_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1307_Sample/req
      -- 
    req_2547_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2547_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2164_elements(47), ack => WPIPE_maxpool_output_pipe_1307_inst_req_0); -- 
    sendB_cp_element_group_47: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_47"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_2164_elements(44) & sendB_CP_2164_elements(46);
      gj_sendB_cp_element_group_47 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2164_elements(47), clk => clk, reset => reset); --
    end block;
    -- CP-element group 48:  transition  input  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (6) 
      -- CP-element group 48: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1307_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1307_update_start_
      -- CP-element group 48: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1307_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1307_Sample/ack
      -- CP-element group 48: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1307_Update/$entry
      -- CP-element group 48: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1307_Update/req
      -- 
    ack_2548_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1307_inst_ack_0, ack => sendB_CP_2164_elements(48)); -- 
    req_2552_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2552_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2164_elements(48), ack => WPIPE_maxpool_output_pipe_1307_inst_req_1); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1307_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1307_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/WPIPE_maxpool_output_pipe_1307_Update/ack
      -- 
    ack_2553_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1307_inst_ack_1, ack => sendB_CP_2164_elements(49)); -- 
    -- CP-element group 50:  branch  join  transition  place  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	5 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (10) 
      -- CP-element group 50: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/$exit
      -- CP-element group 50: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320__exit__
      -- CP-element group 50: 	 branch_block_stmt_1142/if_stmt_1321__entry__
      -- CP-element group 50: 	 branch_block_stmt_1142/if_stmt_1321_dead_link/$entry
      -- CP-element group 50: 	 branch_block_stmt_1142/if_stmt_1321_eval_test/$entry
      -- CP-element group 50: 	 branch_block_stmt_1142/if_stmt_1321_eval_test/$exit
      -- CP-element group 50: 	 branch_block_stmt_1142/if_stmt_1321_eval_test/branch_req
      -- CP-element group 50: 	 branch_block_stmt_1142/R_exitcond1_1322_place
      -- CP-element group 50: 	 branch_block_stmt_1142/if_stmt_1321_if_link/$entry
      -- CP-element group 50: 	 branch_block_stmt_1142/if_stmt_1321_else_link/$entry
      -- 
    branch_req_2561_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2561_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2164_elements(50), ack => if_stmt_1321_branch_req_0); -- 
    sendB_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_2164_elements(5) & sendB_CP_2164_elements(49);
      gj_sendB_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2164_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  merge  transition  place  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	59 
    -- CP-element group 51:  members (13) 
      -- CP-element group 51: 	 branch_block_stmt_1142/merge_stmt_1327__exit__
      -- CP-element group 51: 	 branch_block_stmt_1142/forx_xendx_xloopexit_forx_xend
      -- CP-element group 51: 	 branch_block_stmt_1142/if_stmt_1321_if_link/$exit
      -- CP-element group 51: 	 branch_block_stmt_1142/if_stmt_1321_if_link/if_choice_transition
      -- CP-element group 51: 	 branch_block_stmt_1142/forx_xbody_forx_xendx_xloopexit
      -- CP-element group 51: 	 branch_block_stmt_1142/forx_xbody_forx_xendx_xloopexit_PhiReq/$entry
      -- CP-element group 51: 	 branch_block_stmt_1142/forx_xbody_forx_xendx_xloopexit_PhiReq/$exit
      -- CP-element group 51: 	 branch_block_stmt_1142/merge_stmt_1327_PhiReqMerge
      -- CP-element group 51: 	 branch_block_stmt_1142/merge_stmt_1327_PhiAck/$entry
      -- CP-element group 51: 	 branch_block_stmt_1142/merge_stmt_1327_PhiAck/$exit
      -- CP-element group 51: 	 branch_block_stmt_1142/merge_stmt_1327_PhiAck/dummy
      -- CP-element group 51: 	 branch_block_stmt_1142/forx_xendx_xloopexit_forx_xend_PhiReq/$entry
      -- CP-element group 51: 	 branch_block_stmt_1142/forx_xendx_xloopexit_forx_xend_PhiReq/$exit
      -- 
    if_choice_transition_2566_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1321_branch_ack_1, ack => sendB_CP_2164_elements(51)); -- 
    -- CP-element group 52:  fork  transition  place  input  output  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52: 	55 
    -- CP-element group 52:  members (12) 
      -- CP-element group 52: 	 branch_block_stmt_1142/if_stmt_1321_else_link/$exit
      -- CP-element group 52: 	 branch_block_stmt_1142/if_stmt_1321_else_link/else_choice_transition
      -- CP-element group 52: 	 branch_block_stmt_1142/forx_xbody_forx_xbody
      -- CP-element group 52: 	 branch_block_stmt_1142/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 52: 	 branch_block_stmt_1142/forx_xbody_forx_xbody_PhiReq/phi_stmt_1193/$entry
      -- CP-element group 52: 	 branch_block_stmt_1142/forx_xbody_forx_xbody_PhiReq/phi_stmt_1193/phi_stmt_1193_sources/$entry
      -- CP-element group 52: 	 branch_block_stmt_1142/forx_xbody_forx_xbody_PhiReq/phi_stmt_1193/phi_stmt_1193_sources/type_cast_1199/$entry
      -- CP-element group 52: 	 branch_block_stmt_1142/forx_xbody_forx_xbody_PhiReq/phi_stmt_1193/phi_stmt_1193_sources/type_cast_1199/SplitProtocol/$entry
      -- CP-element group 52: 	 branch_block_stmt_1142/forx_xbody_forx_xbody_PhiReq/phi_stmt_1193/phi_stmt_1193_sources/type_cast_1199/SplitProtocol/Sample/$entry
      -- CP-element group 52: 	 branch_block_stmt_1142/forx_xbody_forx_xbody_PhiReq/phi_stmt_1193/phi_stmt_1193_sources/type_cast_1199/SplitProtocol/Sample/rr
      -- CP-element group 52: 	 branch_block_stmt_1142/forx_xbody_forx_xbody_PhiReq/phi_stmt_1193/phi_stmt_1193_sources/type_cast_1199/SplitProtocol/Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_1142/forx_xbody_forx_xbody_PhiReq/phi_stmt_1193/phi_stmt_1193_sources/type_cast_1199/SplitProtocol/Update/cr
      -- 
    else_choice_transition_2570_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1321_branch_ack_0, ack => sendB_CP_2164_elements(52)); -- 
    rr_2614_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2614_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2164_elements(52), ack => type_cast_1199_inst_req_0); -- 
    cr_2619_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2619_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2164_elements(52), ack => type_cast_1199_inst_req_1); -- 
    -- CP-element group 53:  transition  output  delay-element  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	4 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	57 
    -- CP-element group 53:  members (5) 
      -- CP-element group 53: 	 branch_block_stmt_1142/bbx_xnph_forx_xbody_PhiReq/$exit
      -- CP-element group 53: 	 branch_block_stmt_1142/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1193/$exit
      -- CP-element group 53: 	 branch_block_stmt_1142/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1193/phi_stmt_1193_sources/$exit
      -- CP-element group 53: 	 branch_block_stmt_1142/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1193/phi_stmt_1193_sources/type_cast_1197_konst_delay_trans
      -- CP-element group 53: 	 branch_block_stmt_1142/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1193/phi_stmt_1193_req
      -- 
    phi_stmt_1193_req_2595_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1193_req_2595_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2164_elements(53), ack => phi_stmt_1193_req_0); -- 
    -- Element group sendB_CP_2164_elements(53) is a control-delay.
    cp_element_53_delay: control_delay_element  generic map(name => " 53_delay", delay_value => 1)  port map(req => sendB_CP_2164_elements(4), ack => sendB_CP_2164_elements(53), clk => clk, reset =>reset);
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	56 
    -- CP-element group 54:  members (2) 
      -- CP-element group 54: 	 branch_block_stmt_1142/forx_xbody_forx_xbody_PhiReq/phi_stmt_1193/phi_stmt_1193_sources/type_cast_1199/SplitProtocol/Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_1142/forx_xbody_forx_xbody_PhiReq/phi_stmt_1193/phi_stmt_1193_sources/type_cast_1199/SplitProtocol/Sample/ra
      -- 
    ra_2615_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1199_inst_ack_0, ack => sendB_CP_2164_elements(54)); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	52 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (2) 
      -- CP-element group 55: 	 branch_block_stmt_1142/forx_xbody_forx_xbody_PhiReq/phi_stmt_1193/phi_stmt_1193_sources/type_cast_1199/SplitProtocol/Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_1142/forx_xbody_forx_xbody_PhiReq/phi_stmt_1193/phi_stmt_1193_sources/type_cast_1199/SplitProtocol/Update/ca
      -- 
    ca_2620_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1199_inst_ack_1, ack => sendB_CP_2164_elements(55)); -- 
    -- CP-element group 56:  join  transition  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	54 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (6) 
      -- CP-element group 56: 	 branch_block_stmt_1142/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 56: 	 branch_block_stmt_1142/forx_xbody_forx_xbody_PhiReq/phi_stmt_1193/$exit
      -- CP-element group 56: 	 branch_block_stmt_1142/forx_xbody_forx_xbody_PhiReq/phi_stmt_1193/phi_stmt_1193_sources/$exit
      -- CP-element group 56: 	 branch_block_stmt_1142/forx_xbody_forx_xbody_PhiReq/phi_stmt_1193/phi_stmt_1193_sources/type_cast_1199/$exit
      -- CP-element group 56: 	 branch_block_stmt_1142/forx_xbody_forx_xbody_PhiReq/phi_stmt_1193/phi_stmt_1193_sources/type_cast_1199/SplitProtocol/$exit
      -- CP-element group 56: 	 branch_block_stmt_1142/forx_xbody_forx_xbody_PhiReq/phi_stmt_1193/phi_stmt_1193_req
      -- 
    phi_stmt_1193_req_2621_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1193_req_2621_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2164_elements(56), ack => phi_stmt_1193_req_1); -- 
    sendB_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_2164_elements(54) & sendB_CP_2164_elements(55);
      gj_sendB_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_2164_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  merge  transition  place  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	53 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (2) 
      -- CP-element group 57: 	 branch_block_stmt_1142/merge_stmt_1192_PhiReqMerge
      -- CP-element group 57: 	 branch_block_stmt_1142/merge_stmt_1192_PhiAck/$entry
      -- 
    sendB_CP_2164_elements(57) <= OrReduce(sendB_CP_2164_elements(53) & sendB_CP_2164_elements(56));
    -- CP-element group 58:  fork  transition  place  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	12 
    -- CP-element group 58: 	16 
    -- CP-element group 58: 	5 
    -- CP-element group 58: 	6 
    -- CP-element group 58: 	8 
    -- CP-element group 58: 	10 
    -- CP-element group 58: 	21 
    -- CP-element group 58: 	26 
    -- CP-element group 58: 	31 
    -- CP-element group 58: 	36 
    -- CP-element group 58: 	41 
    -- CP-element group 58: 	46 
    -- CP-element group 58:  members (53) 
      -- CP-element group 58: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/array_obj_ref_1205_index_scale_1/scale_rename_req
      -- CP-element group 58: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/array_obj_ref_1205_final_index_sum_regn_Sample/req
      -- CP-element group 58: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/array_obj_ref_1205_index_resize_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/ptr_deref_1210_Update/word_access_complete/$entry
      -- CP-element group 58: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/array_obj_ref_1205_index_scale_1/scale_rename_ack
      -- CP-element group 58: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/ptr_deref_1210_Update/word_access_complete/word_0/$entry
      -- CP-element group 58: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/array_obj_ref_1205_final_index_sum_regn_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/addr_of_1206_update_start_
      -- CP-element group 58: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/array_obj_ref_1205_index_computed_1
      -- CP-element group 58: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/$entry
      -- CP-element group 58: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/array_obj_ref_1205_final_index_sum_regn_update_start
      -- CP-element group 58: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/array_obj_ref_1205_index_scale_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/array_obj_ref_1205_index_resize_1/index_resize_req
      -- CP-element group 58: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/array_obj_ref_1205_final_index_sum_regn_Update/req
      -- CP-element group 58: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/addr_of_1206_complete/$entry
      -- CP-element group 58: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/array_obj_ref_1205_index_resize_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/addr_of_1206_complete/req
      -- CP-element group 58: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/array_obj_ref_1205_index_resized_1
      -- CP-element group 58: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/array_obj_ref_1205_index_resize_1/index_resize_ack
      -- CP-element group 58: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/array_obj_ref_1205_final_index_sum_regn_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/array_obj_ref_1205_index_scaled_1
      -- CP-element group 58: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1256_update_start_
      -- CP-element group 58: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/ptr_deref_1210_update_start_
      -- CP-element group 58: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/ptr_deref_1210_Update/word_access_complete/word_0/cr
      -- CP-element group 58: 	 branch_block_stmt_1142/merge_stmt_1192__exit__
      -- CP-element group 58: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320__entry__
      -- CP-element group 58: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1256_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/array_obj_ref_1205_index_scale_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/ptr_deref_1210_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1256_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1263_update_start_
      -- CP-element group 58: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1263_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1263_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1270_update_start_
      -- CP-element group 58: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1270_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1270_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1277_update_start_
      -- CP-element group 58: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1277_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1277_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1284_update_start_
      -- CP-element group 58: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1284_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1284_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1291_update_start_
      -- CP-element group 58: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1291_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1291_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1298_update_start_
      -- CP-element group 58: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1298_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1298_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1305_update_start_
      -- CP-element group 58: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1305_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_1142/assign_stmt_1207_to_assign_stmt_1320/type_cast_1305_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_1142/merge_stmt_1192_PhiAck/$exit
      -- CP-element group 58: 	 branch_block_stmt_1142/merge_stmt_1192_PhiAck/phi_stmt_1193_ack
      -- 
    phi_stmt_1193_ack_2626_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1193_ack_0, ack => sendB_CP_2164_elements(58)); -- 
    req_2258_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2258_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2164_elements(58), ack => array_obj_ref_1205_index_offset_req_0); -- 
    req_2263_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2263_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2164_elements(58), ack => array_obj_ref_1205_index_offset_req_1); -- 
    req_2278_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2278_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2164_elements(58), ack => addr_of_1206_final_reg_req_1); -- 
    cr_2323_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2323_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2164_elements(58), ack => ptr_deref_1210_load_0_req_1); -- 
    cr_2342_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2342_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2164_elements(58), ack => type_cast_1256_inst_req_1); -- 
    cr_2370_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2370_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2164_elements(58), ack => type_cast_1263_inst_req_1); -- 
    cr_2398_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2398_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2164_elements(58), ack => type_cast_1270_inst_req_1); -- 
    cr_2426_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2426_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2164_elements(58), ack => type_cast_1277_inst_req_1); -- 
    cr_2454_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2454_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2164_elements(58), ack => type_cast_1284_inst_req_1); -- 
    cr_2482_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2482_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2164_elements(58), ack => type_cast_1291_inst_req_1); -- 
    cr_2510_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2510_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2164_elements(58), ack => type_cast_1298_inst_req_1); -- 
    cr_2538_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2538_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_2164_elements(58), ack => type_cast_1305_inst_req_1); -- 
    -- CP-element group 59:  merge  transition  place  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	2 
    -- CP-element group 59: 	51 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (16) 
      -- CP-element group 59: 	 $exit
      -- CP-element group 59: 	 branch_block_stmt_1142/branch_block_stmt_1142__exit__
      -- CP-element group 59: 	 branch_block_stmt_1142/return__
      -- CP-element group 59: 	 branch_block_stmt_1142/merge_stmt_1329__exit__
      -- CP-element group 59: 	 branch_block_stmt_1142/$exit
      -- CP-element group 59: 	 branch_block_stmt_1142/merge_stmt_1331__exit__
      -- CP-element group 59: 	 branch_block_stmt_1142/merge_stmt_1329_PhiReqMerge
      -- CP-element group 59: 	 branch_block_stmt_1142/merge_stmt_1329_PhiAck/$entry
      -- CP-element group 59: 	 branch_block_stmt_1142/merge_stmt_1329_PhiAck/$exit
      -- CP-element group 59: 	 branch_block_stmt_1142/merge_stmt_1329_PhiAck/dummy
      -- CP-element group 59: 	 branch_block_stmt_1142/return___PhiReq/$entry
      -- CP-element group 59: 	 branch_block_stmt_1142/return___PhiReq/$exit
      -- CP-element group 59: 	 branch_block_stmt_1142/merge_stmt_1331_PhiReqMerge
      -- CP-element group 59: 	 branch_block_stmt_1142/merge_stmt_1331_PhiAck/$entry
      -- CP-element group 59: 	 branch_block_stmt_1142/merge_stmt_1331_PhiAck/$exit
      -- CP-element group 59: 	 branch_block_stmt_1142/merge_stmt_1331_PhiAck/dummy
      -- 
    sendB_CP_2164_elements(59) <= OrReduce(sendB_CP_2164_elements(2) & sendB_CP_2164_elements(51));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_indvar_1204_resized : std_logic_vector(13 downto 0);
    signal R_indvar_1204_scaled : std_logic_vector(13 downto 0);
    signal array_obj_ref_1205_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1205_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1205_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1205_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1205_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1205_root_address : std_logic_vector(13 downto 0);
    signal arrayidx_1207 : std_logic_vector(31 downto 0);
    signal cmp76_1148 : std_logic_vector(0 downto 0);
    signal conv52_1257 : std_logic_vector(7 downto 0);
    signal conv55_1264 : std_logic_vector(7 downto 0);
    signal conv58_1271 : std_logic_vector(7 downto 0);
    signal conv61_1278 : std_logic_vector(7 downto 0);
    signal conv64_1285 : std_logic_vector(7 downto 0);
    signal conv67_1292 : std_logic_vector(7 downto 0);
    signal conv70_1299 : std_logic_vector(7 downto 0);
    signal conv73_1306 : std_logic_vector(7 downto 0);
    signal exitcond1_1320 : std_logic_vector(0 downto 0);
    signal iNsTr_1_1177 : std_logic_vector(63 downto 0);
    signal indvar_1193 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_1315 : std_logic_vector(63 downto 0);
    signal ptr_deref_1210_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1210_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1210_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1210_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1210_word_offset_0 : std_logic_vector(13 downto 0);
    signal shr15_1223 : std_logic_vector(63 downto 0);
    signal shr21_1229 : std_logic_vector(63 downto 0);
    signal shr27_1235 : std_logic_vector(63 downto 0);
    signal shr33_1241 : std_logic_vector(63 downto 0);
    signal shr39_1247 : std_logic_vector(63 downto 0);
    signal shr45_1253 : std_logic_vector(63 downto 0);
    signal shr9_1217 : std_logic_vector(63 downto 0);
    signal shr_1161 : std_logic_vector(31 downto 0);
    signal shrx_xop_1173 : std_logic_vector(31 downto 0);
    signal tmp4_1211 : std_logic_vector(63 downto 0);
    signal tmp80_1190 : std_logic_vector(63 downto 0);
    signal tmp_1167 : std_logic_vector(0 downto 0);
    signal type_cast_1146_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1159_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1165_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1171_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1181_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1188_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1197_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1199_wire : std_logic_vector(63 downto 0);
    signal type_cast_1215_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1221_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1227_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1233_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1239_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1245_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1251_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1313_wire_constant : std_logic_vector(63 downto 0);
    signal xx_xop_1183 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    array_obj_ref_1205_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1205_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1205_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1205_resized_base_address <= "00000000000000";
    ptr_deref_1210_word_offset_0 <= "00000000000000";
    type_cast_1146_wire_constant <= "00000000000000000000000000000011";
    type_cast_1159_wire_constant <= "00000000000000000000000000000010";
    type_cast_1165_wire_constant <= "00000000000000000000000000000001";
    type_cast_1171_wire_constant <= "11111111111111111111111111111111";
    type_cast_1181_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1188_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1197_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1215_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1221_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1227_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1233_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1239_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1245_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1251_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1313_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    phi_stmt_1193: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1197_wire_constant & type_cast_1199_wire;
      req <= phi_stmt_1193_req_0 & phi_stmt_1193_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1193",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1193_ack_0,
          idata => idata,
          odata => indvar_1193,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1193
    -- flow-through select operator MUX_1189_inst
    tmp80_1190 <= xx_xop_1183 when (tmp_1167(0) /=  '0') else type_cast_1188_wire_constant;
    addr_of_1206_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1206_final_reg_req_0;
      addr_of_1206_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1206_final_reg_req_1;
      addr_of_1206_final_reg_ack_1<= rack(0);
      addr_of_1206_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1206_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1205_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_1207,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1176_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1176_inst_req_0;
      type_cast_1176_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1176_inst_req_1;
      type_cast_1176_inst_ack_1<= rack(0);
      type_cast_1176_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1176_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shrx_xop_1173,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_1_1177,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1199_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1199_inst_req_0;
      type_cast_1199_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1199_inst_req_1;
      type_cast_1199_inst_ack_1<= rack(0);
      type_cast_1199_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1199_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1315,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1199_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1256_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1256_inst_req_0;
      type_cast_1256_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1256_inst_req_1;
      type_cast_1256_inst_ack_1<= rack(0);
      type_cast_1256_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1256_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr45_1253,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv52_1257,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1263_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1263_inst_req_0;
      type_cast_1263_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1263_inst_req_1;
      type_cast_1263_inst_ack_1<= rack(0);
      type_cast_1263_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1263_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr39_1247,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv55_1264,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1270_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1270_inst_req_0;
      type_cast_1270_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1270_inst_req_1;
      type_cast_1270_inst_ack_1<= rack(0);
      type_cast_1270_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1270_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr33_1241,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv58_1271,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1277_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1277_inst_req_0;
      type_cast_1277_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1277_inst_req_1;
      type_cast_1277_inst_ack_1<= rack(0);
      type_cast_1277_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1277_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr27_1235,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv61_1278,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1284_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1284_inst_req_0;
      type_cast_1284_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1284_inst_req_1;
      type_cast_1284_inst_ack_1<= rack(0);
      type_cast_1284_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1284_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr21_1229,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv64_1285,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1291_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1291_inst_req_0;
      type_cast_1291_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1291_inst_req_1;
      type_cast_1291_inst_ack_1<= rack(0);
      type_cast_1291_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1291_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr15_1223,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv67_1292,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1298_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1298_inst_req_0;
      type_cast_1298_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1298_inst_req_1;
      type_cast_1298_inst_ack_1<= rack(0);
      type_cast_1298_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1298_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr9_1217,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv70_1299,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1305_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1305_inst_req_0;
      type_cast_1305_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1305_inst_req_1;
      type_cast_1305_inst_ack_1<= rack(0);
      type_cast_1305_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1305_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp4_1211,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv73_1306,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1205_index_1_rename
    process(R_indvar_1204_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_1204_resized;
      ov(13 downto 0) := iv;
      R_indvar_1204_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1205_index_1_resize
    process(indvar_1193) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_1193;
      ov := iv(13 downto 0);
      R_indvar_1204_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1205_root_address_inst
    process(array_obj_ref_1205_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1205_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1205_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1210_addr_0
    process(ptr_deref_1210_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1210_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1210_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1210_base_resize
    process(arrayidx_1207) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_1207;
      ov := iv(13 downto 0);
      ptr_deref_1210_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1210_gather_scatter
    process(ptr_deref_1210_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1210_data_0;
      ov(63 downto 0) := iv;
      tmp4_1211 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1210_root_address_inst
    process(ptr_deref_1210_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1210_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1210_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1149_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp76_1148;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1149_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1149_branch_req_0,
          ack0 => if_stmt_1149_branch_ack_0,
          ack1 => if_stmt_1149_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1321_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond1_1320;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1321_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1321_branch_req_0,
          ack0 => if_stmt_1321_branch_ack_0,
          ack1 => if_stmt_1321_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u32_u32_1172_inst
    process(shr_1161) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shr_1161, type_cast_1171_wire_constant, tmp_var);
      shrx_xop_1173 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1182_inst
    process(iNsTr_1_1177) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_1_1177, type_cast_1181_wire_constant, tmp_var);
      xx_xop_1183 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1314_inst
    process(indvar_1193) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1193, type_cast_1313_wire_constant, tmp_var);
      indvarx_xnext_1315 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1319_inst
    process(indvarx_xnext_1315, tmp80_1190) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_1315, tmp80_1190, tmp_var);
      exitcond1_1320 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1160_inst
    process(size_buffer) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(size_buffer, type_cast_1159_wire_constant, tmp_var);
      shr_1161 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1216_inst
    process(tmp4_1211) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_1211, type_cast_1215_wire_constant, tmp_var);
      shr9_1217 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1222_inst
    process(tmp4_1211) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_1211, type_cast_1221_wire_constant, tmp_var);
      shr15_1223 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1228_inst
    process(tmp4_1211) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_1211, type_cast_1227_wire_constant, tmp_var);
      shr21_1229 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1234_inst
    process(tmp4_1211) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_1211, type_cast_1233_wire_constant, tmp_var);
      shr27_1235 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1240_inst
    process(tmp4_1211) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_1211, type_cast_1239_wire_constant, tmp_var);
      shr33_1241 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1246_inst
    process(tmp4_1211) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_1211, type_cast_1245_wire_constant, tmp_var);
      shr39_1247 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1252_inst
    process(tmp4_1211) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_1211, type_cast_1251_wire_constant, tmp_var);
      shr45_1253 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1147_inst
    process(size_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(size_buffer, type_cast_1146_wire_constant, tmp_var);
      cmp76_1148 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1166_inst
    process(shr_1161) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(shr_1161, type_cast_1165_wire_constant, tmp_var);
      tmp_1167 <= tmp_var; --
    end process;
    -- shared split operator group (14) : array_obj_ref_1205_index_offset 
    ApIntAdd_group_14: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_1204_scaled;
      array_obj_ref_1205_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1205_index_offset_req_0;
      array_obj_ref_1205_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1205_index_offset_req_1;
      array_obj_ref_1205_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_14_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_14_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_14",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 14
    -- shared load operator group (0) : ptr_deref_1210_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1210_load_0_req_0;
      ptr_deref_1210_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1210_load_0_req_1;
      ptr_deref_1210_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1210_word_address_0;
      ptr_deref_1210_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 3,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(13 downto 0),
          mtag => memory_space_0_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared outport operator group (0) : WPIPE_maxpool_output_pipe_1279_inst WPIPE_maxpool_output_pipe_1265_inst WPIPE_maxpool_output_pipe_1272_inst WPIPE_maxpool_output_pipe_1286_inst WPIPE_maxpool_output_pipe_1293_inst WPIPE_maxpool_output_pipe_1300_inst WPIPE_maxpool_output_pipe_1258_inst WPIPE_maxpool_output_pipe_1307_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 7 downto 0);
      signal update_req, update_ack : BooleanArray( 7 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 7 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 7 downto 0);
      signal guard_vector : std_logic_vector( 7 downto 0);
      constant inBUFs : IntegerArray(7 downto 0) := (7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(7 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false);
      constant guardBuffering: IntegerArray(7 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2);
      -- 
    begin -- 
      sample_req_unguarded(7) <= WPIPE_maxpool_output_pipe_1279_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_maxpool_output_pipe_1265_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_maxpool_output_pipe_1272_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_maxpool_output_pipe_1286_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_maxpool_output_pipe_1293_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_maxpool_output_pipe_1300_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_maxpool_output_pipe_1258_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_maxpool_output_pipe_1307_inst_req_0;
      WPIPE_maxpool_output_pipe_1279_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_maxpool_output_pipe_1265_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_maxpool_output_pipe_1272_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_maxpool_output_pipe_1286_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_maxpool_output_pipe_1293_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_maxpool_output_pipe_1300_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_maxpool_output_pipe_1258_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_maxpool_output_pipe_1307_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(7) <= WPIPE_maxpool_output_pipe_1279_inst_req_1;
      update_req_unguarded(6) <= WPIPE_maxpool_output_pipe_1265_inst_req_1;
      update_req_unguarded(5) <= WPIPE_maxpool_output_pipe_1272_inst_req_1;
      update_req_unguarded(4) <= WPIPE_maxpool_output_pipe_1286_inst_req_1;
      update_req_unguarded(3) <= WPIPE_maxpool_output_pipe_1293_inst_req_1;
      update_req_unguarded(2) <= WPIPE_maxpool_output_pipe_1300_inst_req_1;
      update_req_unguarded(1) <= WPIPE_maxpool_output_pipe_1258_inst_req_1;
      update_req_unguarded(0) <= WPIPE_maxpool_output_pipe_1307_inst_req_1;
      WPIPE_maxpool_output_pipe_1279_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_maxpool_output_pipe_1265_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_maxpool_output_pipe_1272_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_maxpool_output_pipe_1286_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_maxpool_output_pipe_1293_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_maxpool_output_pipe_1300_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_maxpool_output_pipe_1258_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_maxpool_output_pipe_1307_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      data_in <= conv61_1278 & conv55_1264 & conv58_1271 & conv64_1285 & conv67_1292 & conv70_1299 & conv52_1257 & conv73_1306;
      maxpool_output_pipe_write_0_gI: SplitGuardInterface generic map(name => "maxpool_output_pipe_write_0_gI", nreqs => 8, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      maxpool_output_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "maxpool_output_pipe", data_width => 8, num_reqs => 8, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => maxpool_output_pipe_pipe_write_req(0),
          oack => maxpool_output_pipe_pipe_write_ack(0),
          odata => maxpool_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end sendB_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timer is -- 
  generic (tag_length : integer); 
  port ( -- 
    c : out  std_logic_vector(63 downto 0);
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timer;
architecture timer_arch of timer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal c_buffer :  std_logic_vector(63 downto 0);
  signal c_update_enable: Boolean;
  signal timer_CP_307_start: Boolean;
  signal timer_CP_307_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal LOAD_count_81_load_0_req_0 : boolean;
  signal LOAD_count_81_load_0_ack_0 : boolean;
  signal LOAD_count_81_load_0_req_1 : boolean;
  signal LOAD_count_81_load_0_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timer_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timer_CP_307_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timer_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= c_buffer;
  c <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_307_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timer_CP_307_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_307_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timer_CP_307: Block -- control-path 
    signal timer_CP_307_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    timer_CP_307_elements(0) <= timer_CP_307_start;
    timer_CP_307_symbol <= timer_CP_307_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (14) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_82/$entry
      -- CP-element group 0: 	 assign_stmt_82/LOAD_count_81_sample_start_
      -- CP-element group 0: 	 assign_stmt_82/LOAD_count_81_update_start_
      -- CP-element group 0: 	 assign_stmt_82/LOAD_count_81_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_82/LOAD_count_81_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_82/LOAD_count_81_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_82/LOAD_count_81_Sample/word_access_start/$entry
      -- CP-element group 0: 	 assign_stmt_82/LOAD_count_81_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_82/LOAD_count_81_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 assign_stmt_82/LOAD_count_81_Update/$entry
      -- CP-element group 0: 	 assign_stmt_82/LOAD_count_81_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_82/LOAD_count_81_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_82/LOAD_count_81_Update/word_access_complete/word_0/cr
      -- 
    cr_339_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_339_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_307_elements(0), ack => LOAD_count_81_load_0_req_1); -- 
    rr_328_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_328_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_307_elements(0), ack => LOAD_count_81_load_0_req_0); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (5) 
      -- CP-element group 1: 	 assign_stmt_82/LOAD_count_81_sample_completed_
      -- CP-element group 1: 	 assign_stmt_82/LOAD_count_81_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_82/LOAD_count_81_Sample/word_access_start/$exit
      -- CP-element group 1: 	 assign_stmt_82/LOAD_count_81_Sample/word_access_start/word_0/$exit
      -- CP-element group 1: 	 assign_stmt_82/LOAD_count_81_Sample/word_access_start/word_0/ra
      -- 
    ra_329_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_count_81_load_0_ack_0, ack => timer_CP_307_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (11) 
      -- CP-element group 2: 	 $exit
      -- CP-element group 2: 	 assign_stmt_82/$exit
      -- CP-element group 2: 	 assign_stmt_82/LOAD_count_81_update_completed_
      -- CP-element group 2: 	 assign_stmt_82/LOAD_count_81_Update/$exit
      -- CP-element group 2: 	 assign_stmt_82/LOAD_count_81_Update/word_access_complete/$exit
      -- CP-element group 2: 	 assign_stmt_82/LOAD_count_81_Update/word_access_complete/word_0/$exit
      -- CP-element group 2: 	 assign_stmt_82/LOAD_count_81_Update/word_access_complete/word_0/ca
      -- CP-element group 2: 	 assign_stmt_82/LOAD_count_81_Update/LOAD_count_81_Merge/$entry
      -- CP-element group 2: 	 assign_stmt_82/LOAD_count_81_Update/LOAD_count_81_Merge/$exit
      -- CP-element group 2: 	 assign_stmt_82/LOAD_count_81_Update/LOAD_count_81_Merge/merge_req
      -- CP-element group 2: 	 assign_stmt_82/LOAD_count_81_Update/LOAD_count_81_Merge/merge_ack
      -- 
    ca_340_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_count_81_load_0_ack_1, ack => timer_CP_307_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal LOAD_count_81_data_0 : std_logic_vector(63 downto 0);
    signal LOAD_count_81_word_address_0 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    LOAD_count_81_word_address_0 <= "0";
    -- equivalence LOAD_count_81_gather_scatter
    process(LOAD_count_81_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_count_81_data_0;
      ov(63 downto 0) := iv;
      c_buffer <= ov(63 downto 0);
      --
    end process;
    -- shared load operator group (0) : LOAD_count_81_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_count_81_load_0_req_0;
      LOAD_count_81_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_count_81_load_0_req_1;
      LOAD_count_81_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_count_81_word_address_0;
      LOAD_count_81_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(0 downto 0),
          mtag => memory_space_2_lr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(63 downto 0),
          mtag => memory_space_2_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- 
  end Block; -- data_path
  -- 
end timer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timerDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(17 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timerDaemon;
architecture timerDaemon_arch of timerDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal timerDaemon_CP_3928_start: Boolean;
  signal timerDaemon_CP_3928_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal phi_stmt_1965_ack_0 : boolean;
  signal phi_stmt_1965_req_0 : boolean;
  signal do_while_stmt_1963_branch_ack_1 : boolean;
  signal do_while_stmt_1963_branch_ack_0 : boolean;
  signal ADD_u64_u64_1971_inst_req_1 : boolean;
  signal ADD_u64_u64_1971_inst_ack_1 : boolean;
  signal do_while_stmt_1963_branch_req_0 : boolean;
  signal phi_stmt_1965_req_1 : boolean;
  signal ADD_u64_u64_1971_inst_ack_0 : boolean;
  signal ADD_u64_u64_1971_inst_req_0 : boolean;
  signal STORE_count_1973_store_0_ack_1 : boolean;
  signal STORE_count_1973_store_0_req_1 : boolean;
  signal STORE_count_1973_store_0_ack_0 : boolean;
  signal STORE_count_1973_store_0_req_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timerDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timerDaemon_CP_3928_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timerDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timerDaemon_CP_3928_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timerDaemon_CP_3928_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timerDaemon_CP_3928_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timerDaemon_CP_3928: Block -- control-path 
    signal timerDaemon_CP_3928_elements: BooleanArray(39 downto 0);
    -- 
  begin -- 
    timerDaemon_CP_3928_elements(0) <= timerDaemon_CP_3928_start;
    timerDaemon_CP_3928_symbol <= timerDaemon_CP_3928_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 branch_block_stmt_1962/do_while_stmt_1963__entry__
      -- CP-element group 0: 	 branch_block_stmt_1962/branch_block_stmt_1962__entry__
      -- CP-element group 0: 	 branch_block_stmt_1962/$entry
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	39 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 branch_block_stmt_1962/branch_block_stmt_1962__exit__
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_1962/do_while_stmt_1963__exit__
      -- CP-element group 1: 	 branch_block_stmt_1962/$exit
      -- 
    timerDaemon_CP_3928_elements(1) <= timerDaemon_CP_3928_elements(39);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963__entry__
      -- CP-element group 2: 	 branch_block_stmt_1962/do_while_stmt_1963/$entry
      -- 
    timerDaemon_CP_3928_elements(2) <= timerDaemon_CP_3928_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	39 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963__exit__
      -- 
    -- Element group timerDaemon_CP_3928_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_1962/do_while_stmt_1963/loop_back
      -- 
    -- Element group timerDaemon_CP_3928_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	37 
    -- CP-element group 5: 	38 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1962/do_while_stmt_1963/loop_taken/$entry
      -- CP-element group 5: 	 branch_block_stmt_1962/do_while_stmt_1963/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_1962/do_while_stmt_1963/condition_done
      -- 
    timerDaemon_CP_3928_elements(5) <= timerDaemon_CP_3928_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	36 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_1962/do_while_stmt_1963/loop_body_done
      -- 
    timerDaemon_CP_3928_elements(6) <= timerDaemon_CP_3928_elements(36);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	16 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/back_edge_to_loop_body
      -- 
    timerDaemon_CP_3928_elements(7) <= timerDaemon_CP_3928_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	18 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/first_time_through_loop_body
      -- 
    timerDaemon_CP_3928_elements(8) <= timerDaemon_CP_3928_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	35 
    -- CP-element group 9: 	31 
    -- CP-element group 9: 	12 
    -- CP-element group 9: 	13 
    -- CP-element group 9:  members (4) 
      -- CP-element group 9: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/STORE_count_1973_word_address_calculated
      -- CP-element group 9: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/STORE_count_1973_root_address_calculated
      -- 
    -- Element group timerDaemon_CP_3928_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	35 
    -- CP-element group 10: 	15 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/condition_evaluated
      -- 
    condition_evaluated_3952_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_3952_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_3928_elements(10), ack => do_while_stmt_1963_branch_req_0); -- 
    timerDaemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 3);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_3928_elements(35) & timerDaemon_CP_3928_elements(15);
      gj_timerDaemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3928_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	12 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	15 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/phi_stmt_1965_sample_start__ps
      -- 
    timerDaemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_3928_elements(12) & timerDaemon_CP_3928_elements(15);
      gj_timerDaemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3928_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	9 
    -- CP-element group 12: marked-predecessors 
    -- CP-element group 12: 	14 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	11 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/phi_stmt_1965_sample_start_
      -- 
    timerDaemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_3928_elements(9) & timerDaemon_CP_3928_elements(14);
      gj_timerDaemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3928_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	9 
    -- CP-element group 13: marked-predecessors 
    -- CP-element group 13: 	33 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/phi_stmt_1965_update_start__ps
      -- CP-element group 13: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/phi_stmt_1965_update_start_
      -- 
    timerDaemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_3928_elements(9) & timerDaemon_CP_3928_elements(33);
      gj_timerDaemon_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3928_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	36 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	12 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/aggregated_phi_sample_ack
      -- CP-element group 14: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/phi_stmt_1965_sample_completed__ps
      -- CP-element group 14: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/phi_stmt_1965_sample_completed_
      -- 
    -- Element group timerDaemon_CP_3928_elements(14) is bound as output of CP function.
    -- CP-element group 15:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	31 
    -- CP-element group 15: 	10 
    -- CP-element group 15: marked-successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/phi_stmt_1965_update_completed__ps
      -- CP-element group 15: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/aggregated_phi_update_ack
      -- CP-element group 15: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/phi_stmt_1965_update_completed_
      -- 
    -- Element group timerDaemon_CP_3928_elements(15) is bound as output of CP function.
    -- CP-element group 16:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	7 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/phi_stmt_1965_loopback_trigger
      -- 
    timerDaemon_CP_3928_elements(16) <= timerDaemon_CP_3928_elements(7);
    -- CP-element group 17:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (2) 
      -- CP-element group 17: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/phi_stmt_1965_loopback_sample_req
      -- CP-element group 17: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/phi_stmt_1965_loopback_sample_req_ps
      -- 
    phi_stmt_1965_loopback_sample_req_3967_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1965_loopback_sample_req_3967_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_3928_elements(17), ack => phi_stmt_1965_req_1); -- 
    -- Element group timerDaemon_CP_3928_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	8 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/phi_stmt_1965_entry_trigger
      -- 
    timerDaemon_CP_3928_elements(18) <= timerDaemon_CP_3928_elements(8);
    -- CP-element group 19:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (2) 
      -- CP-element group 19: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/phi_stmt_1965_entry_sample_req
      -- CP-element group 19: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/phi_stmt_1965_entry_sample_req_ps
      -- 
    phi_stmt_1965_entry_sample_req_3970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1965_entry_sample_req_3970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_3928_elements(19), ack => phi_stmt_1965_req_0); -- 
    -- Element group timerDaemon_CP_3928_elements(19) is bound as output of CP function.
    -- CP-element group 20:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/phi_stmt_1965_phi_mux_ack
      -- CP-element group 20: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/phi_stmt_1965_phi_mux_ack_ps
      -- 
    phi_stmt_1965_phi_mux_ack_3973_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1965_ack_0, ack => timerDaemon_CP_3928_elements(20)); -- 
    -- CP-element group 21:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (4) 
      -- CP-element group 21: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/type_cast_1968_sample_start__ps
      -- CP-element group 21: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/type_cast_1968_sample_completed__ps
      -- CP-element group 21: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/type_cast_1968_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/type_cast_1968_sample_completed_
      -- 
    -- Element group timerDaemon_CP_3928_elements(21) is bound as output of CP function.
    -- CP-element group 22:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	24 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/type_cast_1968_update_start__ps
      -- CP-element group 22: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/type_cast_1968_update_start_
      -- 
    -- Element group timerDaemon_CP_3928_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	24 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/type_cast_1968_update_completed__ps
      -- 
    timerDaemon_CP_3928_elements(23) <= timerDaemon_CP_3928_elements(24);
    -- CP-element group 24:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	22 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	23 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/type_cast_1968_update_completed_
      -- 
    -- Element group timerDaemon_CP_3928_elements(24) is a control-delay.
    cp_element_24_delay: control_delay_element  generic map(name => " 24_delay", delay_value => 1)  port map(req => timerDaemon_CP_3928_elements(22), ack => timerDaemon_CP_3928_elements(24), clk => clk, reset =>reset);
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/ADD_u64_u64_1971_sample_start__ps
      -- 
    -- Element group timerDaemon_CP_3928_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	28 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/ADD_u64_u64_1971_update_start__ps
      -- 
    -- Element group timerDaemon_CP_3928_elements(26) is bound as output of CP function.
    -- CP-element group 27:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: marked-predecessors 
    -- CP-element group 27: 	29 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/ADD_u64_u64_1971_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/ADD_u64_u64_1971_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/ADD_u64_u64_1971_Sample/rr
      -- 
    rr_3994_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3994_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_3928_elements(27), ack => ADD_u64_u64_1971_inst_req_0); -- 
    timerDaemon_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_3928_elements(25) & timerDaemon_CP_3928_elements(29);
      gj_timerDaemon_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3928_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: marked-predecessors 
    -- CP-element group 28: 	30 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/ADD_u64_u64_1971_Update/cr
      -- CP-element group 28: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/ADD_u64_u64_1971_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/ADD_u64_u64_1971_update_start_
      -- 
    cr_3999_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3999_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_3928_elements(28), ack => ADD_u64_u64_1971_inst_req_1); -- 
    timerDaemon_cp_element_group_28: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_28"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_3928_elements(26) & timerDaemon_CP_3928_elements(30);
      gj_timerDaemon_cp_element_group_28 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3928_elements(28), clk => clk, reset => reset); --
    end block;
    -- CP-element group 29:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29: marked-successors 
    -- CP-element group 29: 	27 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/ADD_u64_u64_1971_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/ADD_u64_u64_1971_sample_completed__ps
      -- CP-element group 29: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/ADD_u64_u64_1971_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/ADD_u64_u64_1971_Sample/ra
      -- 
    ra_3995_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_1971_inst_ack_0, ack => timerDaemon_CP_3928_elements(29)); -- 
    -- CP-element group 30:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30: marked-successors 
    -- CP-element group 30: 	28 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/ADD_u64_u64_1971_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/ADD_u64_u64_1971_Update/ca
      -- CP-element group 30: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/ADD_u64_u64_1971_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/ADD_u64_u64_1971_update_completed__ps
      -- 
    ca_4000_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u64_u64_1971_inst_ack_1, ack => timerDaemon_CP_3928_elements(30)); -- 
    -- CP-element group 31:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	9 
    -- CP-element group 31: 	15 
    -- CP-element group 31: marked-predecessors 
    -- CP-element group 31: 	33 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (9) 
      -- CP-element group 31: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/STORE_count_1973_Sample/STORE_count_1973_Split/$exit
      -- CP-element group 31: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/STORE_count_1973_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/STORE_count_1973_Sample/STORE_count_1973_Split/split_req
      -- CP-element group 31: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/STORE_count_1973_Sample/STORE_count_1973_Split/split_ack
      -- CP-element group 31: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/STORE_count_1973_Sample/word_access_start/$entry
      -- CP-element group 31: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/STORE_count_1973_Sample/word_access_start/word_0/$entry
      -- CP-element group 31: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/STORE_count_1973_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/STORE_count_1973_Sample/STORE_count_1973_Split/$entry
      -- CP-element group 31: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/STORE_count_1973_Sample/word_access_start/word_0/rr
      -- 
    rr_4022_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4022_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_3928_elements(31), ack => STORE_count_1973_store_0_req_0); -- 
    timerDaemon_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 3,1 => 3,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= timerDaemon_CP_3928_elements(9) & timerDaemon_CP_3928_elements(15) & timerDaemon_CP_3928_elements(33);
      gj_timerDaemon_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3928_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	34 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	34 
    -- CP-element group 32:  members (5) 
      -- CP-element group 32: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/STORE_count_1973_update_start_
      -- CP-element group 32: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/STORE_count_1973_Update/word_access_complete/word_0/cr
      -- CP-element group 32: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/STORE_count_1973_Update/word_access_complete/word_0/$entry
      -- CP-element group 32: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/STORE_count_1973_Update/word_access_complete/$entry
      -- CP-element group 32: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/STORE_count_1973_Update/$entry
      -- 
    cr_4033_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4033_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_3928_elements(32), ack => STORE_count_1973_store_0_req_1); -- 
    timerDaemon_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= timerDaemon_CP_3928_elements(34);
      gj_timerDaemon_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3928_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33: marked-successors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: 	13 
    -- CP-element group 33:  members (5) 
      -- CP-element group 33: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/STORE_count_1973_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/STORE_count_1973_Sample/word_access_start/word_0/$exit
      -- CP-element group 33: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/STORE_count_1973_Sample/word_access_start/$exit
      -- CP-element group 33: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/STORE_count_1973_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/STORE_count_1973_Sample/word_access_start/word_0/ra
      -- 
    ra_4023_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_count_1973_store_0_ack_0, ack => timerDaemon_CP_3928_elements(33)); -- 
    -- CP-element group 34:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	32 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34: marked-successors 
    -- CP-element group 34: 	32 
    -- CP-element group 34:  members (5) 
      -- CP-element group 34: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/STORE_count_1973_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/STORE_count_1973_Update/word_access_complete/word_0/ca
      -- CP-element group 34: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/STORE_count_1973_Update/word_access_complete/word_0/$exit
      -- CP-element group 34: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/STORE_count_1973_Update/word_access_complete/$exit
      -- CP-element group 34: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/STORE_count_1973_Update/$exit
      -- 
    ca_4034_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_count_1973_store_0_ack_1, ack => timerDaemon_CP_3928_elements(34)); -- 
    -- CP-element group 35:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	9 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	10 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group timerDaemon_CP_3928_elements(35) is a control-delay.
    cp_element_35_delay: control_delay_element  generic map(name => " 35_delay", delay_value => 1)  port map(req => timerDaemon_CP_3928_elements(9), ack => timerDaemon_CP_3928_elements(35), clk => clk, reset =>reset);
    -- CP-element group 36:  join  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: 	14 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	6 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_1962/do_while_stmt_1963/do_while_stmt_1963_loop_body/$exit
      -- 
    timerDaemon_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 3,1 => 3);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_3928_elements(34) & timerDaemon_CP_3928_elements(14);
      gj_timerDaemon_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_3928_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  transition  input  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	5 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (2) 
      -- CP-element group 37: 	 branch_block_stmt_1962/do_while_stmt_1963/loop_exit/$exit
      -- CP-element group 37: 	 branch_block_stmt_1962/do_while_stmt_1963/loop_exit/ack
      -- 
    ack_4039_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1963_branch_ack_0, ack => timerDaemon_CP_3928_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	5 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (2) 
      -- CP-element group 38: 	 branch_block_stmt_1962/do_while_stmt_1963/loop_taken/$exit
      -- CP-element group 38: 	 branch_block_stmt_1962/do_while_stmt_1963/loop_taken/ack
      -- 
    ack_4043_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1963_branch_ack_1, ack => timerDaemon_CP_3928_elements(38)); -- 
    -- CP-element group 39:  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	3 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	1 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_1962/do_while_stmt_1963/$exit
      -- 
    timerDaemon_CP_3928_elements(39) <= timerDaemon_CP_3928_elements(3);
    timerDaemon_do_while_stmt_1963_terminator_4044: loop_terminator -- 
      generic map (name => " timerDaemon_do_while_stmt_1963_terminator_4044", max_iterations_in_flight =>3) 
      port map(loop_body_exit => timerDaemon_CP_3928_elements(6),loop_continue => timerDaemon_CP_3928_elements(38),loop_terminate => timerDaemon_CP_3928_elements(37),loop_back => timerDaemon_CP_3928_elements(4),loop_exit => timerDaemon_CP_3928_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_1965_phi_seq_4001_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= timerDaemon_CP_3928_elements(18);
      timerDaemon_CP_3928_elements(21)<= src_sample_reqs(0);
      src_sample_acks(0)  <= timerDaemon_CP_3928_elements(21);
      timerDaemon_CP_3928_elements(22)<= src_update_reqs(0);
      src_update_acks(0)  <= timerDaemon_CP_3928_elements(23);
      timerDaemon_CP_3928_elements(19) <= phi_mux_reqs(0);
      triggers(1)  <= timerDaemon_CP_3928_elements(16);
      timerDaemon_CP_3928_elements(25)<= src_sample_reqs(1);
      src_sample_acks(1)  <= timerDaemon_CP_3928_elements(29);
      timerDaemon_CP_3928_elements(26)<= src_update_reqs(1);
      src_update_acks(1)  <= timerDaemon_CP_3928_elements(30);
      timerDaemon_CP_3928_elements(17) <= phi_mux_reqs(1);
      phi_stmt_1965_phi_seq_4001 : phi_sequencer_v2-- 
        generic map (place_capacity => 3, ntriggers => 2, name => "phi_stmt_1965_phi_seq_4001") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => timerDaemon_CP_3928_elements(11), 
          phi_sample_ack => timerDaemon_CP_3928_elements(14), 
          phi_update_req => timerDaemon_CP_3928_elements(13), 
          phi_update_ack => timerDaemon_CP_3928_elements(15), 
          phi_mux_ack => timerDaemon_CP_3928_elements(20), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_3953_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= timerDaemon_CP_3928_elements(7);
        preds(1)  <= timerDaemon_CP_3928_elements(8);
        entry_tmerge_3953 : transition_merge -- 
          generic map(name => " entry_tmerge_3953")
          port map (preds => preds, symbol_out => timerDaemon_CP_3928_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u64_u64_1971_wire : std_logic_vector(63 downto 0);
    signal STORE_count_1973_data_0 : std_logic_vector(63 downto 0);
    signal STORE_count_1973_word_address_0 : std_logic_vector(0 downto 0);
    signal konst_1970_wire_constant : std_logic_vector(63 downto 0);
    signal konst_1977_wire_constant : std_logic_vector(0 downto 0);
    signal ncount_1965 : std_logic_vector(63 downto 0);
    signal type_cast_1968_wire_constant : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    STORE_count_1973_word_address_0 <= "0";
    konst_1970_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    konst_1977_wire_constant <= "1";
    type_cast_1968_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    phi_stmt_1965: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1968_wire_constant & ADD_u64_u64_1971_wire;
      req <= phi_stmt_1965_req_0 & phi_stmt_1965_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1965",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1965_ack_0,
          idata => idata,
          odata => ncount_1965,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1965
    -- equivalence STORE_count_1973_gather_scatter
    process(ncount_1965) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ncount_1965;
      ov(63 downto 0) := iv;
      STORE_count_1973_data_0 <= ov(63 downto 0);
      --
    end process;
    do_while_stmt_1963_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_1977_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1963_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1963_branch_req_0,
          ack0 => do_while_stmt_1963_branch_ack_0,
          ack1 => do_while_stmt_1963_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : ADD_u64_u64_1971_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ncount_1965;
      ADD_u64_u64_1971_wire <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u64_u64_1971_inst_req_0;
      ADD_u64_u64_1971_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u64_u64_1971_inst_req_1;
      ADD_u64_u64_1971_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000000001",
          constant_width => 64,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared store operator group (0) : STORE_count_1973_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 3);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= STORE_count_1973_store_0_req_0;
      STORE_count_1973_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= STORE_count_1973_store_0_req_1;
      STORE_count_1973_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_count_1973_word_address_0;
      data_in <= STORE_count_1973_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 1,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(0 downto 0),
          mdata => memory_space_2_sr_data(63 downto 0),
          mtag => memory_space_2_sr_tag(17 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end timerDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    elapsed_time_pipe_pipe_read_data: out std_logic_vector(63 downto 0);
    elapsed_time_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    elapsed_time_pipe_pipe_read_ack : out std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_write_data: in std_logic_vector(7 downto 0);
    maxpool_input_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_read_data: out std_logic_vector(7 downto 0);
    maxpool_output_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(19 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(2 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(19 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(2 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(19 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(255 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(2 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(255 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(19 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(2 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_2_lr_tag : std_logic_vector(17 downto 0);
  signal memory_space_2_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_2_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(17 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(0 downto 0);
  -- declarations related to module fill_T
  component fill_T is -- 
    generic (tag_length : integer); 
    port ( -- 
      addr : in  std_logic_vector(63 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(255 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(2 downto 0);
      maxpool_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      maxpool_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      maxpool_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module fill_T
  signal fill_T_addr :  std_logic_vector(63 downto 0);
  signal fill_T_in_args    : std_logic_vector(63 downto 0);
  signal fill_T_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal fill_T_tag_out   : std_logic_vector(1 downto 0);
  signal fill_T_start_req : std_logic;
  signal fill_T_start_ack : std_logic;
  signal fill_T_fin_req   : std_logic;
  signal fill_T_fin_ack : std_logic;
  -- caller side aggregated signals for module fill_T
  signal fill_T_call_reqs: std_logic_vector(0 downto 0);
  signal fill_T_call_acks: std_logic_vector(0 downto 0);
  signal fill_T_return_reqs: std_logic_vector(0 downto 0);
  signal fill_T_return_acks: std_logic_vector(0 downto 0);
  signal fill_T_call_data: std_logic_vector(63 downto 0);
  signal fill_T_call_tag: std_logic_vector(0 downto 0);
  signal fill_T_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module maxPool3D
  component maxPool3D is -- 
    generic (tag_length : integer); 
    port ( -- 
      maxpool_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      maxpool_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      maxpool_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      elapsed_time_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      elapsed_time_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      elapsed_time_pipe_pipe_write_data : out  std_logic_vector(63 downto 0);
      maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      fill_T_call_reqs : out  std_logic_vector(0 downto 0);
      fill_T_call_acks : in   std_logic_vector(0 downto 0);
      fill_T_call_data : out  std_logic_vector(63 downto 0);
      fill_T_call_tag  :  out  std_logic_vector(0 downto 0);
      fill_T_return_reqs : out  std_logic_vector(0 downto 0);
      fill_T_return_acks : in   std_logic_vector(0 downto 0);
      fill_T_return_tag :  in   std_logic_vector(0 downto 0);
      timer_call_reqs : out  std_logic_vector(0 downto 0);
      timer_call_acks : in   std_logic_vector(0 downto 0);
      timer_call_tag  :  out  std_logic_vector(1 downto 0);
      timer_return_reqs : out  std_logic_vector(0 downto 0);
      timer_return_acks : in   std_logic_vector(0 downto 0);
      timer_return_data : in   std_logic_vector(63 downto 0);
      timer_return_tag :  in   std_logic_vector(1 downto 0);
      maxPool4_call_reqs : out  std_logic_vector(0 downto 0);
      maxPool4_call_acks : in   std_logic_vector(0 downto 0);
      maxPool4_call_data : out  std_logic_vector(159 downto 0);
      maxPool4_call_tag  :  out  std_logic_vector(0 downto 0);
      maxPool4_return_reqs : out  std_logic_vector(0 downto 0);
      maxPool4_return_acks : in   std_logic_vector(0 downto 0);
      maxPool4_return_data : in   std_logic_vector(7 downto 0);
      maxPool4_return_tag :  in   std_logic_vector(0 downto 0);
      sendB_call_reqs : out  std_logic_vector(0 downto 0);
      sendB_call_acks : in   std_logic_vector(0 downto 0);
      sendB_call_data : out  std_logic_vector(31 downto 0);
      sendB_call_tag  :  out  std_logic_vector(0 downto 0);
      sendB_return_reqs : out  std_logic_vector(0 downto 0);
      sendB_return_acks : in   std_logic_vector(0 downto 0);
      sendB_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module maxPool3D
  signal maxPool3D_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal maxPool3D_tag_out   : std_logic_vector(1 downto 0);
  signal maxPool3D_start_req : std_logic;
  signal maxPool3D_start_ack : std_logic;
  signal maxPool3D_fin_req   : std_logic;
  signal maxPool3D_fin_ack : std_logic;
  -- declarations related to module maxPool4
  component maxPool4 is -- 
    generic (tag_length : integer); 
    port ( -- 
      addr : in  std_logic_vector(31 downto 0);
      addr1 : in  std_logic_vector(31 downto 0);
      addr2 : in  std_logic_vector(31 downto 0);
      addr3 : in  std_logic_vector(31 downto 0);
      addr4 : in  std_logic_vector(31 downto 0);
      output : out  std_logic_vector(7 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(255 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module maxPool4
  signal maxPool4_addr :  std_logic_vector(31 downto 0);
  signal maxPool4_addr1 :  std_logic_vector(31 downto 0);
  signal maxPool4_addr2 :  std_logic_vector(31 downto 0);
  signal maxPool4_addr3 :  std_logic_vector(31 downto 0);
  signal maxPool4_addr4 :  std_logic_vector(31 downto 0);
  signal maxPool4_output :  std_logic_vector(7 downto 0);
  signal maxPool4_in_args    : std_logic_vector(159 downto 0);
  signal maxPool4_out_args   : std_logic_vector(7 downto 0);
  signal maxPool4_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal maxPool4_tag_out   : std_logic_vector(1 downto 0);
  signal maxPool4_start_req : std_logic;
  signal maxPool4_start_ack : std_logic;
  signal maxPool4_fin_req   : std_logic;
  signal maxPool4_fin_ack : std_logic;
  -- caller side aggregated signals for module maxPool4
  signal maxPool4_call_reqs: std_logic_vector(0 downto 0);
  signal maxPool4_call_acks: std_logic_vector(0 downto 0);
  signal maxPool4_return_reqs: std_logic_vector(0 downto 0);
  signal maxPool4_return_acks: std_logic_vector(0 downto 0);
  signal maxPool4_call_data: std_logic_vector(159 downto 0);
  signal maxPool4_call_tag: std_logic_vector(0 downto 0);
  signal maxPool4_return_data: std_logic_vector(7 downto 0);
  signal maxPool4_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module sendB
  component sendB is -- 
    generic (tag_length : integer); 
    port ( -- 
      size : in  std_logic_vector(31 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
      maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module sendB
  signal sendB_size :  std_logic_vector(31 downto 0);
  signal sendB_in_args    : std_logic_vector(31 downto 0);
  signal sendB_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal sendB_tag_out   : std_logic_vector(1 downto 0);
  signal sendB_start_req : std_logic;
  signal sendB_start_ack : std_logic;
  signal sendB_fin_req   : std_logic;
  signal sendB_fin_ack : std_logic;
  -- caller side aggregated signals for module sendB
  signal sendB_call_reqs: std_logic_vector(0 downto 0);
  signal sendB_call_acks: std_logic_vector(0 downto 0);
  signal sendB_return_reqs: std_logic_vector(0 downto 0);
  signal sendB_return_acks: std_logic_vector(0 downto 0);
  signal sendB_call_data: std_logic_vector(31 downto 0);
  signal sendB_call_tag: std_logic_vector(0 downto 0);
  signal sendB_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module timer
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      c : out  std_logic_vector(63 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timer
  signal timer_c :  std_logic_vector(63 downto 0);
  signal timer_out_args   : std_logic_vector(63 downto 0);
  signal timer_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal timer_tag_out   : std_logic_vector(2 downto 0);
  signal timer_start_req : std_logic;
  signal timer_start_ack : std_logic;
  signal timer_fin_req   : std_logic;
  signal timer_fin_ack : std_logic;
  -- caller side aggregated signals for module timer
  signal timer_call_reqs: std_logic_vector(0 downto 0);
  signal timer_call_acks: std_logic_vector(0 downto 0);
  signal timer_return_reqs: std_logic_vector(0 downto 0);
  signal timer_return_acks: std_logic_vector(0 downto 0);
  signal timer_call_tag: std_logic_vector(1 downto 0);
  signal timer_return_data: std_logic_vector(63 downto 0);
  signal timer_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module timerDaemon
  component timerDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(17 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timerDaemon
  signal timerDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal timerDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal timerDaemon_start_req : std_logic;
  signal timerDaemon_start_ack : std_logic;
  signal timerDaemon_fin_req   : std_logic;
  signal timerDaemon_fin_ack : std_logic;
  -- aggregate signals for write to pipe elapsed_time_pipe
  signal elapsed_time_pipe_pipe_write_data: std_logic_vector(63 downto 0);
  signal elapsed_time_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal elapsed_time_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe maxpool_input_pipe
  signal maxpool_input_pipe_pipe_read_data: std_logic_vector(15 downto 0);
  signal maxpool_input_pipe_pipe_read_req: std_logic_vector(1 downto 0);
  signal maxpool_input_pipe_pipe_read_ack: std_logic_vector(1 downto 0);
  -- aggregate signals for write to pipe maxpool_output_pipe
  signal maxpool_output_pipe_pipe_write_data: std_logic_vector(15 downto 0);
  signal maxpool_output_pipe_pipe_write_req: std_logic_vector(1 downto 0);
  signal maxpool_output_pipe_pipe_write_ack: std_logic_vector(1 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module fill_T
  fill_T_addr <= fill_T_in_args(63 downto 0);
  -- call arbiter for module fill_T
  fill_T_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => fill_T_call_reqs,
      call_acks => fill_T_call_acks,
      return_reqs => fill_T_return_reqs,
      return_acks => fill_T_return_acks,
      call_data  => fill_T_call_data,
      call_tag  => fill_T_call_tag,
      return_tag  => fill_T_return_tag,
      call_mtag => fill_T_tag_in,
      return_mtag => fill_T_tag_out,
      call_mreq => fill_T_start_req,
      call_mack => fill_T_start_ack,
      return_mreq => fill_T_fin_req,
      return_mack => fill_T_fin_ack,
      call_mdata => fill_T_in_args,
      clk => clk, 
      reset => reset --
    ); --
  fill_T_instance:fill_T-- 
    generic map(tag_length => 2)
    port map(-- 
      addr => fill_T_addr,
      start_req => fill_T_start_req,
      start_ack => fill_T_start_ack,
      fin_req => fill_T_fin_req,
      fin_ack => fill_T_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(13 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(255 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(19 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(2 downto 0),
      maxpool_input_pipe_pipe_read_req => maxpool_input_pipe_pipe_read_req(1 downto 1),
      maxpool_input_pipe_pipe_read_ack => maxpool_input_pipe_pipe_read_ack(1 downto 1),
      maxpool_input_pipe_pipe_read_data => maxpool_input_pipe_pipe_read_data(15 downto 8),
      tag_in => fill_T_tag_in,
      tag_out => fill_T_tag_out-- 
    ); -- 
  -- module maxPool3D
  maxPool3D_instance:maxPool3D-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => maxPool3D_start_req,
      start_ack => maxPool3D_start_ack,
      fin_req => maxPool3D_fin_req,
      fin_ack => maxPool3D_fin_ack,
      clk => clk,
      reset => reset,
      maxpool_input_pipe_pipe_read_req => maxpool_input_pipe_pipe_read_req(0 downto 0),
      maxpool_input_pipe_pipe_read_ack => maxpool_input_pipe_pipe_read_ack(0 downto 0),
      maxpool_input_pipe_pipe_read_data => maxpool_input_pipe_pipe_read_data(7 downto 0),
      elapsed_time_pipe_pipe_write_req => elapsed_time_pipe_pipe_write_req(0 downto 0),
      elapsed_time_pipe_pipe_write_ack => elapsed_time_pipe_pipe_write_ack(0 downto 0),
      elapsed_time_pipe_pipe_write_data => elapsed_time_pipe_pipe_write_data(63 downto 0),
      maxpool_output_pipe_pipe_write_req => maxpool_output_pipe_pipe_write_req(0 downto 0),
      maxpool_output_pipe_pipe_write_ack => maxpool_output_pipe_pipe_write_ack(0 downto 0),
      maxpool_output_pipe_pipe_write_data => maxpool_output_pipe_pipe_write_data(7 downto 0),
      fill_T_call_reqs => fill_T_call_reqs(0 downto 0),
      fill_T_call_acks => fill_T_call_acks(0 downto 0),
      fill_T_call_data => fill_T_call_data(63 downto 0),
      fill_T_call_tag => fill_T_call_tag(0 downto 0),
      fill_T_return_reqs => fill_T_return_reqs(0 downto 0),
      fill_T_return_acks => fill_T_return_acks(0 downto 0),
      fill_T_return_tag => fill_T_return_tag(0 downto 0),
      timer_call_reqs => timer_call_reqs(0 downto 0),
      timer_call_acks => timer_call_acks(0 downto 0),
      timer_call_tag => timer_call_tag(1 downto 0),
      timer_return_reqs => timer_return_reqs(0 downto 0),
      timer_return_acks => timer_return_acks(0 downto 0),
      timer_return_data => timer_return_data(63 downto 0),
      timer_return_tag => timer_return_tag(1 downto 0),
      maxPool4_call_reqs => maxPool4_call_reqs(0 downto 0),
      maxPool4_call_acks => maxPool4_call_acks(0 downto 0),
      maxPool4_call_data => maxPool4_call_data(159 downto 0),
      maxPool4_call_tag => maxPool4_call_tag(0 downto 0),
      maxPool4_return_reqs => maxPool4_return_reqs(0 downto 0),
      maxPool4_return_acks => maxPool4_return_acks(0 downto 0),
      maxPool4_return_data => maxPool4_return_data(7 downto 0),
      maxPool4_return_tag => maxPool4_return_tag(0 downto 0),
      sendB_call_reqs => sendB_call_reqs(0 downto 0),
      sendB_call_acks => sendB_call_acks(0 downto 0),
      sendB_call_data => sendB_call_data(31 downto 0),
      sendB_call_tag => sendB_call_tag(0 downto 0),
      sendB_return_reqs => sendB_return_reqs(0 downto 0),
      sendB_return_acks => sendB_return_acks(0 downto 0),
      sendB_return_tag => sendB_return_tag(0 downto 0),
      tag_in => maxPool3D_tag_in,
      tag_out => maxPool3D_tag_out-- 
    ); -- 
  -- module will be run forever 
  maxPool3D_tag_in <= (others => '0');
  maxPool3D_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => maxPool3D_start_req, start_ack => maxPool3D_start_ack,  fin_req => maxPool3D_fin_req,  fin_ack => maxPool3D_fin_ack);
  -- module maxPool4
  maxPool4_addr <= maxPool4_in_args(159 downto 128);
  maxPool4_addr1 <= maxPool4_in_args(127 downto 96);
  maxPool4_addr2 <= maxPool4_in_args(95 downto 64);
  maxPool4_addr3 <= maxPool4_in_args(63 downto 32);
  maxPool4_addr4 <= maxPool4_in_args(31 downto 0);
  maxPool4_out_args <= maxPool4_output ;
  -- call arbiter for module maxPool4
  maxPool4_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 160,
      return_data_width => 8,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => maxPool4_call_reqs,
      call_acks => maxPool4_call_acks,
      return_reqs => maxPool4_return_reqs,
      return_acks => maxPool4_return_acks,
      call_data  => maxPool4_call_data,
      call_tag  => maxPool4_call_tag,
      return_tag  => maxPool4_return_tag,
      call_mtag => maxPool4_tag_in,
      return_mtag => maxPool4_tag_out,
      return_data =>maxPool4_return_data,
      call_mreq => maxPool4_start_req,
      call_mack => maxPool4_start_ack,
      return_mreq => maxPool4_fin_req,
      return_mack => maxPool4_fin_ack,
      call_mdata => maxPool4_in_args,
      return_mdata => maxPool4_out_args,
      clk => clk, 
      reset => reset --
    ); --
  maxPool4_instance:maxPool4-- 
    generic map(tag_length => 2)
    port map(-- 
      addr => maxPool4_addr,
      addr1 => maxPool4_addr1,
      addr2 => maxPool4_addr2,
      addr3 => maxPool4_addr3,
      addr4 => maxPool4_addr4,
      output => maxPool4_output,
      start_req => maxPool4_start_req,
      start_ack => maxPool4_start_ack,
      fin_req => maxPool4_fin_req,
      fin_ack => maxPool4_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(13 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(19 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(255 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(2 downto 0),
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(13 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(63 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(19 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(2 downto 0),
      tag_in => maxPool4_tag_in,
      tag_out => maxPool4_tag_out-- 
    ); -- 
  -- module sendB
  sendB_size <= sendB_in_args(31 downto 0);
  -- call arbiter for module sendB
  sendB_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 32,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => sendB_call_reqs,
      call_acks => sendB_call_acks,
      return_reqs => sendB_return_reqs,
      return_acks => sendB_return_acks,
      call_data  => sendB_call_data,
      call_tag  => sendB_call_tag,
      return_tag  => sendB_return_tag,
      call_mtag => sendB_tag_in,
      return_mtag => sendB_tag_out,
      call_mreq => sendB_start_req,
      call_mack => sendB_start_ack,
      return_mreq => sendB_fin_req,
      return_mack => sendB_fin_ack,
      call_mdata => sendB_in_args,
      clk => clk, 
      reset => reset --
    ); --
  sendB_instance:sendB-- 
    generic map(tag_length => 2)
    port map(-- 
      size => sendB_size,
      start_req => sendB_start_req,
      start_ack => sendB_start_ack,
      fin_req => sendB_fin_req,
      fin_ack => sendB_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(13 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(19 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(2 downto 0),
      maxpool_output_pipe_pipe_write_req => maxpool_output_pipe_pipe_write_req(1 downto 1),
      maxpool_output_pipe_pipe_write_ack => maxpool_output_pipe_pipe_write_ack(1 downto 1),
      maxpool_output_pipe_pipe_write_data => maxpool_output_pipe_pipe_write_data(15 downto 8),
      tag_in => sendB_tag_in,
      tag_out => sendB_tag_out-- 
    ); -- 
  -- module timer
  timer_out_args <= timer_c ;
  -- call arbiter for module timer
  timer_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargs", num_reqs => 1,
      return_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => timer_call_reqs,
      call_acks => timer_call_acks,
      return_reqs => timer_return_reqs,
      return_acks => timer_return_acks,
      call_tag  => timer_call_tag,
      return_tag  => timer_return_tag,
      call_mtag => timer_tag_in,
      return_mtag => timer_tag_out,
      return_data =>timer_return_data,
      call_mreq => timer_start_req,
      call_mack => timer_start_ack,
      return_mreq => timer_fin_req,
      return_mack => timer_fin_ack,
      return_mdata => timer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  timer_instance:timer-- 
    generic map(tag_length => 3)
    port map(-- 
      c => timer_c,
      start_req => timer_start_req,
      start_ack => timer_start_ack,
      fin_req => timer_fin_req,
      fin_ack => timer_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_2_lr_req => memory_space_2_lr_req(0 downto 0),
      memory_space_2_lr_ack => memory_space_2_lr_ack(0 downto 0),
      memory_space_2_lr_addr => memory_space_2_lr_addr(0 downto 0),
      memory_space_2_lr_tag => memory_space_2_lr_tag(17 downto 0),
      memory_space_2_lc_req => memory_space_2_lc_req(0 downto 0),
      memory_space_2_lc_ack => memory_space_2_lc_ack(0 downto 0),
      memory_space_2_lc_data => memory_space_2_lc_data(63 downto 0),
      memory_space_2_lc_tag => memory_space_2_lc_tag(0 downto 0),
      tag_in => timer_tag_in,
      tag_out => timer_tag_out-- 
    ); -- 
  -- module timerDaemon
  timerDaemon_instance:timerDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => timerDaemon_start_req,
      start_ack => timerDaemon_start_ack,
      fin_req => timerDaemon_fin_req,
      fin_ack => timerDaemon_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_2_sr_req => memory_space_2_sr_req(0 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(0 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(0 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(63 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(17 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(0 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(0 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(0 downto 0),
      tag_in => timerDaemon_tag_in,
      tag_out => timerDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  timerDaemon_tag_in <= (others => '0');
  timerDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => timerDaemon_start_req, start_ack => timerDaemon_start_ack,  fin_req => timerDaemon_fin_req,  fin_ack => timerDaemon_fin_ack);
  elapsed_time_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe elapsed_time_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => elapsed_time_pipe_pipe_read_req,
      read_ack => elapsed_time_pipe_pipe_read_ack,
      read_data => elapsed_time_pipe_pipe_read_data,
      write_req => elapsed_time_pipe_pipe_write_req,
      write_ack => elapsed_time_pipe_pipe_write_ack,
      write_data => elapsed_time_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  maxpool_input_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe maxpool_input_pipe",
      num_reads => 2,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => maxpool_input_pipe_pipe_read_req,
      read_ack => maxpool_input_pipe_pipe_read_ack,
      read_data => maxpool_input_pipe_pipe_read_data,
      write_req => maxpool_input_pipe_pipe_write_req,
      write_ack => maxpool_input_pipe_pipe_write_ack,
      write_data => maxpool_input_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  maxpool_output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe maxpool_output_pipe",
      num_reads => 1,
      num_writes => 2,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => maxpool_output_pipe_pipe_read_req,
      read_ack => maxpool_output_pipe_pipe_read_ack,
      read_data => maxpool_output_pipe_pipe_read_data,
      write_req => maxpool_output_pipe_pipe_write_req,
      write_ack => maxpool_output_pipe_pipe_write_ack,
      write_data => maxpool_output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  MemorySpace_memory_space_0: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 3,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_1: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 256,
      tag_width => 3,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 256
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_2: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_2",
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_2_lr_addr,
      lr_req_in => memory_space_2_lr_req,
      lr_ack_out => memory_space_2_lr_ack,
      lr_tag_in => memory_space_2_lr_tag,
      lc_req_in => memory_space_2_lc_req,
      lc_ack_out => memory_space_2_lc_ack,
      lc_data_out => memory_space_2_lc_data,
      lc_tag_out => memory_space_2_lc_tag,
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
